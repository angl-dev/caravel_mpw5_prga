VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2600.000 BY 2600.000 ;
  PIN ipin_x0y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END ipin_x0y1_0
  PIN ipin_x0y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END ipin_x0y1_1
  PIN ipin_x0y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END ipin_x0y2_0
  PIN ipin_x0y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END ipin_x0y2_1
  PIN ipin_x0y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END ipin_x0y3_0
  PIN ipin_x0y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END ipin_x0y3_1
  PIN ipin_x0y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END ipin_x0y4_0
  PIN ipin_x0y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END ipin_x0y4_1
  PIN ipin_x0y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END ipin_x0y5_0
  PIN ipin_x0y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END ipin_x0y5_1
  PIN ipin_x0y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END ipin_x0y6_0
  PIN ipin_x0y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END ipin_x0y6_1
  PIN ipin_x0y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END ipin_x0y7_0
  PIN ipin_x0y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END ipin_x0y7_1
  PIN ipin_x0y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END ipin_x0y8_0
  PIN ipin_x0y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END ipin_x0y8_1
  PIN ipin_x1y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 2596.000 27.050 2600.000 ;
    END
  END ipin_x1y9_0
  PIN ipin_x1y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 2596.000 80.870 2600.000 ;
    END
  END ipin_x1y9_1
  PIN ipin_x2y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 2596.000 135.150 2600.000 ;
    END
  END ipin_x2y9_0
  PIN ipin_x2y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 2596.000 189.430 2600.000 ;
    END
  END ipin_x2y9_1
  PIN ipin_x3y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 2596.000 243.710 2600.000 ;
    END
  END ipin_x3y9_0
  PIN ipin_x3y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 2596.000 297.530 2600.000 ;
    END
  END ipin_x3y9_1
  PIN ipin_x4y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 2596.000 351.810 2600.000 ;
    END
  END ipin_x4y9_0
  PIN ipin_x4y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 2596.000 406.090 2600.000 ;
    END
  END ipin_x4y9_1
  PIN ipin_x5y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 2596.000 460.370 2600.000 ;
    END
  END ipin_x5y9_0
  PIN ipin_x5y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 2596.000 514.190 2600.000 ;
    END
  END ipin_x5y9_1
  PIN ipin_x6y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 2596.000 568.470 2600.000 ;
    END
  END ipin_x6y9_0
  PIN ipin_x6y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 2596.000 622.750 2600.000 ;
    END
  END ipin_x6y9_1
  PIN ipin_x7y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 2596.000 677.030 2600.000 ;
    END
  END ipin_x7y9_0
  PIN ipin_x7y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 2596.000 730.850 2600.000 ;
    END
  END ipin_x7y9_1
  PIN ipin_x8y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 2596.000 785.130 2600.000 ;
    END
  END ipin_x8y9_0
  PIN ipin_x8y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 2596.000 839.410 2600.000 ;
    END
  END ipin_x8y9_1
  PIN ipin_x9y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 26.560 2600.000 27.160 ;
    END
  END ipin_x9y1_0
  PIN ipin_x9y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 80.280 2600.000 80.880 ;
    END
  END ipin_x9y1_1
  PIN ipin_x9y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 134.680 2600.000 135.280 ;
    END
  END ipin_x9y2_0
  PIN ipin_x9y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 189.080 2600.000 189.680 ;
    END
  END ipin_x9y2_1
  PIN ipin_x9y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 242.800 2600.000 243.400 ;
    END
  END ipin_x9y3_0
  PIN ipin_x9y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 297.200 2600.000 297.800 ;
    END
  END ipin_x9y3_1
  PIN ipin_x9y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 351.600 2600.000 352.200 ;
    END
  END ipin_x9y4_0
  PIN ipin_x9y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 405.320 2600.000 405.920 ;
    END
  END ipin_x9y4_1
  PIN ipin_x9y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 459.720 2600.000 460.320 ;
    END
  END ipin_x9y5_0
  PIN ipin_x9y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 514.120 2600.000 514.720 ;
    END
  END ipin_x9y5_1
  PIN ipin_x9y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 567.840 2600.000 568.440 ;
    END
  END ipin_x9y6_0
  PIN ipin_x9y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 622.240 2600.000 622.840 ;
    END
  END ipin_x9y6_1
  PIN ipin_x9y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 676.640 2600.000 677.240 ;
    END
  END ipin_x9y7_0
  PIN ipin_x9y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 730.360 2600.000 730.960 ;
    END
  END ipin_x9y7_1
  PIN ipin_x9y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 784.760 2600.000 785.360 ;
    END
  END ipin_x9y8_0
  PIN ipin_x9y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 839.160 2600.000 839.760 ;
    END
  END ipin_x9y8_1
  PIN oe_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1759.880 4.000 1760.480 ;
    END
  END oe_x0y1_0
  PIN oe_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1814.280 4.000 1814.880 ;
    END
  END oe_x0y1_1
  PIN oe_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1868.000 4.000 1868.600 ;
    END
  END oe_x0y2_0
  PIN oe_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1922.400 4.000 1923.000 ;
    END
  END oe_x0y2_1
  PIN oe_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1976.800 4.000 1977.400 ;
    END
  END oe_x0y3_0
  PIN oe_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2030.520 4.000 2031.120 ;
    END
  END oe_x0y3_1
  PIN oe_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2084.920 4.000 2085.520 ;
    END
  END oe_x0y4_0
  PIN oe_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2139.320 4.000 2139.920 ;
    END
  END oe_x0y4_1
  PIN oe_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2193.040 4.000 2193.640 ;
    END
  END oe_x0y5_0
  PIN oe_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2247.440 4.000 2248.040 ;
    END
  END oe_x0y5_1
  PIN oe_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2301.840 4.000 2302.440 ;
    END
  END oe_x0y6_0
  PIN oe_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2355.560 4.000 2356.160 ;
    END
  END oe_x0y6_1
  PIN oe_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2409.960 4.000 2410.560 ;
    END
  END oe_x0y7_0
  PIN oe_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2464.360 4.000 2464.960 ;
    END
  END oe_x0y7_1
  PIN oe_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2518.080 4.000 2518.680 ;
    END
  END oe_x0y8_0
  PIN oe_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2572.480 4.000 2573.080 ;
    END
  END oe_x0y8_1
  PIN oe_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.050 2596.000 1760.330 2600.000 ;
    END
  END oe_x1y9_0
  PIN oe_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.870 2596.000 1814.150 2600.000 ;
    END
  END oe_x1y9_1
  PIN oe_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 2596.000 1868.430 2600.000 ;
    END
  END oe_x2y9_0
  PIN oe_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 2596.000 1922.710 2600.000 ;
    END
  END oe_x2y9_1
  PIN oe_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.710 2596.000 1976.990 2600.000 ;
    END
  END oe_x3y9_0
  PIN oe_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.530 2596.000 2030.810 2600.000 ;
    END
  END oe_x3y9_1
  PIN oe_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.810 2596.000 2085.090 2600.000 ;
    END
  END oe_x4y9_0
  PIN oe_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.090 2596.000 2139.370 2600.000 ;
    END
  END oe_x4y9_1
  PIN oe_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.370 2596.000 2193.650 2600.000 ;
    END
  END oe_x5y9_0
  PIN oe_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.190 2596.000 2247.470 2600.000 ;
    END
  END oe_x5y9_1
  PIN oe_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.470 2596.000 2301.750 2600.000 ;
    END
  END oe_x6y9_0
  PIN oe_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.750 2596.000 2356.030 2600.000 ;
    END
  END oe_x6y9_1
  PIN oe_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.030 2596.000 2410.310 2600.000 ;
    END
  END oe_x7y9_0
  PIN oe_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.850 2596.000 2464.130 2600.000 ;
    END
  END oe_x7y9_1
  PIN oe_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.130 2596.000 2518.410 2600.000 ;
    END
  END oe_x8y9_0
  PIN oe_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2572.410 2596.000 2572.690 2600.000 ;
    END
  END oe_x8y9_1
  PIN oe_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1759.880 2600.000 1760.480 ;
    END
  END oe_x9y1_0
  PIN oe_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1814.280 2600.000 1814.880 ;
    END
  END oe_x9y1_1
  PIN oe_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1868.000 2600.000 1868.600 ;
    END
  END oe_x9y2_0
  PIN oe_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1922.400 2600.000 1923.000 ;
    END
  END oe_x9y2_1
  PIN oe_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1976.800 2600.000 1977.400 ;
    END
  END oe_x9y3_0
  PIN oe_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2030.520 2600.000 2031.120 ;
    END
  END oe_x9y3_1
  PIN oe_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2084.920 2600.000 2085.520 ;
    END
  END oe_x9y4_0
  PIN oe_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2139.320 2600.000 2139.920 ;
    END
  END oe_x9y4_1
  PIN oe_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2193.040 2600.000 2193.640 ;
    END
  END oe_x9y5_0
  PIN oe_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2247.440 2600.000 2248.040 ;
    END
  END oe_x9y5_1
  PIN oe_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2301.840 2600.000 2302.440 ;
    END
  END oe_x9y6_0
  PIN oe_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2355.560 2600.000 2356.160 ;
    END
  END oe_x9y6_1
  PIN oe_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2409.960 2600.000 2410.560 ;
    END
  END oe_x9y7_0
  PIN oe_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2464.360 2600.000 2464.960 ;
    END
  END oe_x9y7_1
  PIN oe_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2518.080 2600.000 2518.680 ;
    END
  END oe_x9y8_0
  PIN oe_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2572.480 2600.000 2573.080 ;
    END
  END oe_x9y8_1
  PIN opin_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END opin_x0y1_0
  PIN opin_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.280 4.000 947.880 ;
    END
  END opin_x0y1_1
  PIN opin_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END opin_x0y2_0
  PIN opin_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1055.400 4.000 1056.000 ;
    END
  END opin_x0y2_1
  PIN opin_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.800 4.000 1110.400 ;
    END
  END opin_x0y3_0
  PIN opin_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1164.200 4.000 1164.800 ;
    END
  END opin_x0y3_1
  PIN opin_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.920 4.000 1218.520 ;
    END
  END opin_x0y4_0
  PIN opin_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1272.320 4.000 1272.920 ;
    END
  END opin_x0y4_1
  PIN opin_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.720 4.000 1327.320 ;
    END
  END opin_x0y5_0
  PIN opin_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END opin_x0y5_1
  PIN opin_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END opin_x0y6_0
  PIN opin_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END opin_x0y6_1
  PIN opin_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1542.960 4.000 1543.560 ;
    END
  END opin_x0y7_0
  PIN opin_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1597.360 4.000 1597.960 ;
    END
  END opin_x0y7_1
  PIN opin_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1651.760 4.000 1652.360 ;
    END
  END opin_x0y8_0
  PIN opin_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1705.480 4.000 1706.080 ;
    END
  END opin_x0y8_1
  PIN opin_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 2596.000 893.690 2600.000 ;
    END
  END opin_x1y9_0
  PIN opin_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 2596.000 947.510 2600.000 ;
    END
  END opin_x1y9_1
  PIN opin_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 2596.000 1001.790 2600.000 ;
    END
  END opin_x2y9_0
  PIN opin_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 2596.000 1056.070 2600.000 ;
    END
  END opin_x2y9_1
  PIN opin_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 2596.000 1110.350 2600.000 ;
    END
  END opin_x3y9_0
  PIN opin_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 2596.000 1164.170 2600.000 ;
    END
  END opin_x3y9_1
  PIN opin_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 2596.000 1218.450 2600.000 ;
    END
  END opin_x4y9_0
  PIN opin_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 2596.000 1272.730 2600.000 ;
    END
  END opin_x4y9_1
  PIN opin_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 2596.000 1327.010 2600.000 ;
    END
  END opin_x5y9_0
  PIN opin_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 2596.000 1380.830 2600.000 ;
    END
  END opin_x5y9_1
  PIN opin_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.830 2596.000 1435.110 2600.000 ;
    END
  END opin_x6y9_0
  PIN opin_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 2596.000 1489.390 2600.000 ;
    END
  END opin_x6y9_1
  PIN opin_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.390 2596.000 1543.670 2600.000 ;
    END
  END opin_x7y9_0
  PIN opin_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 2596.000 1597.490 2600.000 ;
    END
  END opin_x7y9_1
  PIN opin_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.490 2596.000 1651.770 2600.000 ;
    END
  END opin_x8y9_0
  PIN opin_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 2596.000 1706.050 2600.000 ;
    END
  END opin_x8y9_1
  PIN opin_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 892.880 2600.000 893.480 ;
    END
  END opin_x9y1_0
  PIN opin_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 947.280 2600.000 947.880 ;
    END
  END opin_x9y1_1
  PIN opin_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1001.680 2600.000 1002.280 ;
    END
  END opin_x9y2_0
  PIN opin_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1055.400 2600.000 1056.000 ;
    END
  END opin_x9y2_1
  PIN opin_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1109.800 2600.000 1110.400 ;
    END
  END opin_x9y3_0
  PIN opin_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1164.200 2600.000 1164.800 ;
    END
  END opin_x9y3_1
  PIN opin_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1217.920 2600.000 1218.520 ;
    END
  END opin_x9y4_0
  PIN opin_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1272.320 2600.000 1272.920 ;
    END
  END opin_x9y4_1
  PIN opin_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1326.720 2600.000 1327.320 ;
    END
  END opin_x9y5_0
  PIN opin_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1380.440 2600.000 1381.040 ;
    END
  END opin_x9y5_1
  PIN opin_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1434.840 2600.000 1435.440 ;
    END
  END opin_x9y6_0
  PIN opin_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1489.240 2600.000 1489.840 ;
    END
  END opin_x9y6_1
  PIN opin_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1542.960 2600.000 1543.560 ;
    END
  END opin_x9y7_0
  PIN opin_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1597.360 2600.000 1597.960 ;
    END
  END opin_x9y7_1
  PIN opin_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1651.760 2600.000 1652.360 ;
    END
  END opin_x9y8_0
  PIN opin_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1705.480 2600.000 1706.080 ;
    END
  END opin_x9y8_1
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END prog_clk
  PIN prog_din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END prog_din
  PIN prog_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END prog_done
  PIN prog_dout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 4.000 ;
    END
  END prog_dout
  PIN prog_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.810 0.000 1671.090 4.000 ;
    END
  END prog_rst
  PIN prog_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.490 0.000 2042.770 4.000 ;
    END
  END prog_we
  PIN prog_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.710 0.000 2413.990 4.000 ;
    END
  END prog_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 2586.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 2586.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 2586.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2595.175 2586.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 2599.390 2587.360 ;
      LAYER met2 ;
        RECT 6.990 2595.720 26.490 2596.650 ;
        RECT 27.330 2595.720 80.310 2596.650 ;
        RECT 81.150 2595.720 134.590 2596.650 ;
        RECT 135.430 2595.720 188.870 2596.650 ;
        RECT 189.710 2595.720 243.150 2596.650 ;
        RECT 243.990 2595.720 296.970 2596.650 ;
        RECT 297.810 2595.720 351.250 2596.650 ;
        RECT 352.090 2595.720 405.530 2596.650 ;
        RECT 406.370 2595.720 459.810 2596.650 ;
        RECT 460.650 2595.720 513.630 2596.650 ;
        RECT 514.470 2595.720 567.910 2596.650 ;
        RECT 568.750 2595.720 622.190 2596.650 ;
        RECT 623.030 2595.720 676.470 2596.650 ;
        RECT 677.310 2595.720 730.290 2596.650 ;
        RECT 731.130 2595.720 784.570 2596.650 ;
        RECT 785.410 2595.720 838.850 2596.650 ;
        RECT 839.690 2595.720 893.130 2596.650 ;
        RECT 893.970 2595.720 946.950 2596.650 ;
        RECT 947.790 2595.720 1001.230 2596.650 ;
        RECT 1002.070 2595.720 1055.510 2596.650 ;
        RECT 1056.350 2595.720 1109.790 2596.650 ;
        RECT 1110.630 2595.720 1163.610 2596.650 ;
        RECT 1164.450 2595.720 1217.890 2596.650 ;
        RECT 1218.730 2595.720 1272.170 2596.650 ;
        RECT 1273.010 2595.720 1326.450 2596.650 ;
        RECT 1327.290 2595.720 1380.270 2596.650 ;
        RECT 1381.110 2595.720 1434.550 2596.650 ;
        RECT 1435.390 2595.720 1488.830 2596.650 ;
        RECT 1489.670 2595.720 1543.110 2596.650 ;
        RECT 1543.950 2595.720 1596.930 2596.650 ;
        RECT 1597.770 2595.720 1651.210 2596.650 ;
        RECT 1652.050 2595.720 1705.490 2596.650 ;
        RECT 1706.330 2595.720 1759.770 2596.650 ;
        RECT 1760.610 2595.720 1813.590 2596.650 ;
        RECT 1814.430 2595.720 1867.870 2596.650 ;
        RECT 1868.710 2595.720 1922.150 2596.650 ;
        RECT 1922.990 2595.720 1976.430 2596.650 ;
        RECT 1977.270 2595.720 2030.250 2596.650 ;
        RECT 2031.090 2595.720 2084.530 2596.650 ;
        RECT 2085.370 2595.720 2138.810 2596.650 ;
        RECT 2139.650 2595.720 2193.090 2596.650 ;
        RECT 2193.930 2595.720 2246.910 2596.650 ;
        RECT 2247.750 2595.720 2301.190 2596.650 ;
        RECT 2302.030 2595.720 2355.470 2596.650 ;
        RECT 2356.310 2595.720 2409.750 2596.650 ;
        RECT 2410.590 2595.720 2463.570 2596.650 ;
        RECT 2464.410 2595.720 2517.850 2596.650 ;
        RECT 2518.690 2595.720 2572.130 2596.650 ;
        RECT 2572.970 2595.720 2599.360 2596.650 ;
        RECT 6.990 4.280 2599.360 2595.720 ;
        RECT 6.990 4.000 185.190 4.280 ;
        RECT 186.030 4.000 556.410 4.280 ;
        RECT 557.250 4.000 927.630 4.280 ;
        RECT 928.470 4.000 1299.310 4.280 ;
        RECT 1300.150 4.000 1670.530 4.280 ;
        RECT 1671.370 4.000 2042.210 4.280 ;
        RECT 2043.050 4.000 2413.430 4.280 ;
        RECT 2414.270 4.000 2599.360 4.280 ;
      LAYER met3 ;
        RECT 4.000 2573.480 2596.000 2586.885 ;
        RECT 4.400 2572.080 2595.600 2573.480 ;
        RECT 4.000 2519.080 2596.000 2572.080 ;
        RECT 4.400 2517.680 2595.600 2519.080 ;
        RECT 4.000 2465.360 2596.000 2517.680 ;
        RECT 4.400 2463.960 2595.600 2465.360 ;
        RECT 4.000 2410.960 2596.000 2463.960 ;
        RECT 4.400 2409.560 2595.600 2410.960 ;
        RECT 4.000 2356.560 2596.000 2409.560 ;
        RECT 4.400 2355.160 2595.600 2356.560 ;
        RECT 4.000 2302.840 2596.000 2355.160 ;
        RECT 4.400 2301.440 2595.600 2302.840 ;
        RECT 4.000 2248.440 2596.000 2301.440 ;
        RECT 4.400 2247.040 2595.600 2248.440 ;
        RECT 4.000 2194.040 2596.000 2247.040 ;
        RECT 4.400 2192.640 2595.600 2194.040 ;
        RECT 4.000 2140.320 2596.000 2192.640 ;
        RECT 4.400 2138.920 2595.600 2140.320 ;
        RECT 4.000 2085.920 2596.000 2138.920 ;
        RECT 4.400 2084.520 2595.600 2085.920 ;
        RECT 4.000 2031.520 2596.000 2084.520 ;
        RECT 4.400 2030.120 2595.600 2031.520 ;
        RECT 4.000 1977.800 2596.000 2030.120 ;
        RECT 4.400 1976.400 2595.600 1977.800 ;
        RECT 4.000 1923.400 2596.000 1976.400 ;
        RECT 4.400 1922.000 2595.600 1923.400 ;
        RECT 4.000 1869.000 2596.000 1922.000 ;
        RECT 4.400 1867.600 2595.600 1869.000 ;
        RECT 4.000 1815.280 2596.000 1867.600 ;
        RECT 4.400 1813.880 2595.600 1815.280 ;
        RECT 4.000 1760.880 2596.000 1813.880 ;
        RECT 4.400 1759.480 2595.600 1760.880 ;
        RECT 4.000 1706.480 2596.000 1759.480 ;
        RECT 4.400 1705.080 2595.600 1706.480 ;
        RECT 4.000 1652.760 2596.000 1705.080 ;
        RECT 4.400 1651.360 2595.600 1652.760 ;
        RECT 4.000 1598.360 2596.000 1651.360 ;
        RECT 4.400 1596.960 2595.600 1598.360 ;
        RECT 4.000 1543.960 2596.000 1596.960 ;
        RECT 4.400 1542.560 2595.600 1543.960 ;
        RECT 4.000 1490.240 2596.000 1542.560 ;
        RECT 4.400 1488.840 2595.600 1490.240 ;
        RECT 4.000 1435.840 2596.000 1488.840 ;
        RECT 4.400 1434.440 2595.600 1435.840 ;
        RECT 4.000 1381.440 2596.000 1434.440 ;
        RECT 4.400 1380.040 2595.600 1381.440 ;
        RECT 4.000 1327.720 2596.000 1380.040 ;
        RECT 4.400 1326.320 2595.600 1327.720 ;
        RECT 4.000 1273.320 2596.000 1326.320 ;
        RECT 4.400 1271.920 2595.600 1273.320 ;
        RECT 4.000 1218.920 2596.000 1271.920 ;
        RECT 4.400 1217.520 2595.600 1218.920 ;
        RECT 4.000 1165.200 2596.000 1217.520 ;
        RECT 4.400 1163.800 2595.600 1165.200 ;
        RECT 4.000 1110.800 2596.000 1163.800 ;
        RECT 4.400 1109.400 2595.600 1110.800 ;
        RECT 4.000 1056.400 2596.000 1109.400 ;
        RECT 4.400 1055.000 2595.600 1056.400 ;
        RECT 4.000 1002.680 2596.000 1055.000 ;
        RECT 4.400 1001.280 2595.600 1002.680 ;
        RECT 4.000 948.280 2596.000 1001.280 ;
        RECT 4.400 946.880 2595.600 948.280 ;
        RECT 4.000 893.880 2596.000 946.880 ;
        RECT 4.400 892.480 2595.600 893.880 ;
        RECT 4.000 840.160 2596.000 892.480 ;
        RECT 4.400 838.760 2595.600 840.160 ;
        RECT 4.000 785.760 2596.000 838.760 ;
        RECT 4.400 784.360 2595.600 785.760 ;
        RECT 4.000 731.360 2596.000 784.360 ;
        RECT 4.400 729.960 2595.600 731.360 ;
        RECT 4.000 677.640 2596.000 729.960 ;
        RECT 4.400 676.240 2595.600 677.640 ;
        RECT 4.000 623.240 2596.000 676.240 ;
        RECT 4.400 621.840 2595.600 623.240 ;
        RECT 4.000 568.840 2596.000 621.840 ;
        RECT 4.400 567.440 2595.600 568.840 ;
        RECT 4.000 515.120 2596.000 567.440 ;
        RECT 4.400 513.720 2595.600 515.120 ;
        RECT 4.000 460.720 2596.000 513.720 ;
        RECT 4.400 459.320 2595.600 460.720 ;
        RECT 4.000 406.320 2596.000 459.320 ;
        RECT 4.400 404.920 2595.600 406.320 ;
        RECT 4.000 352.600 2596.000 404.920 ;
        RECT 4.400 351.200 2595.600 352.600 ;
        RECT 4.000 298.200 2596.000 351.200 ;
        RECT 4.400 296.800 2595.600 298.200 ;
        RECT 4.000 243.800 2596.000 296.800 ;
        RECT 4.400 242.400 2595.600 243.800 ;
        RECT 4.000 190.080 2596.000 242.400 ;
        RECT 4.400 188.680 2595.600 190.080 ;
        RECT 4.000 135.680 2596.000 188.680 ;
        RECT 4.400 134.280 2595.600 135.680 ;
        RECT 4.000 81.280 2596.000 134.280 ;
        RECT 4.400 79.880 2595.600 81.280 ;
        RECT 4.000 27.560 2596.000 79.880 ;
        RECT 4.400 26.160 2595.600 27.560 ;
        RECT 4.000 10.715 2596.000 26.160 ;
      LAYER met4 ;
        RECT 44.455 34.175 97.440 2553.225 ;
        RECT 99.840 34.175 174.240 2553.225 ;
        RECT 176.640 34.175 251.040 2553.225 ;
        RECT 253.440 34.175 327.840 2553.225 ;
        RECT 330.240 34.175 404.640 2553.225 ;
        RECT 407.040 34.175 481.440 2553.225 ;
        RECT 483.840 34.175 558.240 2553.225 ;
        RECT 560.640 34.175 635.040 2553.225 ;
        RECT 637.440 34.175 711.840 2553.225 ;
        RECT 714.240 34.175 788.640 2553.225 ;
        RECT 791.040 34.175 865.440 2553.225 ;
        RECT 867.840 34.175 942.240 2553.225 ;
        RECT 944.640 34.175 1019.040 2553.225 ;
        RECT 1021.440 34.175 1095.840 2553.225 ;
        RECT 1098.240 34.175 1172.640 2553.225 ;
        RECT 1175.040 34.175 1249.440 2553.225 ;
        RECT 1251.840 34.175 1326.240 2553.225 ;
        RECT 1328.640 34.175 1403.040 2553.225 ;
        RECT 1405.440 34.175 1479.840 2553.225 ;
        RECT 1482.240 34.175 1556.640 2553.225 ;
        RECT 1559.040 34.175 1633.440 2553.225 ;
        RECT 1635.840 34.175 1710.240 2553.225 ;
        RECT 1712.640 34.175 1787.040 2553.225 ;
        RECT 1789.440 34.175 1863.840 2553.225 ;
        RECT 1866.240 34.175 1940.640 2553.225 ;
        RECT 1943.040 34.175 2017.440 2553.225 ;
        RECT 2019.840 34.175 2094.240 2553.225 ;
        RECT 2096.640 34.175 2171.040 2553.225 ;
        RECT 2173.440 34.175 2247.840 2553.225 ;
        RECT 2250.240 34.175 2324.640 2553.225 ;
        RECT 2327.040 34.175 2401.440 2553.225 ;
        RECT 2403.840 34.175 2478.240 2553.225 ;
        RECT 2480.640 34.175 2555.040 2553.225 ;
        RECT 2557.440 34.175 2586.745 2553.225 ;
  END
END top
END LIBRARY

