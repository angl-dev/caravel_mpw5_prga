magic
tech sky130A
magscale 1 2
timestamp 1647052296
<< locali >>
rect 22845 45883 22879 45985
rect 9781 44183 9815 44489
rect 7297 33303 7331 33541
rect 25329 32895 25363 33065
rect 19073 32215 19107 32385
rect 21373 32215 21407 32521
rect 26341 31195 26375 31433
rect 6193 28475 6227 28577
rect 17141 26775 17175 27081
rect 23029 25347 23063 25449
rect 2329 25143 2363 25245
rect 25053 24599 25087 24701
rect 8769 18139 8803 18309
rect 6193 15351 6227 15589
rect 13277 14807 13311 15045
rect 18061 14807 18095 15113
rect 3065 14331 3099 14433
rect 5641 10659 5675 10761
rect 16129 7327 16163 7497
rect 5273 7191 5307 7293
rect 19257 5151 19291 5321
rect 19073 3927 19107 4029
rect 19441 3587 19475 3689
<< viali >>
rect 1409 48161 1443 48195
rect 9137 48161 9171 48195
rect 15853 48161 15887 48195
rect 25145 48161 25179 48195
rect 31125 48161 31159 48195
rect 8953 48025 8987 48059
rect 15393 48025 15427 48059
rect 24961 48025 24995 48059
rect 1593 47957 1627 47991
rect 11713 47957 11747 47991
rect 15945 47957 15979 47991
rect 16957 47957 16991 47991
rect 18153 47957 18187 47991
rect 19533 47957 19567 47991
rect 20085 47957 20119 47991
rect 31309 47957 31343 47991
rect 1409 47753 1443 47787
rect 14197 47753 14231 47787
rect 14933 47685 14967 47719
rect 13277 47617 13311 47651
rect 8309 47549 8343 47583
rect 10517 47549 10551 47583
rect 13001 47549 13035 47583
rect 13185 47549 13219 47583
rect 13369 47549 13403 47583
rect 13553 47549 13587 47583
rect 15393 47549 15427 47583
rect 17325 47549 17359 47583
rect 21097 47549 21131 47583
rect 21833 47549 21867 47583
rect 8042 47481 8076 47515
rect 10784 47481 10818 47515
rect 15660 47481 15694 47515
rect 17592 47481 17626 47515
rect 20852 47481 20886 47515
rect 22100 47481 22134 47515
rect 6929 47413 6963 47447
rect 11897 47413 11931 47447
rect 12817 47413 12851 47447
rect 16773 47413 16807 47447
rect 18705 47413 18739 47447
rect 19717 47413 19751 47447
rect 23213 47413 23247 47447
rect 15393 47209 15427 47243
rect 22569 47209 22603 47243
rect 24777 47209 24811 47243
rect 31309 47209 31343 47243
rect 12440 47141 12474 47175
rect 23664 47141 23698 47175
rect 25237 47141 25271 47175
rect 7757 47073 7791 47107
rect 8013 47073 8047 47107
rect 9597 47073 9631 47107
rect 9864 47073 9898 47107
rect 14269 47073 14303 47107
rect 16129 47073 16163 47107
rect 17794 47073 17828 47107
rect 18061 47073 18095 47107
rect 18705 47073 18739 47107
rect 18961 47073 18995 47107
rect 21097 47073 21131 47107
rect 21833 47073 21867 47107
rect 22017 47073 22051 47107
rect 22385 47073 22419 47107
rect 31125 47073 31159 47107
rect 12173 47005 12207 47039
rect 14013 47005 14047 47039
rect 22109 47005 22143 47039
rect 22201 47005 22235 47039
rect 23397 47005 23431 47039
rect 11621 46937 11655 46971
rect 16037 46937 16071 46971
rect 20637 46937 20671 46971
rect 21189 46937 21223 46971
rect 9137 46869 9171 46903
rect 10977 46869 11011 46903
rect 13553 46869 13587 46903
rect 16681 46869 16715 46903
rect 20085 46869 20119 46903
rect 30665 46869 30699 46903
rect 8401 46665 8435 46699
rect 13553 46665 13587 46699
rect 17877 46665 17911 46699
rect 18337 46665 18371 46699
rect 8033 46529 8067 46563
rect 9505 46529 9539 46563
rect 22477 46529 22511 46563
rect 24679 46529 24713 46563
rect 7665 46461 7699 46495
rect 7849 46461 7883 46495
rect 7941 46461 7975 46495
rect 8217 46461 8251 46495
rect 9137 46461 9171 46495
rect 9321 46461 9355 46495
rect 9413 46461 9447 46495
rect 9689 46461 9723 46495
rect 10333 46461 10367 46495
rect 12173 46461 12207 46495
rect 14381 46461 14415 46495
rect 16221 46461 16255 46495
rect 17141 46461 17175 46495
rect 17325 46461 17359 46495
rect 17417 46461 17451 46495
rect 17509 46461 17543 46495
rect 17693 46461 17727 46495
rect 24409 46461 24443 46495
rect 24593 46461 24627 46495
rect 24777 46461 24811 46495
rect 24961 46461 24995 46495
rect 25605 46461 25639 46495
rect 9873 46393 9907 46427
rect 10578 46393 10612 46427
rect 12440 46393 12474 46427
rect 14648 46393 14682 46427
rect 20269 46393 20303 46427
rect 22722 46393 22756 46427
rect 11713 46325 11747 46359
rect 15761 46325 15795 46359
rect 16313 46325 16347 46359
rect 19809 46325 19843 46359
rect 21557 46325 21591 46359
rect 23857 46325 23891 46359
rect 25145 46325 25179 46359
rect 25697 46325 25731 46359
rect 9781 46121 9815 46155
rect 10977 46121 11011 46155
rect 13369 46121 13403 46155
rect 14565 46121 14599 46155
rect 15761 46121 15795 46155
rect 17417 46121 17451 46155
rect 18797 46121 18831 46155
rect 20729 46121 20763 46155
rect 23204 46053 23238 46087
rect 1397 45985 1431 46019
rect 6377 45985 6411 46019
rect 6644 45985 6678 46019
rect 8401 45985 8435 46019
rect 9045 45985 9079 46019
rect 9229 45985 9263 46019
rect 9413 45985 9447 46019
rect 9597 45985 9631 46019
rect 10241 45985 10275 46019
rect 10425 45985 10459 46019
rect 10793 45985 10827 46019
rect 11689 45985 11723 46019
rect 12633 45985 12667 46019
rect 12817 45985 12851 46019
rect 13185 45985 13219 46019
rect 13829 45985 13863 46019
rect 14013 45985 14047 46019
rect 14381 45985 14415 46019
rect 15025 45985 15059 46019
rect 15209 45985 15243 46019
rect 15577 45985 15611 46019
rect 16681 45985 16715 46019
rect 16865 45985 16899 46019
rect 16957 45985 16991 46019
rect 17233 45985 17267 46019
rect 17877 45985 17911 46019
rect 18981 45985 19015 46019
rect 19349 45985 19383 46019
rect 19533 45985 19567 46019
rect 19993 45985 20027 46019
rect 20177 45985 20211 46019
rect 20269 45985 20303 46019
rect 20545 45985 20579 46019
rect 21189 45985 21223 46019
rect 22017 45985 22051 46019
rect 22109 45985 22143 46019
rect 22385 45985 22419 46019
rect 22845 45985 22879 46019
rect 25890 45985 25924 46019
rect 30665 45985 30699 46019
rect 31125 45985 31159 46019
rect 9321 45917 9355 45951
rect 10517 45917 10551 45951
rect 10609 45917 10643 45951
rect 12909 45917 12943 45951
rect 13001 45917 13035 45951
rect 14105 45917 14139 45951
rect 14197 45917 14231 45951
rect 15301 45917 15335 45951
rect 15393 45917 15427 45951
rect 17049 45917 17083 45951
rect 19165 45917 19199 45951
rect 19257 45917 19291 45951
rect 20361 45917 20395 45951
rect 22937 45917 22971 45951
rect 26157 45917 26191 45951
rect 7757 45849 7791 45883
rect 22293 45849 22327 45883
rect 22845 45849 22879 45883
rect 31309 45849 31343 45883
rect 1593 45781 1627 45815
rect 8493 45781 8527 45815
rect 11621 45781 11655 45815
rect 17969 45781 18003 45815
rect 21833 45781 21867 45815
rect 24317 45781 24351 45815
rect 24777 45781 24811 45815
rect 1409 45577 1443 45611
rect 9413 45577 9447 45611
rect 26249 45577 26283 45611
rect 8033 45509 8067 45543
rect 16405 45509 16439 45543
rect 21097 45509 21131 45543
rect 22385 45509 22419 45543
rect 7573 45441 7607 45475
rect 12817 45441 12851 45475
rect 14105 45441 14139 45475
rect 14473 45441 14507 45475
rect 14565 45441 14599 45475
rect 23397 45441 23431 45475
rect 24409 45441 24443 45475
rect 6837 45373 6871 45407
rect 7297 45373 7331 45407
rect 7485 45373 7519 45407
rect 7665 45373 7699 45407
rect 7849 45373 7883 45407
rect 10057 45373 10091 45407
rect 10885 45373 10919 45407
rect 11437 45373 11471 45407
rect 12081 45373 12115 45407
rect 12541 45373 12575 45407
rect 14289 45373 14323 45407
rect 14657 45373 14691 45407
rect 14841 45373 14875 45407
rect 15301 45373 15335 45407
rect 16129 45373 16163 45407
rect 16221 45373 16255 45407
rect 16497 45373 16531 45407
rect 17325 45373 17359 45407
rect 20637 45373 20671 45407
rect 21281 45373 21315 45407
rect 21465 45373 21499 45407
rect 21557 45373 21591 45407
rect 21649 45373 21683 45407
rect 21833 45373 21867 45407
rect 22293 45373 22327 45407
rect 23121 45373 23155 45407
rect 23305 45375 23339 45409
rect 23489 45373 23523 45407
rect 23673 45373 23707 45407
rect 26801 45373 26835 45407
rect 9505 45305 9539 45339
rect 17592 45305 17626 45339
rect 20392 45305 20426 45339
rect 23857 45305 23891 45339
rect 24654 45305 24688 45339
rect 6745 45237 6779 45271
rect 10149 45237 10183 45271
rect 10793 45237 10827 45271
rect 11989 45237 12023 45271
rect 15393 45237 15427 45271
rect 15945 45237 15979 45271
rect 18705 45237 18739 45271
rect 19257 45237 19291 45271
rect 25789 45237 25823 45271
rect 7205 45033 7239 45067
rect 17969 45033 18003 45067
rect 18521 45033 18555 45067
rect 22569 45033 22603 45067
rect 24133 45033 24167 45067
rect 12265 44965 12299 44999
rect 7389 44897 7423 44931
rect 7757 44897 7791 44931
rect 7941 44897 7975 44931
rect 10241 44897 10275 44931
rect 10425 44897 10459 44931
rect 10793 44897 10827 44931
rect 11713 44897 11747 44931
rect 12173 44897 12207 44931
rect 13553 44897 13587 44931
rect 14657 44897 14691 44931
rect 14749 44897 14783 44931
rect 15025 44897 15059 44931
rect 15485 44897 15519 44931
rect 15669 44897 15703 44931
rect 15761 44897 15795 44931
rect 16037 44897 16071 44931
rect 17233 44897 17267 44931
rect 17417 44897 17451 44931
rect 17785 44897 17819 44931
rect 18613 44897 18647 44931
rect 19073 44897 19107 44931
rect 19809 44897 19843 44931
rect 21005 44897 21039 44931
rect 21833 44897 21867 44931
rect 22017 44897 22051 44931
rect 22201 44897 22235 44931
rect 22385 44897 22419 44931
rect 23397 44897 23431 44931
rect 23569 44895 23603 44929
rect 23667 44897 23701 44931
rect 23949 44897 23983 44931
rect 24593 44897 24627 44931
rect 24869 44897 24903 44931
rect 24961 44897 24995 44931
rect 28098 44897 28132 44931
rect 7573 44829 7607 44863
rect 7665 44829 7699 44863
rect 9137 44829 9171 44863
rect 9413 44829 9447 44863
rect 10517 44829 10551 44863
rect 10609 44829 10643 44863
rect 13829 44829 13863 44863
rect 17509 44829 17543 44863
rect 17601 44829 17635 44863
rect 21281 44829 21315 44863
rect 22109 44829 22143 44863
rect 23765 44829 23799 44863
rect 26157 44829 26191 44863
rect 28365 44829 28399 44863
rect 10977 44761 11011 44795
rect 14473 44761 14507 44795
rect 19165 44761 19199 44795
rect 25605 44761 25639 44795
rect 11621 44693 11655 44727
rect 14933 44693 14967 44727
rect 15945 44693 15979 44727
rect 16773 44693 16807 44727
rect 19901 44693 19935 44727
rect 24685 44693 24719 44727
rect 25145 44693 25179 44727
rect 26985 44693 27019 44727
rect 30941 44693 30975 44727
rect 9781 44489 9815 44523
rect 27997 44489 28031 44523
rect 7205 44421 7239 44455
rect 8309 44353 8343 44387
rect 5825 44285 5859 44319
rect 8033 44285 8067 44319
rect 8125 44285 8159 44319
rect 8401 44285 8435 44319
rect 1869 44217 1903 44251
rect 6092 44217 6126 44251
rect 24501 44421 24535 44455
rect 28549 44421 28583 44455
rect 14105 44353 14139 44387
rect 14381 44353 14415 44387
rect 15853 44353 15887 44387
rect 20729 44353 20763 44387
rect 21005 44353 21039 44387
rect 22661 44353 22695 44387
rect 12081 44285 12115 44319
rect 12348 44285 12382 44319
rect 15485 44285 15519 44319
rect 15669 44285 15703 44319
rect 15761 44285 15795 44319
rect 16037 44285 16071 44319
rect 16865 44285 16899 44319
rect 17049 44285 17083 44319
rect 17141 44285 17175 44319
rect 17233 44285 17267 44319
rect 17417 44285 17451 44319
rect 18245 44285 18279 44319
rect 19257 44285 19291 44319
rect 21465 44285 21499 44319
rect 22477 44285 22511 44319
rect 22753 44285 22787 44319
rect 22845 44285 22879 44319
rect 23029 44285 23063 44319
rect 23673 44285 23707 44319
rect 24409 44285 24443 44319
rect 26985 44285 27019 44319
rect 31125 44285 31159 44319
rect 9873 44217 9907 44251
rect 11621 44217 11655 44251
rect 18153 44217 18187 44251
rect 26718 44217 26752 44251
rect 2145 44149 2179 44183
rect 7849 44149 7883 44183
rect 9229 44149 9263 44183
rect 9781 44149 9815 44183
rect 13461 44149 13495 44183
rect 16221 44149 16255 44183
rect 17601 44149 17635 44183
rect 19349 44149 19383 44183
rect 21557 44149 21591 44183
rect 22293 44149 22327 44183
rect 23581 44149 23615 44183
rect 25145 44149 25179 44183
rect 25605 44149 25639 44183
rect 27445 44149 27479 44183
rect 30665 44149 30699 44183
rect 31309 44149 31343 44183
rect 6837 43945 6871 43979
rect 11805 43945 11839 43979
rect 18613 43945 18647 43979
rect 24593 43945 24627 43979
rect 26433 43945 26467 43979
rect 29377 43945 29411 43979
rect 1593 43877 1627 43911
rect 17500 43877 17534 43911
rect 7021 43809 7055 43843
rect 7389 43809 7423 43843
rect 7573 43809 7607 43843
rect 8861 43809 8895 43843
rect 10885 43809 10919 43843
rect 11897 43809 11931 43843
rect 12624 43809 12658 43843
rect 14197 43809 14231 43843
rect 14381 43809 14415 43843
rect 14749 43809 14783 43843
rect 14933 43809 14967 43843
rect 15577 43809 15611 43843
rect 15853 43809 15887 43843
rect 15945 43809 15979 43843
rect 16129 43809 16163 43843
rect 16773 43809 16807 43843
rect 19349 43809 19383 43843
rect 20361 43809 20395 43843
rect 20545 43809 20579 43843
rect 20729 43809 20763 43843
rect 20913 43809 20947 43843
rect 22017 43809 22051 43843
rect 22385 43809 22419 43843
rect 22569 43809 22603 43843
rect 23489 43809 23523 43843
rect 24685 43809 24719 43843
rect 25697 43809 25731 43843
rect 25881 43809 25915 43843
rect 26249 43809 26283 43843
rect 27701 43809 27735 43843
rect 7205 43741 7239 43775
rect 7297 43741 7331 43775
rect 8585 43741 8619 43775
rect 9321 43741 9355 43775
rect 9597 43741 9631 43775
rect 12357 43741 12391 43775
rect 14565 43741 14599 43775
rect 14657 43741 14691 43775
rect 15761 43741 15795 43775
rect 17233 43741 17267 43775
rect 19073 43741 19107 43775
rect 20637 43741 20671 43775
rect 22201 43741 22235 43775
rect 22293 43741 22327 43775
rect 23213 43741 23247 43775
rect 25973 43741 26007 43775
rect 26065 43741 26099 43775
rect 27445 43741 27479 43775
rect 13737 43673 13771 43707
rect 2145 43605 2179 43639
rect 5825 43605 5859 43639
rect 10793 43605 10827 43639
rect 15393 43605 15427 43639
rect 21097 43605 21131 43639
rect 21833 43605 21867 43639
rect 25237 43605 25271 43639
rect 28825 43605 28859 43639
rect 30481 43605 30515 43639
rect 31033 43605 31067 43639
rect 23857 43401 23891 43435
rect 27169 43401 27203 43435
rect 30665 43401 30699 43435
rect 31309 43401 31343 43435
rect 6009 43265 6043 43299
rect 10977 43265 11011 43299
rect 12449 43265 12483 43299
rect 12725 43265 12759 43299
rect 16589 43265 16623 43299
rect 18429 43265 18463 43299
rect 20913 43265 20947 43299
rect 22477 43265 22511 43299
rect 22753 43265 22787 43299
rect 26801 43265 26835 43299
rect 8217 43197 8251 43231
rect 9413 43197 9447 43231
rect 9689 43197 9723 43231
rect 10701 43197 10735 43231
rect 10885 43197 10919 43231
rect 11069 43197 11103 43231
rect 11253 43197 11287 43231
rect 15485 43197 15519 43231
rect 16313 43197 16347 43231
rect 18705 43197 18739 43231
rect 19533 43197 19567 43231
rect 20637 43197 20671 43231
rect 21465 43197 21499 43231
rect 24409 43197 24443 43231
rect 26433 43197 26467 43231
rect 26617 43197 26651 43231
rect 26709 43197 26743 43231
rect 26985 43197 27019 43231
rect 27629 43197 27663 43231
rect 31125 43197 31159 43231
rect 6276 43129 6310 43163
rect 11897 43129 11931 43163
rect 15240 43129 15274 43163
rect 24654 43129 24688 43163
rect 27896 43129 27930 43163
rect 1501 43061 1535 43095
rect 1961 43061 1995 43095
rect 2605 43061 2639 43095
rect 3065 43061 3099 43095
rect 4905 43061 4939 43095
rect 5549 43061 5583 43095
rect 7389 43061 7423 43095
rect 8309 43061 8343 43095
rect 11437 43061 11471 43095
rect 14105 43061 14139 43095
rect 19441 43061 19475 43095
rect 21557 43061 21591 43095
rect 25789 43061 25823 43095
rect 29009 43061 29043 43095
rect 29561 43061 29595 43095
rect 15393 42857 15427 42891
rect 28273 42857 28307 42891
rect 11796 42789 11830 42823
rect 5733 42721 5767 42755
rect 7297 42721 7331 42755
rect 8217 42721 8251 42755
rect 9229 42721 9263 42755
rect 9413 42721 9447 42755
rect 9505 42721 9539 42755
rect 9781 42721 9815 42755
rect 10609 42721 10643 42755
rect 10701 42721 10735 42755
rect 10977 42721 11011 42755
rect 11529 42721 11563 42755
rect 13645 42721 13679 42755
rect 14657 42721 14691 42755
rect 14841 42721 14875 42755
rect 15209 42721 15243 42755
rect 15853 42721 15887 42755
rect 16957 42721 16991 42755
rect 17141 42721 17175 42755
rect 17509 42721 17543 42755
rect 18613 42721 18647 42755
rect 18880 42721 18914 42755
rect 20453 42721 20487 42755
rect 22385 42721 22419 42755
rect 22569 42721 22603 42755
rect 22753 42721 22787 42755
rect 22845 42721 22879 42755
rect 22937 42721 22971 42755
rect 23121 42721 23155 42755
rect 23569 42731 23603 42765
rect 23765 42721 23799 42755
rect 23857 42721 23891 42755
rect 24133 42721 24167 42755
rect 26249 42721 26283 42755
rect 27537 42721 27571 42755
rect 27721 42721 27755 42755
rect 28089 42721 28123 42755
rect 28733 42721 28767 42755
rect 29377 42721 29411 42755
rect 30941 42721 30975 42755
rect 4537 42653 4571 42687
rect 6837 42653 6871 42687
rect 7941 42653 7975 42687
rect 9597 42653 9631 42687
rect 13369 42653 13403 42687
rect 14933 42653 14967 42687
rect 15025 42653 15059 42687
rect 17233 42653 17267 42687
rect 17325 42653 17359 42687
rect 20729 42653 20763 42687
rect 23949 42653 23983 42687
rect 24961 42653 24995 42687
rect 25237 42653 25271 42687
rect 27813 42653 27847 42687
rect 27905 42653 27939 42687
rect 15945 42585 15979 42619
rect 29469 42585 29503 42619
rect 1501 42517 1535 42551
rect 2053 42517 2087 42551
rect 2513 42517 2547 42551
rect 3065 42517 3099 42551
rect 3985 42517 4019 42551
rect 5181 42517 5215 42551
rect 7389 42517 7423 42551
rect 9965 42517 9999 42551
rect 10425 42517 10459 42551
rect 10885 42517 10919 42551
rect 12909 42517 12943 42551
rect 17693 42517 17727 42551
rect 19993 42517 20027 42551
rect 21833 42517 21867 42551
rect 24317 42517 24351 42551
rect 26341 42517 26375 42551
rect 26985 42517 27019 42551
rect 28825 42517 28859 42551
rect 30113 42517 30147 42551
rect 4997 42313 5031 42347
rect 7297 42313 7331 42347
rect 11621 42313 11655 42347
rect 21281 42313 21315 42347
rect 22937 42313 22971 42347
rect 26985 42313 27019 42347
rect 3249 42245 3283 42279
rect 13461 42245 13495 42279
rect 23397 42245 23431 42279
rect 3893 42177 3927 42211
rect 7748 42177 7782 42211
rect 9321 42177 9355 42211
rect 10419 42177 10453 42211
rect 12173 42177 12207 42211
rect 14473 42177 14507 42211
rect 16304 42177 16338 42211
rect 18429 42177 18463 42211
rect 22017 42177 22051 42211
rect 22109 42177 22143 42211
rect 29837 42177 29871 42211
rect 29929 42177 29963 42211
rect 1869 42109 1903 42143
rect 2237 42109 2271 42143
rect 6653 42109 6687 42143
rect 7481 42109 7515 42143
rect 7665 42109 7699 42143
rect 7849 42107 7883 42141
rect 8033 42109 8067 42143
rect 8953 42109 8987 42143
rect 9137 42109 9171 42143
rect 9229 42109 9263 42143
rect 9505 42109 9539 42143
rect 10149 42109 10183 42143
rect 10333 42111 10367 42145
rect 10517 42109 10551 42143
rect 10701 42109 10735 42143
rect 11529 42109 11563 42143
rect 12449 42109 12483 42143
rect 14289 42109 14323 42143
rect 14565 42109 14599 42143
rect 14657 42109 14691 42143
rect 14841 42109 14875 42143
rect 16037 42109 16071 42143
rect 16221 42109 16255 42143
rect 16405 42111 16439 42145
rect 16589 42109 16623 42143
rect 18162 42109 18196 42143
rect 19257 42109 19291 42143
rect 19901 42109 19935 42143
rect 21741 42109 21775 42143
rect 21925 42109 21959 42143
rect 22304 42109 22338 42143
rect 23121 42109 23155 42143
rect 23213 42109 23247 42143
rect 23489 42109 23523 42143
rect 24409 42109 24443 42143
rect 26249 42099 26283 42133
rect 26437 42111 26471 42145
rect 26525 42109 26559 42143
rect 26663 42109 26697 42143
rect 26801 42109 26835 42143
rect 27445 42109 27479 42143
rect 28273 42109 28307 42143
rect 29009 42109 29043 42143
rect 29561 42109 29595 42143
rect 29745 42109 29779 42143
rect 30113 42109 30147 42143
rect 31125 42109 31159 42143
rect 5641 42041 5675 42075
rect 20168 42041 20202 42075
rect 24654 42041 24688 42075
rect 28181 42041 28215 42075
rect 4445 41973 4479 42007
rect 6101 41973 6135 42007
rect 6745 41973 6779 42007
rect 9689 41973 9723 42007
rect 10885 41973 10919 42007
rect 14105 41973 14139 42007
rect 15393 41973 15427 42007
rect 15853 41973 15887 42007
rect 17049 41973 17083 42007
rect 19349 41973 19383 42007
rect 22477 41973 22511 42007
rect 25789 41973 25823 42007
rect 27537 41973 27571 42007
rect 28917 41973 28951 42007
rect 30297 41973 30331 42007
rect 31309 41973 31343 42007
rect 2697 41769 2731 41803
rect 9413 41769 9447 41803
rect 17877 41769 17911 41803
rect 23949 41769 23983 41803
rect 30021 41769 30055 41803
rect 31033 41769 31067 41803
rect 2145 41701 2179 41735
rect 7512 41701 7546 41735
rect 8217 41701 8251 41735
rect 14197 41701 14231 41735
rect 22201 41701 22235 41735
rect 28908 41701 28942 41735
rect 3709 41633 3743 41667
rect 3976 41633 4010 41667
rect 8401 41633 8435 41667
rect 8585 41633 8619 41667
rect 8769 41633 8803 41667
rect 8953 41633 8987 41667
rect 9597 41633 9631 41667
rect 9689 41633 9723 41667
rect 9965 41633 9999 41667
rect 10793 41633 10827 41667
rect 12081 41633 12115 41667
rect 13093 41633 13127 41667
rect 13369 41633 13403 41667
rect 16681 41633 16715 41667
rect 16865 41633 16899 41667
rect 16957 41633 16991 41667
rect 17233 41633 17267 41667
rect 18981 41633 19015 41667
rect 20269 41633 20303 41667
rect 21005 41633 21039 41667
rect 21833 41633 21867 41667
rect 22017 41633 22051 41667
rect 23213 41633 23247 41667
rect 23397 41633 23431 41667
rect 23857 41633 23891 41667
rect 25053 41633 25087 41667
rect 25320 41633 25354 41667
rect 27077 41633 27111 41667
rect 28181 41633 28215 41667
rect 5733 41565 5767 41599
rect 7757 41565 7791 41599
rect 8677 41565 8711 41599
rect 10701 41565 10735 41599
rect 17049 41565 17083 41599
rect 19257 41565 19291 41599
rect 20545 41565 20579 41599
rect 28641 41565 28675 41599
rect 6377 41497 6411 41531
rect 11989 41497 12023 41531
rect 1593 41429 1627 41463
rect 3249 41429 3283 41463
rect 5089 41429 5123 41463
rect 9873 41429 9907 41463
rect 10425 41429 10459 41463
rect 10793 41429 10827 41463
rect 15485 41429 15519 41463
rect 17417 41429 17451 41463
rect 21097 41429 21131 41463
rect 23029 41429 23063 41463
rect 24593 41429 24627 41463
rect 26433 41429 26467 41463
rect 27169 41429 27203 41463
rect 28089 41429 28123 41463
rect 30481 41429 30515 41463
rect 2053 41225 2087 41259
rect 4077 41225 4111 41259
rect 8309 41225 8343 41259
rect 13093 41225 13127 41259
rect 16313 41225 16347 41259
rect 16957 41225 16991 41259
rect 18613 41225 18647 41259
rect 19257 41225 19291 41259
rect 22569 41225 22603 41259
rect 23305 41225 23339 41259
rect 25789 41225 25823 41259
rect 10517 41157 10551 41191
rect 14105 41157 14139 41191
rect 17785 41157 17819 41191
rect 11713 41089 11747 41123
rect 19708 41089 19742 41123
rect 20821 41089 20855 41123
rect 23213 41089 23247 41123
rect 26157 41089 26191 41123
rect 28641 41089 28675 41123
rect 29653 41089 29687 41123
rect 3893 41021 3927 41055
rect 4077 41021 4111 41055
rect 4537 41021 4571 41055
rect 4721 41021 4755 41055
rect 4813 41021 4847 41055
rect 4905 41021 4939 41055
rect 5641 41021 5675 41055
rect 5825 41021 5859 41055
rect 8217 41021 8251 41055
rect 8953 41021 8987 41055
rect 9229 41021 9263 41055
rect 10241 41021 10275 41055
rect 10425 41021 10459 41055
rect 10609 41021 10643 41055
rect 10701 41021 10735 41055
rect 15485 41021 15519 41055
rect 15945 41021 15979 41055
rect 16313 41021 16347 41055
rect 17141 41021 17175 41055
rect 19441 41021 19475 41055
rect 19625 41021 19659 41055
rect 19809 41021 19843 41055
rect 19993 41021 20027 41055
rect 21097 41021 21131 41055
rect 22385 41021 22419 41055
rect 22661 41021 22695 41055
rect 23121 41021 23155 41055
rect 24409 41021 24443 41055
rect 24685 41021 24719 41055
rect 25973 41021 26007 41055
rect 26249 41021 26283 41055
rect 26341 41021 26375 41055
rect 26525 41021 26559 41055
rect 26985 41021 27019 41055
rect 29920 41021 29954 41055
rect 1501 40953 1535 40987
rect 5181 40953 5215 40987
rect 7757 40953 7791 40987
rect 11980 40953 12014 40987
rect 15218 40953 15252 40987
rect 17325 40953 17359 40987
rect 17969 40953 18003 40987
rect 18153 40953 18187 40987
rect 2513 40885 2547 40919
rect 3249 40885 3283 40919
rect 5733 40885 5767 40919
rect 6653 40885 6687 40919
rect 7113 40885 7147 40919
rect 10885 40885 10919 40919
rect 16497 40885 16531 40919
rect 22109 40885 22143 40919
rect 23489 40885 23523 40919
rect 31033 40885 31067 40919
rect 4077 40681 4111 40715
rect 7849 40681 7883 40715
rect 10793 40681 10827 40715
rect 12265 40681 12299 40715
rect 14841 40681 14875 40715
rect 20729 40681 20763 40715
rect 26341 40681 26375 40715
rect 13728 40613 13762 40647
rect 15945 40613 15979 40647
rect 16129 40613 16163 40647
rect 19594 40613 19628 40647
rect 21833 40613 21867 40647
rect 1869 40545 1903 40579
rect 2964 40545 2998 40579
rect 4537 40545 4571 40579
rect 4721 40545 4755 40579
rect 4813 40545 4847 40579
rect 4951 40545 4985 40579
rect 5825 40545 5859 40579
rect 6469 40545 6503 40579
rect 6736 40545 6770 40579
rect 8493 40545 8527 40579
rect 8769 40545 8803 40579
rect 8861 40545 8895 40579
rect 9045 40545 9079 40579
rect 9505 40545 9539 40579
rect 9689 40545 9723 40579
rect 10149 40545 10183 40579
rect 10609 40545 10643 40579
rect 11713 40545 11747 40579
rect 12449 40545 12483 40579
rect 12817 40545 12851 40579
rect 13001 40545 13035 40579
rect 16865 40545 16899 40579
rect 17049 40545 17083 40579
rect 17233 40545 17267 40579
rect 17417 40545 17451 40579
rect 19349 40545 19383 40579
rect 22017 40545 22051 40579
rect 22201 40545 22235 40579
rect 22293 40545 22327 40579
rect 22477 40545 22511 40579
rect 24326 40545 24360 40579
rect 25053 40545 25087 40579
rect 25237 40545 25271 40579
rect 25605 40545 25639 40579
rect 26249 40545 26283 40579
rect 27169 40545 27203 40579
rect 27261 40545 27295 40579
rect 27537 40545 27571 40579
rect 29561 40545 29595 40579
rect 29828 40545 29862 40579
rect 2697 40477 2731 40511
rect 8309 40477 8343 40511
rect 8677 40477 8711 40511
rect 10333 40477 10367 40511
rect 10425 40477 10459 40511
rect 12633 40477 12667 40511
rect 12725 40477 12759 40511
rect 13461 40477 13495 40511
rect 17141 40477 17175 40511
rect 18613 40477 18647 40511
rect 18889 40477 18923 40511
rect 22109 40477 22143 40511
rect 24593 40477 24627 40511
rect 25329 40477 25363 40511
rect 25421 40477 25455 40511
rect 28181 40477 28215 40511
rect 28457 40477 28491 40511
rect 10517 40409 10551 40443
rect 11621 40409 11655 40443
rect 26985 40409 27019 40443
rect 1961 40341 1995 40375
rect 5181 40341 5215 40375
rect 5733 40341 5767 40375
rect 9689 40341 9723 40375
rect 15761 40341 15795 40375
rect 17601 40341 17635 40375
rect 21189 40341 21223 40375
rect 23213 40341 23247 40375
rect 25789 40341 25823 40375
rect 27445 40341 27479 40375
rect 30941 40341 30975 40375
rect 3157 40137 3191 40171
rect 9965 40137 9999 40171
rect 15761 40137 15795 40171
rect 16865 40137 16899 40171
rect 23121 40137 23155 40171
rect 30297 40137 30331 40171
rect 10425 40069 10459 40103
rect 2145 40001 2179 40035
rect 4077 40001 4111 40035
rect 4537 40001 4571 40035
rect 5457 40001 5491 40035
rect 12449 40001 12483 40035
rect 14105 40001 14139 40035
rect 22109 40001 22143 40035
rect 23489 40001 23523 40035
rect 27629 40001 27663 40035
rect 27905 40001 27939 40035
rect 1869 39933 1903 39967
rect 2053 39933 2087 39967
rect 2237 39933 2271 39967
rect 2421 39933 2455 39967
rect 3249 39933 3283 39967
rect 3801 39933 3835 39967
rect 3985 39933 4019 39967
rect 4169 39933 4203 39967
rect 4353 39933 4387 39967
rect 5549 39933 5583 39967
rect 7205 39933 7239 39967
rect 8217 39933 8251 39967
rect 9229 39933 9263 39967
rect 9413 39933 9447 39967
rect 9499 39933 9533 39967
rect 9597 39933 9631 39967
rect 9781 39933 9815 39967
rect 10793 39933 10827 39967
rect 11345 39933 11379 39967
rect 11437 39933 11471 39967
rect 12725 39933 12759 39967
rect 13277 39933 13311 39967
rect 14289 39933 14323 39967
rect 14473 39933 14507 39967
rect 14562 39933 14596 39967
rect 14657 39933 14691 39967
rect 14841 39933 14875 39967
rect 15945 39933 15979 39967
rect 17978 39933 18012 39967
rect 18245 39933 18279 39967
rect 21833 39933 21867 39967
rect 22017 39933 22051 39967
rect 22201 39933 22235 39967
rect 22385 39933 22419 39967
rect 23305 39933 23339 39967
rect 23581 39933 23615 39967
rect 23673 39933 23707 39967
rect 23857 39933 23891 39967
rect 24409 39933 24443 39967
rect 24593 39933 24627 39967
rect 25053 39933 25087 39967
rect 25320 39933 25354 39967
rect 28549 39933 28583 39967
rect 29561 39933 29595 39967
rect 29745 39933 29779 39967
rect 29837 39933 29871 39967
rect 29929 39933 29963 39967
rect 30113 39933 30147 39967
rect 31125 39933 31159 39967
rect 6653 39865 6687 39899
rect 10609 39865 10643 39899
rect 16129 39865 16163 39899
rect 19625 39865 19659 39899
rect 1685 39797 1719 39831
rect 5641 39797 5675 39831
rect 6009 39797 6043 39831
rect 6561 39797 6595 39831
rect 7297 39797 7331 39831
rect 8309 39797 8343 39831
rect 13369 39797 13403 39831
rect 20913 39797 20947 39831
rect 22569 39797 22603 39831
rect 24409 39797 24443 39831
rect 26433 39797 26467 39831
rect 28457 39797 28491 39831
rect 31309 39797 31343 39831
rect 3249 39593 3283 39627
rect 10149 39593 10183 39627
rect 14473 39593 14507 39627
rect 22109 39593 22143 39627
rect 24317 39593 24351 39627
rect 29009 39593 29043 39627
rect 23397 39525 23431 39559
rect 23581 39525 23615 39559
rect 26157 39525 26191 39559
rect 29653 39525 29687 39559
rect 29837 39525 29871 39559
rect 30849 39525 30883 39559
rect 1409 39457 1443 39491
rect 1676 39457 1710 39491
rect 3433 39457 3467 39491
rect 3801 39457 3835 39491
rect 3985 39457 4019 39491
rect 4997 39457 5031 39491
rect 5365 39457 5399 39491
rect 5641 39457 5675 39491
rect 6745 39457 6779 39491
rect 7021 39457 7055 39491
rect 7481 39457 7515 39491
rect 8309 39457 8343 39491
rect 8565 39457 8599 39491
rect 10333 39457 10367 39491
rect 10517 39457 10551 39491
rect 11805 39457 11839 39491
rect 14381 39457 14415 39491
rect 15669 39457 15703 39491
rect 15853 39457 15887 39491
rect 18254 39457 18288 39491
rect 20554 39457 20588 39491
rect 22293 39457 22327 39491
rect 22569 39457 22603 39491
rect 22753 39457 22787 39491
rect 24225 39457 24259 39491
rect 25421 39457 25455 39491
rect 25697 39457 25731 39491
rect 26341 39457 26375 39491
rect 27169 39457 27203 39491
rect 27537 39457 27571 39491
rect 27721 39457 27755 39491
rect 28273 39457 28307 39491
rect 28457 39457 28491 39491
rect 28549 39457 28583 39491
rect 28825 39457 28859 39491
rect 3617 39389 3651 39423
rect 3709 39389 3743 39423
rect 5181 39389 5215 39423
rect 5825 39389 5859 39423
rect 7205 39389 7239 39423
rect 12081 39389 12115 39423
rect 13645 39389 13679 39423
rect 13921 39389 13955 39423
rect 18521 39389 18555 39423
rect 20821 39389 20855 39423
rect 22477 39389 22511 39423
rect 27353 39389 27387 39423
rect 27445 39389 27479 39423
rect 28641 39389 28675 39423
rect 7849 39321 7883 39355
rect 22385 39321 22419 39355
rect 2789 39253 2823 39287
rect 4445 39253 4479 39287
rect 9689 39253 9723 39287
rect 15485 39253 15519 39287
rect 15669 39253 15703 39287
rect 17141 39253 17175 39287
rect 19441 39253 19475 39287
rect 26985 39253 27019 39287
rect 29469 39253 29503 39287
rect 30389 39253 30423 39287
rect 5825 39049 5859 39083
rect 6745 39049 6779 39083
rect 6929 39049 6963 39083
rect 8401 39049 8435 39083
rect 9045 39049 9079 39083
rect 14473 39049 14507 39083
rect 17969 39049 18003 39083
rect 20545 39049 20579 39083
rect 22293 39049 22327 39083
rect 26709 39049 26743 39083
rect 27169 39049 27203 39083
rect 29745 39049 29779 39083
rect 31309 39049 31343 39083
rect 9873 38981 9907 39015
rect 15301 38981 15335 39015
rect 28917 38981 28951 39015
rect 1409 38913 1443 38947
rect 7941 38913 7975 38947
rect 12357 38913 12391 38947
rect 13277 38913 13311 38947
rect 16497 38913 16531 38947
rect 16773 38913 16807 38947
rect 18429 38913 18463 38947
rect 20913 38913 20947 38947
rect 21005 38913 21039 38947
rect 23397 38913 23431 38947
rect 23489 38913 23523 38947
rect 25053 38913 25087 38947
rect 28089 38913 28123 38947
rect 3801 38845 3835 38879
rect 4537 38845 4571 38879
rect 7665 38845 7699 38879
rect 7849 38845 7883 38879
rect 8033 38845 8067 38879
rect 8217 38845 8251 38879
rect 9229 38845 9263 38879
rect 10057 38845 10091 38879
rect 13001 38845 13035 38879
rect 13185 38845 13219 38879
rect 13369 38845 13403 38879
rect 13553 38845 13587 38879
rect 14565 38845 14599 38879
rect 15025 38845 15059 38879
rect 15209 38845 15243 38879
rect 15393 38845 15427 38879
rect 15485 38845 15519 38879
rect 18153 38845 18187 38879
rect 18337 38845 18371 38879
rect 18521 38845 18555 38879
rect 18705 38845 18739 38879
rect 19809 38845 19843 38879
rect 20085 38845 20119 38879
rect 20729 38845 20763 38879
rect 21097 38845 21131 38879
rect 21281 38845 21315 38879
rect 22385 38845 22419 38879
rect 23121 38845 23155 38879
rect 23305 38845 23339 38879
rect 23673 38845 23707 38879
rect 25973 38845 26007 38879
rect 26617 38845 26651 38879
rect 26985 38845 27019 38879
rect 27721 38845 27755 38879
rect 27905 38845 27939 38879
rect 27997 38845 28031 38879
rect 28273 38845 28307 38879
rect 30481 38845 30515 38879
rect 31125 38845 31159 38879
rect 1676 38777 1710 38811
rect 6897 38777 6931 38811
rect 7113 38777 7147 38811
rect 9413 38777 9447 38811
rect 10241 38777 10275 38811
rect 12112 38777 12146 38811
rect 12817 38777 12851 38811
rect 24869 38777 24903 38811
rect 25789 38777 25823 38811
rect 26157 38777 26191 38811
rect 29653 38777 29687 38811
rect 2789 38709 2823 38743
rect 10977 38709 11011 38743
rect 15669 38709 15703 38743
rect 23857 38709 23891 38743
rect 28457 38709 28491 38743
rect 30389 38709 30423 38743
rect 1777 38505 1811 38539
rect 5273 38505 5307 38539
rect 8125 38505 8159 38539
rect 9781 38505 9815 38539
rect 11621 38505 11655 38539
rect 14749 38505 14783 38539
rect 15577 38505 15611 38539
rect 16037 38505 16071 38539
rect 16839 38505 16873 38539
rect 18245 38505 18279 38539
rect 31217 38505 31251 38539
rect 10885 38437 10919 38471
rect 12909 38437 12943 38471
rect 13614 38437 13648 38471
rect 15669 38437 15703 38471
rect 17049 38437 17083 38471
rect 23958 38437 23992 38471
rect 26249 38437 26283 38471
rect 27537 38437 27571 38471
rect 27721 38437 27755 38471
rect 28917 38437 28951 38471
rect 29622 38437 29656 38471
rect 1961 38369 1995 38403
rect 2237 38369 2271 38403
rect 2329 38369 2363 38403
rect 2513 38369 2547 38403
rect 3249 38369 3283 38403
rect 3893 38369 3927 38403
rect 4077 38369 4111 38403
rect 4169 38369 4203 38403
rect 4445 38369 4479 38403
rect 5549 38369 5583 38403
rect 6745 38369 6779 38403
rect 7012 38369 7046 38403
rect 8585 38369 8619 38403
rect 8769 38369 8803 38403
rect 9045 38369 9079 38403
rect 9137 38369 9171 38403
rect 9321 38369 9355 38403
rect 10057 38369 10091 38403
rect 10333 38369 10367 38403
rect 10977 38369 11011 38403
rect 11529 38369 11563 38403
rect 12173 38369 12207 38403
rect 12357 38369 12391 38403
rect 12541 38369 12575 38403
rect 12725 38369 12759 38403
rect 17509 38369 17543 38403
rect 17693 38369 17727 38403
rect 17877 38369 17911 38403
rect 18061 38369 18095 38403
rect 18705 38369 18739 38403
rect 18889 38369 18923 38403
rect 20076 38369 20110 38403
rect 22109 38369 22143 38403
rect 24685 38369 24719 38403
rect 24869 38369 24903 38403
rect 24961 38369 24995 38403
rect 25237 38369 25271 38403
rect 26433 38369 26467 38403
rect 27353 38369 27387 38403
rect 28181 38369 28215 38403
rect 28365 38369 28399 38403
rect 28457 38369 28491 38403
rect 28733 38369 28767 38403
rect 2145 38301 2179 38335
rect 4261 38301 4295 38335
rect 5273 38301 5307 38335
rect 8953 38301 8987 38335
rect 12449 38301 12483 38335
rect 13369 38301 13403 38335
rect 15485 38301 15519 38335
rect 17785 38301 17819 38335
rect 19809 38301 19843 38335
rect 24225 38301 24259 38335
rect 25053 38301 25087 38335
rect 28549 38301 28583 38335
rect 29377 38301 29411 38335
rect 3341 38233 3375 38267
rect 5457 38233 5491 38267
rect 16681 38233 16715 38267
rect 18705 38233 18739 38267
rect 4629 38165 4663 38199
rect 10057 38165 10091 38199
rect 16865 38165 16899 38199
rect 21189 38165 21223 38199
rect 22201 38165 22235 38199
rect 22845 38165 22879 38199
rect 25421 38165 25455 38199
rect 26065 38165 26099 38199
rect 30757 38165 30791 38199
rect 5549 37961 5583 37995
rect 7021 37961 7055 37995
rect 9045 37961 9079 37995
rect 9689 37961 9723 37995
rect 15301 37961 15335 37995
rect 20085 37961 20119 37995
rect 20637 37961 20671 37995
rect 22477 37961 22511 37995
rect 24777 37961 24811 37995
rect 26709 37961 26743 37995
rect 27353 37961 27387 37995
rect 14749 37893 14783 37927
rect 18613 37893 18647 37927
rect 21281 37893 21315 37927
rect 4261 37825 4295 37859
rect 7113 37825 7147 37859
rect 10885 37825 10919 37859
rect 10977 37825 11011 37859
rect 11989 37825 12023 37859
rect 15761 37825 15795 37859
rect 17325 37825 17359 37859
rect 19625 37825 19659 37859
rect 21833 37825 21867 37859
rect 23406 37825 23440 37859
rect 23857 37825 23891 37859
rect 29561 37825 29595 37859
rect 1869 37757 1903 37791
rect 3985 37757 4019 37791
rect 4169 37757 4203 37791
rect 4353 37757 4387 37791
rect 4537 37757 4571 37791
rect 6837 37757 6871 37791
rect 6929 37757 6963 37791
rect 7573 37757 7607 37791
rect 8953 37757 8987 37791
rect 9873 37757 9907 37791
rect 10701 37757 10735 37791
rect 11069 37757 11103 37791
rect 11253 37757 11287 37791
rect 11713 37757 11747 37791
rect 11897 37757 11931 37791
rect 12081 37757 12115 37791
rect 12265 37757 12299 37791
rect 13001 37757 13035 37791
rect 14657 37757 14691 37791
rect 15485 37757 15519 37791
rect 15577 37757 15611 37791
rect 15669 37757 15703 37791
rect 15945 37757 15979 37791
rect 17141 37757 17175 37791
rect 17417 37757 17451 37791
rect 17509 37757 17543 37791
rect 17693 37757 17727 37791
rect 18521 37757 18555 37791
rect 19349 37757 19383 37791
rect 19533 37757 19567 37791
rect 19717 37757 19751 37791
rect 19901 37757 19935 37791
rect 21097 37757 21131 37791
rect 22109 37757 22143 37791
rect 23121 37757 23155 37791
rect 23305 37757 23339 37791
rect 23489 37757 23523 37791
rect 23673 37757 23707 37791
rect 25890 37757 25924 37791
rect 26157 37757 26191 37791
rect 26801 37757 26835 37791
rect 27261 37757 27295 37791
rect 27537 37757 27571 37791
rect 27629 37757 27663 37791
rect 28273 37757 28307 37791
rect 28457 37757 28491 37791
rect 28543 37757 28577 37791
rect 28687 37757 28721 37791
rect 28825 37757 28859 37791
rect 2237 37689 2271 37723
rect 10057 37689 10091 37723
rect 16497 37689 16531 37723
rect 29009 37689 29043 37723
rect 29806 37689 29840 37723
rect 2697 37621 2731 37655
rect 3801 37621 3835 37655
rect 5089 37621 5123 37655
rect 6377 37621 6411 37655
rect 8125 37621 8159 37655
rect 10517 37621 10551 37655
rect 12449 37621 12483 37655
rect 13461 37621 13495 37655
rect 14105 37621 14139 37655
rect 16957 37621 16991 37655
rect 22017 37621 22051 37655
rect 27813 37621 27847 37655
rect 30941 37621 30975 37655
rect 2513 37417 2547 37451
rect 5825 37417 5859 37451
rect 8033 37417 8067 37451
rect 8493 37417 8527 37451
rect 13461 37417 13495 37451
rect 14933 37417 14967 37451
rect 15761 37417 15795 37451
rect 21005 37417 21039 37451
rect 21833 37417 21867 37451
rect 22017 37417 22051 37451
rect 22201 37417 22235 37451
rect 23045 37417 23079 37451
rect 25789 37417 25823 37451
rect 26433 37417 26467 37451
rect 29745 37417 29779 37451
rect 30389 37417 30423 37451
rect 31309 37417 31343 37451
rect 3648 37349 3682 37383
rect 15577 37349 15611 37383
rect 16957 37349 16991 37383
rect 22845 37349 22879 37383
rect 23857 37349 23891 37383
rect 27077 37349 27111 37383
rect 2053 37281 2087 37315
rect 3893 37281 3927 37315
rect 4445 37281 4479 37315
rect 4712 37281 4746 37315
rect 6653 37281 6687 37315
rect 6920 37281 6954 37315
rect 9617 37281 9651 37315
rect 9873 37281 9907 37315
rect 10517 37281 10551 37315
rect 11529 37281 11563 37315
rect 12081 37281 12115 37315
rect 12348 37281 12382 37315
rect 15393 37281 15427 37315
rect 16865 37281 16899 37315
rect 17693 37281 17727 37315
rect 17960 37281 17994 37315
rect 19625 37281 19659 37315
rect 19892 37281 19926 37315
rect 22109 37281 22143 37315
rect 23765 37281 23799 37315
rect 24409 37281 24443 37315
rect 24665 37281 24699 37315
rect 27169 37281 27203 37315
rect 27629 37281 27663 37315
rect 27813 37281 27847 37315
rect 28365 37281 28399 37315
rect 28641 37281 28675 37315
rect 29837 37281 29871 37315
rect 31125 37281 31159 37315
rect 19073 37145 19107 37179
rect 22385 37145 22419 37179
rect 1501 37077 1535 37111
rect 10517 37077 10551 37111
rect 14105 37077 14139 37111
rect 23029 37077 23063 37111
rect 23213 37077 23247 37111
rect 27629 37077 27663 37111
rect 7205 36873 7239 36907
rect 7665 36873 7699 36907
rect 9689 36873 9723 36907
rect 11897 36873 11931 36907
rect 19993 36873 20027 36907
rect 21005 36873 21039 36907
rect 22109 36873 22143 36907
rect 23305 36873 23339 36907
rect 30205 36873 30239 36907
rect 14657 36805 14691 36839
rect 26893 36805 26927 36839
rect 2053 36737 2087 36771
rect 4077 36737 4111 36771
rect 5273 36737 5307 36771
rect 12817 36737 12851 36771
rect 24777 36737 24811 36771
rect 28181 36737 28215 36771
rect 1869 36669 1903 36703
rect 2145 36669 2179 36703
rect 2237 36669 2271 36703
rect 2421 36669 2455 36703
rect 3801 36669 3835 36703
rect 8953 36669 8987 36703
rect 9137 36669 9171 36703
rect 9223 36669 9257 36703
rect 9321 36669 9355 36703
rect 9505 36669 9539 36703
rect 10517 36669 10551 36703
rect 12449 36669 12483 36703
rect 12633 36669 12667 36703
rect 12725 36669 12759 36703
rect 13001 36669 13035 36703
rect 16313 36669 16347 36703
rect 16580 36669 16614 36703
rect 19257 36669 19291 36703
rect 19441 36669 19475 36703
rect 19533 36669 19567 36703
rect 19625 36669 19659 36703
rect 19809 36669 19843 36703
rect 21097 36669 21131 36703
rect 22937 36669 22971 36703
rect 23581 36669 23615 36703
rect 24593 36669 24627 36703
rect 26065 36669 26099 36703
rect 26525 36669 26559 36703
rect 26709 36669 26743 36703
rect 26801 36669 26835 36703
rect 26985 36669 27019 36703
rect 27169 36669 27203 36703
rect 27905 36669 27939 36703
rect 28089 36669 28123 36703
rect 28273 36669 28307 36703
rect 28457 36669 28491 36703
rect 29653 36669 29687 36703
rect 29745 36669 29779 36703
rect 5518 36601 5552 36635
rect 10784 36601 10818 36635
rect 21281 36601 21315 36635
rect 21741 36601 21775 36635
rect 21925 36601 21959 36635
rect 23314 36601 23348 36635
rect 1685 36533 1719 36567
rect 3065 36533 3099 36567
rect 6653 36533 6687 36567
rect 8401 36533 8435 36567
rect 13185 36533 13219 36567
rect 14105 36533 14139 36567
rect 15577 36533 15611 36567
rect 17693 36533 17727 36567
rect 18153 36533 18187 36567
rect 24409 36533 24443 36567
rect 25237 36533 25271 36567
rect 25881 36533 25915 36567
rect 28641 36533 28675 36567
rect 30849 36533 30883 36567
rect 5089 36329 5123 36363
rect 7113 36329 7147 36363
rect 10609 36329 10643 36363
rect 10977 36329 11011 36363
rect 11913 36329 11947 36363
rect 18245 36329 18279 36363
rect 21189 36329 21223 36363
rect 26065 36329 26099 36363
rect 26157 36329 26191 36363
rect 26985 36329 27019 36363
rect 10517 36261 10551 36295
rect 11713 36261 11747 36295
rect 15853 36261 15887 36295
rect 21833 36261 21867 36295
rect 22201 36261 22235 36295
rect 23581 36261 23615 36295
rect 24501 36261 24535 36295
rect 1409 36193 1443 36227
rect 1676 36193 1710 36227
rect 3801 36193 3835 36227
rect 4353 36193 4387 36227
rect 4537 36193 4571 36227
rect 4905 36193 4939 36227
rect 6561 36193 6595 36227
rect 7297 36193 7331 36227
rect 7665 36193 7699 36227
rect 7849 36193 7883 36227
rect 8309 36193 8343 36227
rect 9229 36193 9263 36227
rect 13001 36193 13035 36227
rect 13268 36193 13302 36227
rect 15577 36193 15611 36227
rect 15945 36193 15979 36227
rect 16865 36193 16899 36227
rect 17509 36193 17543 36227
rect 17693 36193 17727 36227
rect 17785 36193 17819 36227
rect 18061 36193 18095 36227
rect 21281 36193 21315 36227
rect 21977 36193 22011 36227
rect 23213 36193 23247 36227
rect 24317 36193 24351 36227
rect 27169 36193 27203 36227
rect 27445 36193 27479 36227
rect 27629 36193 27663 36227
rect 28273 36193 28307 36227
rect 28365 36193 28399 36227
rect 28641 36193 28675 36227
rect 29193 36193 29227 36227
rect 29285 36193 29319 36227
rect 31125 36193 31159 36227
rect 4629 36125 4663 36159
rect 4721 36125 4755 36159
rect 6377 36125 6411 36159
rect 7481 36125 7515 36159
rect 7573 36125 7607 36159
rect 8953 36125 8987 36159
rect 10333 36125 10367 36159
rect 15485 36125 15519 36159
rect 17049 36125 17083 36159
rect 17877 36125 17911 36159
rect 18797 36125 18831 36159
rect 26341 36125 26375 36159
rect 27353 36125 27387 36159
rect 27261 36057 27295 36091
rect 28549 36057 28583 36091
rect 2789 35989 2823 36023
rect 3709 35989 3743 36023
rect 5549 35989 5583 36023
rect 11897 35989 11931 36023
rect 12081 35989 12115 36023
rect 14381 35989 14415 36023
rect 16681 35989 16715 36023
rect 19257 35989 19291 36023
rect 20361 35989 20395 36023
rect 22753 35989 22787 36023
rect 23581 35989 23615 36023
rect 23765 35989 23799 36023
rect 25145 35989 25179 36023
rect 25697 35989 25731 36023
rect 28089 35989 28123 36023
rect 29745 35989 29779 36023
rect 30389 35989 30423 36023
rect 31309 35989 31343 36023
rect 1593 35785 1627 35819
rect 17785 35785 17819 35819
rect 21373 35785 21407 35819
rect 27537 35785 27571 35819
rect 28825 35785 28859 35819
rect 26709 35717 26743 35751
rect 2605 35649 2639 35683
rect 4261 35649 4295 35683
rect 6837 35649 6871 35683
rect 9965 35649 9999 35683
rect 11805 35649 11839 35683
rect 13001 35649 13035 35683
rect 18521 35649 18555 35683
rect 23397 35649 23431 35683
rect 23857 35649 23891 35683
rect 25053 35649 25087 35683
rect 27997 35649 28031 35683
rect 29929 35649 29963 35683
rect 2881 35581 2915 35615
rect 3985 35581 4019 35615
rect 4169 35581 4203 35615
rect 4353 35581 4387 35615
rect 4537 35581 4571 35615
rect 6377 35581 6411 35615
rect 7113 35581 7147 35615
rect 8125 35581 8159 35615
rect 9689 35581 9723 35615
rect 9873 35581 9907 35615
rect 10057 35581 10091 35615
rect 10241 35581 10275 35615
rect 11989 35581 12023 35615
rect 13185 35581 13219 35615
rect 14381 35581 14415 35615
rect 16221 35581 16255 35615
rect 16773 35581 16807 35615
rect 17417 35581 17451 35615
rect 18061 35581 18095 35615
rect 19257 35581 19291 35615
rect 21281 35581 21315 35615
rect 21465 35581 21499 35615
rect 22201 35581 22235 35615
rect 23673 35581 23707 35615
rect 24869 35581 24903 35615
rect 25697 35581 25731 35615
rect 27077 35581 27111 35615
rect 27721 35581 27755 35615
rect 27905 35581 27939 35615
rect 28089 35581 28123 35615
rect 28273 35581 28307 35615
rect 28917 35581 28951 35615
rect 29561 35581 29595 35615
rect 29745 35581 29779 35615
rect 29837 35581 29871 35615
rect 30113 35581 30147 35615
rect 5181 35513 5215 35547
rect 13553 35513 13587 35547
rect 14289 35513 14323 35547
rect 15954 35513 15988 35547
rect 19524 35513 19558 35547
rect 22845 35513 22879 35547
rect 26893 35513 26927 35547
rect 3801 35445 3835 35479
rect 5089 35445 5123 35479
rect 6285 35445 6319 35479
rect 8217 35445 8251 35479
rect 9229 35445 9263 35479
rect 10425 35445 10459 35479
rect 10885 35445 10919 35479
rect 12173 35445 12207 35479
rect 13277 35445 13311 35479
rect 13369 35445 13403 35479
rect 14841 35445 14875 35479
rect 16957 35445 16991 35479
rect 17794 35445 17828 35479
rect 20637 35445 20671 35479
rect 22385 35445 22419 35479
rect 25605 35445 25639 35479
rect 30297 35445 30331 35479
rect 30757 35445 30791 35479
rect 2053 35241 2087 35275
rect 9505 35241 9539 35275
rect 13829 35241 13863 35275
rect 15485 35241 15519 35275
rect 23857 35241 23891 35275
rect 24869 35241 24903 35275
rect 26985 35241 27019 35275
rect 2145 35173 2179 35207
rect 10618 35173 10652 35207
rect 13124 35173 13158 35207
rect 18705 35173 18739 35207
rect 2697 35105 2731 35139
rect 3341 35105 3375 35139
rect 3608 35105 3642 35139
rect 5365 35105 5399 35139
rect 6377 35105 6411 35139
rect 7113 35105 7147 35139
rect 7573 35105 7607 35139
rect 7840 35105 7874 35139
rect 10885 35105 10919 35139
rect 13369 35105 13403 35139
rect 14013 35105 14047 35139
rect 14749 35105 14783 35139
rect 14933 35105 14967 35139
rect 15117 35105 15151 35139
rect 15301 35105 15335 35139
rect 16681 35105 16715 35139
rect 16948 35105 16982 35139
rect 19073 35105 19107 35139
rect 19625 35105 19659 35139
rect 19809 35105 19843 35139
rect 19901 35105 19935 35139
rect 20177 35105 20211 35139
rect 21097 35105 21131 35139
rect 21925 35105 21959 35139
rect 22017 35105 22051 35139
rect 22733 35105 22767 35139
rect 25982 35105 26016 35139
rect 27353 35105 27387 35139
rect 27997 35105 28031 35139
rect 30674 35105 30708 35139
rect 15025 35037 15059 35071
rect 19993 35037 20027 35071
rect 22477 35037 22511 35071
rect 26249 35037 26283 35071
rect 27261 35037 27295 35071
rect 28273 35037 28307 35071
rect 30941 35037 30975 35071
rect 4721 34969 4755 35003
rect 15945 34969 15979 35003
rect 18061 34969 18095 35003
rect 21189 34969 21223 35003
rect 2789 34901 2823 34935
rect 5273 34901 5307 34935
rect 6469 34901 6503 34935
rect 8953 34901 8987 34935
rect 11989 34901 12023 34935
rect 18521 34901 18555 34935
rect 18705 34901 18739 34935
rect 20361 34901 20395 34935
rect 24317 34901 24351 34935
rect 27261 34901 27295 34935
rect 29561 34901 29595 34935
rect 7941 34697 7975 34731
rect 10333 34697 10367 34731
rect 11713 34697 11747 34731
rect 13369 34697 13403 34731
rect 13553 34697 13587 34731
rect 14749 34697 14783 34731
rect 14933 34697 14967 34731
rect 15393 34697 15427 34731
rect 26157 34697 26191 34731
rect 29561 34697 29595 34731
rect 2973 34629 3007 34663
rect 5457 34629 5491 34663
rect 11069 34629 11103 34663
rect 13001 34629 13035 34663
rect 25605 34629 25639 34663
rect 6745 34561 6779 34595
rect 7481 34561 7515 34595
rect 8953 34561 8987 34595
rect 15761 34561 15795 34595
rect 16865 34561 16899 34595
rect 17785 34561 17819 34595
rect 18705 34561 18739 34595
rect 19349 34561 19383 34595
rect 25145 34561 25179 34595
rect 28733 34561 28767 34595
rect 30941 34561 30975 34595
rect 1593 34493 1627 34527
rect 2053 34493 2087 34527
rect 2237 34493 2271 34527
rect 4537 34493 4571 34527
rect 4813 34493 4847 34527
rect 5273 34493 5307 34527
rect 5457 34493 5491 34527
rect 6469 34493 6503 34527
rect 6561 34493 6595 34527
rect 7205 34493 7239 34527
rect 7389 34493 7423 34527
rect 7573 34493 7607 34527
rect 7757 34493 7791 34527
rect 9229 34493 9263 34527
rect 10977 34493 11011 34527
rect 14381 34493 14415 34527
rect 15577 34493 15611 34527
rect 15853 34493 15887 34527
rect 15945 34493 15979 34527
rect 16129 34493 16163 34527
rect 18061 34493 18095 34527
rect 18429 34493 18463 34527
rect 20177 34493 20211 34527
rect 22017 34493 22051 34527
rect 22273 34493 22307 34527
rect 24869 34493 24903 34527
rect 25053 34493 25087 34527
rect 25237 34493 25271 34527
rect 25421 34493 25455 34527
rect 26065 34493 26099 34527
rect 29009 34493 29043 34527
rect 30674 34493 30708 34527
rect 2789 34425 2823 34459
rect 10425 34425 10459 34459
rect 11989 34425 12023 34459
rect 13369 34425 13403 34459
rect 16681 34425 16715 34459
rect 20444 34425 20478 34459
rect 27261 34425 27295 34459
rect 2145 34357 2179 34391
rect 5917 34357 5951 34391
rect 6745 34357 6779 34391
rect 14749 34357 14783 34391
rect 21557 34357 21591 34391
rect 23397 34357 23431 34391
rect 27169 34357 27203 34391
rect 6377 34153 6411 34187
rect 6837 34153 6871 34187
rect 15761 34153 15795 34187
rect 19441 34153 19475 34187
rect 20729 34153 20763 34187
rect 23857 34153 23891 34187
rect 27537 34153 27571 34187
rect 28181 34153 28215 34187
rect 29745 34153 29779 34187
rect 30297 34153 30331 34187
rect 2605 34085 2639 34119
rect 4629 34085 4663 34119
rect 6745 34085 6779 34119
rect 9045 34085 9079 34119
rect 10393 34085 10427 34119
rect 10609 34085 10643 34119
rect 13461 34085 13495 34119
rect 23673 34085 23707 34119
rect 24317 34085 24351 34119
rect 25789 34085 25823 34119
rect 26166 34085 26200 34119
rect 1409 34017 1443 34051
rect 2697 34017 2731 34051
rect 3985 34017 4019 34051
rect 4537 34017 4571 34051
rect 4721 34017 4755 34051
rect 5181 34017 5215 34051
rect 5365 34017 5399 34051
rect 5457 34017 5491 34051
rect 5595 34017 5629 34051
rect 7941 34017 7975 34051
rect 12357 34017 12391 34051
rect 15853 34017 15887 34051
rect 18705 34017 18739 34051
rect 18889 34017 18923 34051
rect 19073 34017 19107 34051
rect 19257 34017 19291 34051
rect 19993 34017 20027 34051
rect 20177 34017 20211 34051
rect 20545 34017 20579 34051
rect 22017 34017 22051 34051
rect 22385 34017 22419 34051
rect 22569 34017 22603 34051
rect 25145 34017 25179 34051
rect 27445 34017 27479 34051
rect 28273 34017 28307 34051
rect 29009 34017 29043 34051
rect 29193 34017 29227 34051
rect 29285 34017 29319 34051
rect 29561 34017 29595 34051
rect 30389 34017 30423 34051
rect 31125 34017 31159 34051
rect 2513 33949 2547 33983
rect 6929 33949 6963 33983
rect 8861 33949 8895 33983
rect 8953 33949 8987 33983
rect 15117 33949 15151 33983
rect 17785 33949 17819 33983
rect 18981 33949 19015 33983
rect 20269 33949 20303 33983
rect 20361 33949 20395 33983
rect 22201 33949 22235 33983
rect 22293 33949 22327 33983
rect 24869 33949 24903 33983
rect 25329 33949 25363 33983
rect 29377 33949 29411 33983
rect 8125 33881 8159 33915
rect 17325 33881 17359 33915
rect 21189 33881 21223 33915
rect 23305 33881 23339 33915
rect 26341 33881 26375 33915
rect 1593 33813 1627 33847
rect 3065 33813 3099 33847
rect 3893 33813 3927 33847
rect 5825 33813 5859 33847
rect 9413 33813 9447 33847
rect 10241 33813 10275 33847
rect 10425 33813 10459 33847
rect 12081 33813 12115 33847
rect 13001 33813 13035 33847
rect 16773 33813 16807 33847
rect 21833 33813 21867 33847
rect 23673 33813 23707 33847
rect 26157 33813 26191 33847
rect 31309 33813 31343 33847
rect 3065 33609 3099 33643
rect 4537 33609 4571 33643
rect 6469 33609 6503 33643
rect 13461 33609 13495 33643
rect 20821 33609 20855 33643
rect 21465 33609 21499 33643
rect 30757 33609 30791 33643
rect 7297 33541 7331 33575
rect 10701 33541 10735 33575
rect 20453 33541 20487 33575
rect 25973 33541 26007 33575
rect 2053 33405 2087 33439
rect 2145 33405 2179 33439
rect 2237 33405 2271 33439
rect 2421 33405 2455 33439
rect 3801 33405 3835 33439
rect 5437 33405 5471 33439
rect 5549 33405 5583 33439
rect 5641 33405 5675 33439
rect 5825 33405 5859 33439
rect 2881 33337 2915 33371
rect 6285 33337 6319 33371
rect 6485 33337 6519 33371
rect 9321 33473 9355 33507
rect 9781 33473 9815 33507
rect 11989 33473 12023 33507
rect 15945 33473 15979 33507
rect 19527 33473 19561 33507
rect 21741 33473 21775 33507
rect 21925 33473 21959 33507
rect 23213 33473 23247 33507
rect 25053 33473 25087 33507
rect 28181 33473 28215 33507
rect 28273 33473 28307 33507
rect 29837 33473 29871 33507
rect 29929 33473 29963 33507
rect 7665 33405 7699 33439
rect 7757 33405 7791 33439
rect 7849 33405 7883 33439
rect 8033 33405 8067 33439
rect 8953 33405 8987 33439
rect 9229 33405 9263 33439
rect 10701 33405 10735 33439
rect 10885 33405 10919 33439
rect 11529 33405 11563 33439
rect 11713 33405 11747 33439
rect 11897 33405 11931 33439
rect 12081 33405 12115 33439
rect 12265 33405 12299 33439
rect 12725 33405 12759 33439
rect 14105 33405 14139 33439
rect 17785 33405 17819 33439
rect 18521 33405 18555 33439
rect 19261 33395 19295 33429
rect 19441 33405 19475 33439
rect 19625 33405 19659 33439
rect 19809 33405 19843 33439
rect 21649 33405 21683 33439
rect 21833 33405 21867 33439
rect 22937 33405 22971 33439
rect 24777 33405 24811 33439
rect 24961 33405 24995 33439
rect 25145 33405 25179 33439
rect 25329 33405 25363 33439
rect 27353 33405 27387 33439
rect 27997 33405 28031 33439
rect 28365 33405 28399 33439
rect 28549 33405 28583 33439
rect 29561 33405 29595 33439
rect 29745 33405 29779 33439
rect 30113 33405 30147 33439
rect 9597 33337 9631 33371
rect 11069 33337 11103 33371
rect 12817 33337 12851 33371
rect 14350 33337 14384 33371
rect 16190 33337 16224 33371
rect 17877 33337 17911 33371
rect 18613 33337 18647 33371
rect 27086 33337 27120 33371
rect 1777 33269 1811 33303
rect 3081 33269 3115 33303
rect 3249 33269 3283 33303
rect 3893 33269 3927 33303
rect 5181 33269 5215 33303
rect 6653 33269 6687 33303
rect 7297 33269 7331 33303
rect 7389 33269 7423 33303
rect 15485 33269 15519 33303
rect 17325 33269 17359 33303
rect 19993 33269 20027 33303
rect 20821 33269 20855 33303
rect 21005 33269 21039 33303
rect 25513 33269 25547 33303
rect 27813 33269 27847 33303
rect 30297 33269 30331 33303
rect 10425 33065 10459 33099
rect 11621 33065 11655 33099
rect 13829 33065 13863 33099
rect 15761 33065 15795 33099
rect 17693 33065 17727 33099
rect 22385 33065 22419 33099
rect 24317 33065 24351 33099
rect 24869 33065 24903 33099
rect 25329 33065 25363 33099
rect 7757 32997 7791 33031
rect 10609 32997 10643 33031
rect 17141 32997 17175 33031
rect 18828 32997 18862 33031
rect 19533 32997 19567 33031
rect 21281 32997 21315 33031
rect 1777 32929 1811 32963
rect 1869 32929 1903 32963
rect 1961 32929 1995 32963
rect 2145 32929 2179 32963
rect 2881 32929 2915 32963
rect 3525 32929 3559 32963
rect 3893 32929 3927 32963
rect 4629 32929 4663 32963
rect 5365 32929 5399 32963
rect 6469 32929 6503 32963
rect 7205 32929 7239 32963
rect 8493 32929 8527 32963
rect 9321 32929 9355 32963
rect 10977 32929 11011 32963
rect 12633 32929 12667 32963
rect 12817 32929 12851 32963
rect 12909 32929 12943 32963
rect 13185 32929 13219 32963
rect 14013 32929 14047 32963
rect 14197 32929 14231 32963
rect 14381 32929 14415 32963
rect 14565 32929 14599 32963
rect 15025 32929 15059 32963
rect 15209 32929 15243 32963
rect 15393 32929 15427 32963
rect 15577 32929 15611 32963
rect 16865 32929 16899 32963
rect 17233 32929 17267 32963
rect 19717 32929 19751 32963
rect 19855 32929 19889 32963
rect 20085 32929 20119 32963
rect 20269 32929 20303 32963
rect 20729 32929 20763 32963
rect 20913 32929 20947 32963
rect 22201 32929 22235 32963
rect 22937 32929 22971 32963
rect 23204 32929 23238 32963
rect 25421 32929 25455 32963
rect 25605 32929 25639 32963
rect 25789 32929 25823 32963
rect 25973 32929 26007 32963
rect 26157 32929 26191 32963
rect 27169 32929 27203 32963
rect 28089 32929 28123 32963
rect 29561 32929 29595 32963
rect 29745 32929 29779 32963
rect 29929 32929 29963 32963
rect 30113 32929 30147 32963
rect 3157 32861 3191 32895
rect 4905 32861 4939 32895
rect 5457 32861 5491 32895
rect 5641 32861 5675 32895
rect 6653 32861 6687 32895
rect 6745 32861 6779 32895
rect 8769 32861 8803 32895
rect 9505 32861 9539 32895
rect 13001 32861 13035 32895
rect 14289 32861 14323 32895
rect 15301 32861 15335 32895
rect 16681 32861 16715 32895
rect 19073 32861 19107 32895
rect 19993 32861 20027 32895
rect 25329 32861 25363 32895
rect 25697 32861 25731 32895
rect 27353 32861 27387 32895
rect 28365 32861 28399 32895
rect 29837 32861 29871 32895
rect 3341 32793 3375 32827
rect 7113 32793 7147 32827
rect 8953 32793 8987 32827
rect 21189 32793 21223 32827
rect 26985 32793 27019 32827
rect 31125 32793 31159 32827
rect 1501 32725 1535 32759
rect 4721 32725 4755 32759
rect 4813 32725 4847 32759
rect 5549 32725 5583 32759
rect 10609 32725 10643 32759
rect 12173 32725 12207 32759
rect 13369 32725 13403 32759
rect 29377 32725 29411 32759
rect 30573 32725 30607 32759
rect 1777 32521 1811 32555
rect 3801 32521 3835 32555
rect 7757 32521 7791 32555
rect 9137 32521 9171 32555
rect 9689 32521 9723 32555
rect 14565 32521 14599 32555
rect 15577 32521 15611 32555
rect 21373 32521 21407 32555
rect 22661 32521 22695 32555
rect 23581 32521 23615 32555
rect 24869 32521 24903 32555
rect 27353 32521 27387 32555
rect 29561 32521 29595 32555
rect 3157 32453 3191 32487
rect 4537 32453 4571 32487
rect 6561 32453 6595 32487
rect 13185 32453 13219 32487
rect 15209 32453 15243 32487
rect 15761 32453 15795 32487
rect 1685 32385 1719 32419
rect 1869 32385 1903 32419
rect 2513 32385 2547 32419
rect 2789 32385 2823 32419
rect 3249 32385 3283 32419
rect 6377 32385 6411 32419
rect 10977 32385 11011 32419
rect 11805 32385 11839 32419
rect 14105 32385 14139 32419
rect 18337 32385 18371 32419
rect 19073 32385 19107 32419
rect 20453 32385 20487 32419
rect 20913 32385 20947 32419
rect 1961 32317 1995 32351
rect 2697 32317 2731 32351
rect 3801 32317 3835 32351
rect 3985 32317 4019 32351
rect 4445 32317 4479 32351
rect 5089 32317 5123 32351
rect 6101 32317 6135 32351
rect 6837 32317 6871 32351
rect 7205 32317 7239 32351
rect 8033 32317 8067 32351
rect 8125 32317 8159 32351
rect 8238 32314 8272 32348
rect 8401 32317 8435 32351
rect 8953 32317 8987 32351
rect 9137 32317 9171 32351
rect 9597 32317 9631 32351
rect 10793 32317 10827 32351
rect 11069 32317 11103 32351
rect 11161 32317 11195 32351
rect 11345 32317 11379 32351
rect 14289 32317 14323 32351
rect 16221 32317 16255 32351
rect 16405 32317 16439 32351
rect 16589 32317 16623 32351
rect 16681 32317 16715 32351
rect 16773 32317 16807 32351
rect 16957 32317 16991 32351
rect 12050 32249 12084 32283
rect 14657 32249 14691 32283
rect 17509 32249 17543 32283
rect 19717 32317 19751 32351
rect 20177 32317 20211 32351
rect 20361 32317 20395 32351
rect 20545 32317 20579 32351
rect 20729 32317 20763 32351
rect 19625 32249 19659 32283
rect 5181 32181 5215 32215
rect 10609 32181 10643 32215
rect 15577 32181 15611 32215
rect 17601 32181 17635 32215
rect 19073 32181 19107 32215
rect 25053 32453 25087 32487
rect 30941 32385 30975 32419
rect 21465 32317 21499 32351
rect 21649 32317 21683 32351
rect 21741 32317 21775 32351
rect 21833 32317 21867 32351
rect 22017 32317 22051 32351
rect 23765 32317 23799 32351
rect 25513 32317 25547 32351
rect 25780 32317 25814 32351
rect 28466 32317 28500 32351
rect 28733 32317 28767 32351
rect 24685 32249 24719 32283
rect 24885 32249 24919 32283
rect 30674 32249 30708 32283
rect 21373 32181 21407 32215
rect 22201 32181 22235 32215
rect 26893 32181 26927 32215
rect 1961 31977 1995 32011
rect 7573 31977 7607 32011
rect 10977 31977 11011 32011
rect 11897 31977 11931 32011
rect 13461 31977 13495 32011
rect 13645 31977 13679 32011
rect 23765 31977 23799 32011
rect 26985 31977 27019 32011
rect 27537 31977 27571 32011
rect 28825 31977 28859 32011
rect 1501 31909 1535 31943
rect 2789 31909 2823 31943
rect 3801 31909 3835 31943
rect 4537 31909 4571 31943
rect 4753 31909 4787 31943
rect 8125 31909 8159 31943
rect 9864 31909 9898 31943
rect 14197 31909 14231 31943
rect 18245 31909 18279 31943
rect 29938 31909 29972 31943
rect 2237 31841 2271 31875
rect 2697 31841 2731 31875
rect 4077 31841 4111 31875
rect 5365 31841 5399 31875
rect 7297 31841 7331 31875
rect 8217 31841 8251 31875
rect 8677 31841 8711 31875
rect 8769 31841 8803 31875
rect 8861 31841 8895 31875
rect 12081 31841 12115 31875
rect 12449 31841 12483 31875
rect 12633 31841 12667 31875
rect 13093 31841 13127 31875
rect 14105 31841 14139 31875
rect 15209 31841 15243 31875
rect 15393 31841 15427 31875
rect 15589 31847 15623 31881
rect 15761 31841 15795 31875
rect 16957 31841 16991 31875
rect 17141 31841 17175 31875
rect 17509 31841 17543 31875
rect 18153 31841 18187 31875
rect 20637 31841 20671 31875
rect 21005 31841 21039 31875
rect 21189 31841 21223 31875
rect 22946 31841 22980 31875
rect 23213 31841 23247 31875
rect 24889 31841 24923 31875
rect 25145 31841 25179 31875
rect 25605 31841 25639 31875
rect 25789 31841 25823 31875
rect 25973 31841 26007 31875
rect 26157 31841 26191 31875
rect 30205 31841 30239 31875
rect 31125 31841 31159 31875
rect 1961 31773 1995 31807
rect 3801 31773 3835 31807
rect 6377 31773 6411 31807
rect 7573 31773 7607 31807
rect 9597 31773 9631 31807
rect 12265 31773 12299 31807
rect 12357 31773 12391 31807
rect 15485 31773 15519 31807
rect 17233 31773 17267 31807
rect 17325 31773 17359 31807
rect 17693 31773 17727 31807
rect 19165 31773 19199 31807
rect 19441 31773 19475 31807
rect 20821 31773 20855 31807
rect 20913 31773 20947 31807
rect 25881 31773 25915 31807
rect 28089 31773 28123 31807
rect 21833 31705 21867 31739
rect 2145 31637 2179 31671
rect 3985 31637 4019 31671
rect 4721 31637 4755 31671
rect 4905 31637 4939 31671
rect 5457 31637 5491 31671
rect 7389 31637 7423 31671
rect 13461 31637 13495 31671
rect 15025 31637 15059 31671
rect 20453 31637 20487 31671
rect 26341 31637 26375 31671
rect 31309 31637 31343 31671
rect 3893 31433 3927 31467
rect 7021 31433 7055 31467
rect 7665 31433 7699 31467
rect 8217 31433 8251 31467
rect 13185 31433 13219 31467
rect 16957 31433 16991 31467
rect 21557 31433 21591 31467
rect 26341 31433 26375 31467
rect 28733 31433 28767 31467
rect 30757 31433 30791 31467
rect 2053 31365 2087 31399
rect 5089 31365 5123 31399
rect 10885 31365 10919 31399
rect 12541 31365 12575 31399
rect 16589 31365 16623 31399
rect 17141 31365 17175 31399
rect 23397 31365 23431 31399
rect 3249 31297 3283 31331
rect 4905 31297 4939 31331
rect 5181 31297 5215 31331
rect 8953 31297 8987 31331
rect 11805 31297 11839 31331
rect 18705 31297 18739 31331
rect 20177 31297 20211 31331
rect 24961 31297 24995 31331
rect 25053 31297 25087 31331
rect 1869 31229 1903 31263
rect 2973 31229 3007 31263
rect 3065 31229 3099 31263
rect 4629 31229 4663 31263
rect 5273 31229 5307 31263
rect 6469 31229 6503 31263
rect 7573 31229 7607 31263
rect 9505 31229 9539 31263
rect 11529 31229 11563 31263
rect 11713 31229 11747 31263
rect 11897 31229 11931 31263
rect 12081 31229 12115 31263
rect 14841 31229 14875 31263
rect 15117 31229 15151 31263
rect 17785 31229 17819 31263
rect 17969 31229 18003 31263
rect 18429 31229 18463 31263
rect 19717 31229 19751 31263
rect 20444 31229 20478 31263
rect 22017 31229 22051 31263
rect 22284 31229 22318 31263
rect 24777 31229 24811 31263
rect 25145 31229 25179 31263
rect 25329 31229 25363 31263
rect 29561 31365 29595 31399
rect 26709 31297 26743 31331
rect 28181 31297 28215 31331
rect 26433 31229 26467 31263
rect 26617 31229 26651 31263
rect 26801 31229 26835 31263
rect 26985 31229 27019 31263
rect 3249 31161 3283 31195
rect 9772 31161 9806 31195
rect 11345 31161 11379 31195
rect 19625 31161 19659 31195
rect 26341 31161 26375 31195
rect 6377 31093 6411 31127
rect 14381 31093 14415 31127
rect 16957 31093 16991 31127
rect 24593 31093 24627 31127
rect 25789 31093 25823 31127
rect 27169 31093 27203 31127
rect 27629 31093 27663 31127
rect 30205 31093 30239 31127
rect 31217 31093 31251 31127
rect 2605 30889 2639 30923
rect 3801 30889 3835 30923
rect 5089 30889 5123 30923
rect 6929 30889 6963 30923
rect 8861 30889 8895 30923
rect 9321 30889 9355 30923
rect 10977 30889 11011 30923
rect 16129 30889 16163 30923
rect 22569 30889 22603 30923
rect 23029 30889 23063 30923
rect 29377 30889 29411 30923
rect 2053 30821 2087 30855
rect 9873 30821 9907 30855
rect 15016 30821 15050 30855
rect 18245 30821 18279 30855
rect 31033 30821 31067 30855
rect 1869 30753 1903 30787
rect 2697 30753 2731 30787
rect 3157 30753 3191 30787
rect 3341 30753 3375 30787
rect 3433 30753 3467 30787
rect 3525 30753 3559 30787
rect 4537 30753 4571 30787
rect 4997 30753 5031 30787
rect 5549 30753 5583 30787
rect 5733 30753 5767 30787
rect 6745 30753 6779 30787
rect 7748 30753 7782 30787
rect 14013 30753 14047 30787
rect 14749 30753 14783 30787
rect 17049 30753 17083 30787
rect 17233 30753 17267 30787
rect 17601 30753 17635 30787
rect 20729 30753 20763 30787
rect 21833 30753 21867 30787
rect 22017 30753 22051 30787
rect 22385 30753 22419 30787
rect 23305 30753 23339 30787
rect 23489 30753 23523 30787
rect 24225 30753 24259 30787
rect 25237 30753 25271 30787
rect 27077 30753 27111 30787
rect 27261 30753 27295 30787
rect 27445 30753 27479 30787
rect 27629 30753 27663 30787
rect 29929 30753 29963 30787
rect 4261 30685 4295 30719
rect 4721 30685 4755 30719
rect 7481 30685 7515 30719
rect 12449 30685 12483 30719
rect 12725 30685 12759 30719
rect 14289 30685 14323 30719
rect 17325 30685 17359 30719
rect 17417 30685 17451 30719
rect 20453 30685 20487 30719
rect 22109 30685 22143 30719
rect 22201 30685 22235 30719
rect 23213 30685 23247 30719
rect 23397 30685 23431 30719
rect 25513 30685 25547 30719
rect 27353 30685 27387 30719
rect 28273 30685 28307 30719
rect 28917 30685 28951 30719
rect 5549 30549 5583 30583
rect 17785 30549 17819 30583
rect 19533 30549 19567 30583
rect 24133 30549 24167 30583
rect 25973 30549 26007 30583
rect 27813 30549 27847 30583
rect 30573 30549 30607 30583
rect 6285 30345 6319 30379
rect 8033 30345 8067 30379
rect 8953 30345 8987 30379
rect 16267 30345 16301 30379
rect 3249 30277 3283 30311
rect 5089 30277 5123 30311
rect 18705 30277 18739 30311
rect 24961 30277 24995 30311
rect 28089 30277 28123 30311
rect 28641 30277 28675 30311
rect 30849 30277 30883 30311
rect 4537 30209 4571 30243
rect 4629 30209 4663 30243
rect 7573 30209 7607 30243
rect 7665 30209 7699 30243
rect 12173 30209 12207 30243
rect 16037 30209 16071 30243
rect 19717 30209 19751 30243
rect 22661 30209 22695 30243
rect 1961 30141 1995 30175
rect 2053 30141 2087 30175
rect 2145 30141 2179 30175
rect 2329 30141 2363 30175
rect 3065 30141 3099 30175
rect 3249 30141 3283 30175
rect 5641 30141 5675 30175
rect 7297 30141 7331 30175
rect 7481 30141 7515 30175
rect 7849 30141 7883 30175
rect 10333 30141 10367 30175
rect 11345 30141 11379 30175
rect 15577 30141 15611 30175
rect 17325 30141 17359 30175
rect 19993 30141 20027 30175
rect 21005 30141 21039 30175
rect 21281 30141 21315 30175
rect 22293 30141 22327 30175
rect 22477 30141 22511 30175
rect 22569 30141 22603 30175
rect 22845 30141 22879 30175
rect 24777 30141 24811 30175
rect 25421 30141 25455 30175
rect 25697 30141 25731 30175
rect 26709 30141 26743 30175
rect 28549 30141 28583 30175
rect 4721 30073 4755 30107
rect 6253 30073 6287 30107
rect 6469 30073 6503 30107
rect 10066 30073 10100 30107
rect 12440 30073 12474 30107
rect 15310 30073 15344 30107
rect 17592 30073 17626 30107
rect 26976 30073 27010 30107
rect 29561 30073 29595 30107
rect 1685 30005 1719 30039
rect 3893 30005 3927 30039
rect 6101 30005 6135 30039
rect 10793 30005 10827 30039
rect 11437 30005 11471 30039
rect 13553 30005 13587 30039
rect 14197 30005 14231 30039
rect 23029 30005 23063 30039
rect 23581 30005 23615 30039
rect 3801 29801 3835 29835
rect 5549 29801 5583 29835
rect 6745 29801 6779 29835
rect 8309 29801 8343 29835
rect 10793 29801 10827 29835
rect 12633 29801 12667 29835
rect 15945 29801 15979 29835
rect 18061 29801 18095 29835
rect 11989 29733 12023 29767
rect 16037 29733 16071 29767
rect 23765 29733 23799 29767
rect 28558 29733 28592 29767
rect 2145 29665 2179 29699
rect 2237 29665 2271 29699
rect 2329 29665 2363 29699
rect 2513 29665 2547 29699
rect 3249 29665 3283 29699
rect 4077 29665 4111 29699
rect 4169 29665 4203 29699
rect 4261 29665 4295 29699
rect 4445 29665 4479 29699
rect 5457 29665 5491 29699
rect 5825 29665 5859 29699
rect 6653 29665 6687 29699
rect 7573 29665 7607 29699
rect 7757 29665 7791 29699
rect 8125 29665 8159 29699
rect 8769 29665 8803 29699
rect 9680 29665 9714 29699
rect 11713 29665 11747 29699
rect 12081 29665 12115 29699
rect 13093 29665 13127 29699
rect 13265 29665 13299 29699
rect 13461 29665 13495 29699
rect 13645 29665 13679 29699
rect 14841 29665 14875 29699
rect 16681 29665 16715 29699
rect 16948 29665 16982 29699
rect 18889 29665 18923 29699
rect 21833 29665 21867 29699
rect 22017 29667 22051 29701
rect 22201 29665 22235 29699
rect 22385 29665 22419 29699
rect 25513 29665 25547 29699
rect 26157 29665 26191 29699
rect 28825 29665 28859 29699
rect 30398 29665 30432 29699
rect 30665 29665 30699 29699
rect 31125 29665 31159 29699
rect 2973 29597 3007 29631
rect 5641 29597 5675 29631
rect 6469 29597 6503 29631
rect 7849 29597 7883 29631
rect 7941 29597 7975 29631
rect 9413 29597 9447 29631
rect 11621 29597 11655 29631
rect 13363 29597 13397 29631
rect 14565 29597 14599 29631
rect 19165 29597 19199 29631
rect 20177 29597 20211 29631
rect 20453 29597 20487 29631
rect 22109 29597 22143 29631
rect 7113 29529 7147 29563
rect 23029 29529 23063 29563
rect 1869 29461 1903 29495
rect 3065 29461 3099 29495
rect 3157 29461 3191 29495
rect 4997 29461 5031 29495
rect 5825 29461 5859 29495
rect 8861 29461 8895 29495
rect 13829 29461 13863 29495
rect 22569 29461 22603 29495
rect 26065 29461 26099 29495
rect 27445 29461 27479 29495
rect 29285 29461 29319 29495
rect 31309 29461 31343 29495
rect 1777 29257 1811 29291
rect 3893 29257 3927 29291
rect 4537 29257 4571 29291
rect 7021 29257 7055 29291
rect 10517 29257 10551 29291
rect 11713 29257 11747 29291
rect 12541 29257 12575 29291
rect 19349 29257 19383 29291
rect 19809 29257 19843 29291
rect 22109 29257 22143 29291
rect 27629 29257 27663 29291
rect 1961 29189 1995 29223
rect 11805 29189 11839 29223
rect 18429 29189 18463 29223
rect 2513 29121 2547 29155
rect 6561 29121 6595 29155
rect 8401 29121 8435 29155
rect 10977 29121 11011 29155
rect 12909 29121 12943 29155
rect 13001 29121 13035 29155
rect 14565 29121 14599 29155
rect 14657 29121 14691 29155
rect 17693 29121 17727 29155
rect 17969 29121 18003 29155
rect 26249 29121 26283 29155
rect 28181 29121 28215 29155
rect 30941 29121 30975 29155
rect 3801 29053 3835 29087
rect 4445 29053 4479 29087
rect 5089 29053 5123 29087
rect 5273 29053 5307 29087
rect 5917 29053 5951 29087
rect 6101 29053 6135 29087
rect 6193 29053 6227 29087
rect 6319 29053 6353 29087
rect 10701 29053 10735 29087
rect 10885 29053 10919 29087
rect 11069 29053 11103 29087
rect 11253 29053 11287 29087
rect 11713 29053 11747 29087
rect 12725 29053 12759 29087
rect 13093 29053 13127 29087
rect 13277 29053 13311 29087
rect 14289 29053 14323 29087
rect 14473 29053 14507 29087
rect 14841 29053 14875 29087
rect 15025 29053 15059 29087
rect 15577 29053 15611 29087
rect 18613 29053 18647 29087
rect 21189 29053 21223 29087
rect 23222 29053 23256 29087
rect 23489 29053 23523 29087
rect 24409 29053 24443 29087
rect 28457 29053 28491 29087
rect 1593 28985 1627 29019
rect 1809 28985 1843 29019
rect 2789 28985 2823 29019
rect 5181 28985 5215 29019
rect 8134 28985 8168 29019
rect 9873 28985 9907 29019
rect 11989 28985 12023 29019
rect 20922 28985 20956 29019
rect 24654 28985 24688 29019
rect 26516 28985 26550 29019
rect 30674 28985 30708 29019
rect 2697 28917 2731 28951
rect 3157 28917 3191 28951
rect 9045 28917 9079 28951
rect 16313 28917 16347 28951
rect 25789 28917 25823 28951
rect 29561 28917 29595 28951
rect 4445 28713 4479 28747
rect 5733 28713 5767 28747
rect 11529 28713 11563 28747
rect 14381 28713 14415 28747
rect 16681 28713 16715 28747
rect 19993 28713 20027 28747
rect 21281 28713 21315 28747
rect 23949 28713 23983 28747
rect 26433 28713 26467 28747
rect 28181 28713 28215 28747
rect 1685 28645 1719 28679
rect 13268 28645 13302 28679
rect 15301 28645 15335 28679
rect 1961 28577 1995 28611
rect 2697 28577 2731 28611
rect 3065 28577 3099 28611
rect 3341 28577 3375 28611
rect 4353 28577 4387 28611
rect 5457 28577 5491 28611
rect 6193 28577 6227 28611
rect 6653 28577 6687 28611
rect 6745 28577 6779 28611
rect 6837 28577 6871 28611
rect 7021 28577 7055 28611
rect 7757 28577 7791 28611
rect 9229 28577 9263 28611
rect 9597 28577 9631 28611
rect 9781 28577 9815 28611
rect 10425 28577 10459 28611
rect 10701 28577 10735 28611
rect 10793 28577 10827 28611
rect 10977 28577 11011 28611
rect 11713 28577 11747 28611
rect 12081 28577 12115 28611
rect 12265 28577 12299 28611
rect 15025 28577 15059 28611
rect 15393 28577 15427 28611
rect 15853 28577 15887 28611
rect 16865 28577 16899 28611
rect 17049 28577 17083 28611
rect 17233 28577 17267 28611
rect 17417 28577 17451 28611
rect 18133 28577 18167 28611
rect 20177 28577 20211 28611
rect 20453 28577 20487 28611
rect 20545 28577 20579 28611
rect 20729 28577 20763 28611
rect 23130 28577 23164 28611
rect 23372 28577 23406 28611
rect 24041 28577 24075 28611
rect 24685 28577 24719 28611
rect 24869 28577 24903 28611
rect 25053 28577 25087 28611
rect 25237 28577 25271 28611
rect 1685 28509 1719 28543
rect 3709 28509 3743 28543
rect 5549 28509 5583 28543
rect 5733 28509 5767 28543
rect 25697 28575 25731 28609
rect 25881 28577 25915 28611
rect 26249 28577 26283 28611
rect 27445 28577 27479 28611
rect 27629 28577 27663 28611
rect 27997 28577 28031 28611
rect 28641 28577 28675 28611
rect 28825 28577 28859 28611
rect 29193 28577 29227 28611
rect 29377 28577 29411 28611
rect 30950 28577 30984 28611
rect 31217 28577 31251 28611
rect 6377 28509 6411 28543
rect 8033 28509 8067 28543
rect 9413 28509 9447 28543
rect 9505 28509 9539 28543
rect 10609 28509 10643 28543
rect 11897 28509 11931 28543
rect 11989 28509 12023 28543
rect 13001 28509 13035 28543
rect 14841 28509 14875 28543
rect 17141 28509 17175 28543
rect 17877 28509 17911 28543
rect 20361 28509 20395 28543
rect 24961 28509 24995 28543
rect 25973 28509 26007 28543
rect 26065 28509 26099 28543
rect 27721 28509 27755 28543
rect 27813 28509 27847 28543
rect 28917 28509 28951 28543
rect 29009 28509 29043 28543
rect 3157 28441 3191 28475
rect 6193 28441 6227 28475
rect 1869 28373 1903 28407
rect 9045 28373 9079 28407
rect 10241 28373 10275 28407
rect 15945 28373 15979 28407
rect 19257 28373 19291 28407
rect 22017 28373 22051 28407
rect 24501 28373 24535 28407
rect 29837 28373 29871 28407
rect 1593 28169 1627 28203
rect 3893 28169 3927 28203
rect 4905 28169 4939 28203
rect 7113 28169 7147 28203
rect 10793 28169 10827 28203
rect 14841 28169 14875 28203
rect 23765 28169 23799 28203
rect 30297 28169 30331 28203
rect 3065 28101 3099 28135
rect 6193 28101 6227 28135
rect 20361 28101 20395 28135
rect 2421 28033 2455 28067
rect 7481 28033 7515 28067
rect 7573 28033 7607 28067
rect 13553 28033 13587 28067
rect 14381 28033 14415 28067
rect 15945 28033 15979 28067
rect 17049 28033 17083 28067
rect 22293 28033 22327 28067
rect 24869 28033 24903 28067
rect 27537 28033 27571 28067
rect 1501 27965 1535 27999
rect 2605 27965 2639 27999
rect 2789 27965 2823 27999
rect 3065 27965 3099 27999
rect 3801 27965 3835 27999
rect 4905 27965 4939 27999
rect 5089 27965 5123 27999
rect 5549 27965 5583 27999
rect 5733 27965 5767 27999
rect 5828 27965 5862 27999
rect 5917 27965 5951 27999
rect 7297 27965 7331 27999
rect 7665 27965 7699 27999
rect 7849 27965 7883 27999
rect 9413 27965 9447 27999
rect 9680 27965 9714 27999
rect 14105 27965 14139 27999
rect 14289 27965 14323 27999
rect 14473 27965 14507 27999
rect 14657 27965 14691 27999
rect 16221 27965 16255 27999
rect 17325 27965 17359 27999
rect 18521 27965 18555 27999
rect 19625 27965 19659 27999
rect 19809 27965 19843 27999
rect 20269 27965 20303 27999
rect 21189 27965 21223 27999
rect 21557 27965 21591 27999
rect 22017 27965 22051 27999
rect 23581 27965 23615 27999
rect 25125 27965 25159 27999
rect 27261 27965 27295 27999
rect 28549 27965 28583 27999
rect 29561 27965 29595 27999
rect 29745 27965 29779 27999
rect 29837 27965 29871 27999
rect 29929 27965 29963 27999
rect 30113 27965 30147 27999
rect 31125 27965 31159 27999
rect 11253 27897 11287 27931
rect 13001 27897 13035 27931
rect 22937 27897 22971 27931
rect 8401 27829 8435 27863
rect 18613 27829 18647 27863
rect 23029 27829 23063 27863
rect 26249 27829 26283 27863
rect 26709 27829 26743 27863
rect 28641 27829 28675 27863
rect 31309 27829 31343 27863
rect 2237 27625 2271 27659
rect 14749 27625 14783 27659
rect 19809 27625 19843 27659
rect 21189 27625 21223 27659
rect 24225 27625 24259 27659
rect 31309 27625 31343 27659
rect 1593 27557 1627 27591
rect 5549 27557 5583 27591
rect 6469 27557 6503 27591
rect 8033 27557 8067 27591
rect 8738 27557 8772 27591
rect 10333 27557 10367 27591
rect 14565 27557 14599 27591
rect 18613 27557 18647 27591
rect 23029 27557 23063 27591
rect 24317 27557 24351 27591
rect 27813 27557 27847 27591
rect 1501 27489 1535 27523
rect 2145 27489 2179 27523
rect 2329 27489 2363 27523
rect 3341 27489 3375 27523
rect 3525 27489 3559 27523
rect 3893 27489 3927 27523
rect 4997 27489 5031 27523
rect 5089 27489 5123 27523
rect 5825 27489 5859 27523
rect 6377 27489 6411 27523
rect 6561 27489 6595 27523
rect 7297 27489 7331 27523
rect 7481 27489 7515 27523
rect 7849 27489 7883 27523
rect 8493 27489 8527 27523
rect 11897 27489 11931 27523
rect 12153 27489 12187 27523
rect 14197 27489 14231 27523
rect 15669 27489 15703 27523
rect 16865 27489 16899 27523
rect 17141 27489 17175 27523
rect 17233 27495 17267 27529
rect 17417 27489 17451 27523
rect 17877 27489 17911 27523
rect 18061 27489 18095 27523
rect 18245 27489 18279 27523
rect 18429 27489 18463 27523
rect 19073 27489 19107 27523
rect 19257 27489 19291 27523
rect 19349 27489 19383 27523
rect 19625 27489 19659 27523
rect 20453 27489 20487 27523
rect 20637 27489 20671 27523
rect 21005 27489 21039 27523
rect 22293 27489 22327 27523
rect 23397 27489 23431 27523
rect 25881 27489 25915 27523
rect 27629 27489 27663 27523
rect 28825 27489 28859 27523
rect 29561 27489 29595 27523
rect 29745 27489 29779 27523
rect 30113 27489 30147 27523
rect 31125 27489 31159 27523
rect 2881 27421 2915 27455
rect 3617 27421 3651 27455
rect 3709 27421 3743 27455
rect 5549 27421 5583 27455
rect 7573 27421 7607 27455
rect 7665 27421 7699 27455
rect 15945 27421 15979 27455
rect 17049 27421 17083 27455
rect 18153 27421 18187 27455
rect 19441 27421 19475 27455
rect 20729 27421 20763 27455
rect 20821 27421 20855 27455
rect 26157 27421 26191 27455
rect 29101 27421 29135 27455
rect 29837 27421 29871 27455
rect 29929 27421 29963 27455
rect 26985 27353 27019 27387
rect 4077 27285 4111 27319
rect 5733 27285 5767 27319
rect 9873 27285 9907 27319
rect 10977 27285 11011 27319
rect 13277 27285 13311 27319
rect 14565 27285 14599 27319
rect 16681 27285 16715 27319
rect 22477 27285 22511 27319
rect 30297 27285 30331 27319
rect 1777 27081 1811 27115
rect 6285 27081 6319 27115
rect 10333 27081 10367 27115
rect 11989 27081 12023 27115
rect 15301 27081 15335 27115
rect 17141 27081 17175 27115
rect 19625 27081 19659 27115
rect 19809 27081 19843 27115
rect 20729 27081 20763 27115
rect 20913 27081 20947 27115
rect 24593 27081 24627 27115
rect 25605 27081 25639 27115
rect 27629 27081 27663 27115
rect 11529 26945 11563 26979
rect 13185 26945 13219 26979
rect 2421 26877 2455 26911
rect 3801 26877 3835 26911
rect 3985 26877 4019 26911
rect 4077 26877 4111 26911
rect 4169 26877 4203 26911
rect 4353 26877 4387 26911
rect 5181 26877 5215 26911
rect 8309 26877 8343 26911
rect 8953 26877 8987 26911
rect 11253 26877 11287 26911
rect 11437 26877 11471 26911
rect 11621 26877 11655 26911
rect 11805 26877 11839 26911
rect 12817 26877 12851 26911
rect 13001 26877 13035 26911
rect 13093 26877 13127 26911
rect 13369 26877 13403 26911
rect 13553 26877 13587 26911
rect 14749 26877 14783 26911
rect 16681 26877 16715 26911
rect 4997 26809 5031 26843
rect 7573 26809 7607 26843
rect 9220 26809 9254 26843
rect 16414 26809 16448 26843
rect 19257 27013 19291 27047
rect 20361 27013 20395 27047
rect 23213 27013 23247 27047
rect 17601 26945 17635 26979
rect 21741 26945 21775 26979
rect 31217 26945 31251 26979
rect 17233 26877 17267 26911
rect 17417 26877 17451 26911
rect 17509 26877 17543 26911
rect 17785 26877 17819 26911
rect 18613 26877 18647 26911
rect 22569 26877 22603 26911
rect 22753 26877 22787 26911
rect 23213 26877 23247 26911
rect 24961 26877 24995 26911
rect 26525 26877 26559 26911
rect 26985 26877 27019 26911
rect 27169 26877 27203 26911
rect 28365 26877 28399 26911
rect 29009 26877 29043 26911
rect 30950 26877 30984 26911
rect 19625 26809 19659 26843
rect 20729 26809 20763 26843
rect 21465 26809 21499 26843
rect 25513 26809 25547 26843
rect 27077 26809 27111 26843
rect 2513 26741 2547 26775
rect 3249 26741 3283 26775
rect 4537 26741 4571 26775
rect 14565 26741 14599 26775
rect 17141 26741 17175 26775
rect 17969 26741 18003 26775
rect 18521 26741 18555 26775
rect 24409 26741 24443 26775
rect 24593 26741 24627 26775
rect 26433 26741 26467 26775
rect 28273 26741 28307 26775
rect 28917 26741 28951 26775
rect 29837 26741 29871 26775
rect 3433 26537 3467 26571
rect 5733 26537 5767 26571
rect 10977 26537 11011 26571
rect 15853 26537 15887 26571
rect 18705 26537 18739 26571
rect 22937 26537 22971 26571
rect 28917 26537 28951 26571
rect 4546 26469 4580 26503
rect 16129 26469 16163 26503
rect 19625 26469 19659 26503
rect 23765 26469 23799 26503
rect 28457 26469 28491 26503
rect 2053 26401 2087 26435
rect 2237 26401 2271 26435
rect 2421 26401 2455 26435
rect 2605 26401 2639 26435
rect 5825 26401 5859 26435
rect 6745 26401 6779 26435
rect 7001 26401 7035 26435
rect 8585 26401 8619 26435
rect 8769 26401 8803 26435
rect 8953 26401 8987 26435
rect 9137 26401 9171 26435
rect 11529 26401 11563 26435
rect 11713 26401 11747 26435
rect 11897 26401 11931 26435
rect 12081 26401 12115 26435
rect 12725 26401 12759 26435
rect 13553 26401 13587 26435
rect 13737 26401 13771 26435
rect 14289 26401 14323 26435
rect 15025 26401 15059 26435
rect 15853 26401 15887 26435
rect 17141 26401 17175 26435
rect 17601 26401 17635 26435
rect 17877 26401 17911 26435
rect 18521 26401 18555 26435
rect 19257 26401 19291 26435
rect 20269 26401 20303 26435
rect 20453 26401 20487 26435
rect 20545 26401 20579 26435
rect 20821 26401 20855 26435
rect 22201 26401 22235 26435
rect 22385 26401 22419 26435
rect 22753 26401 22787 26435
rect 23397 26401 23431 26435
rect 23581 26401 23615 26435
rect 24593 26401 24627 26435
rect 24869 26401 24903 26435
rect 25881 26401 25915 26435
rect 26985 26401 27019 26435
rect 27721 26401 27755 26435
rect 27905 26401 27939 26435
rect 28273 26401 28307 26435
rect 29469 26401 29503 26435
rect 29653 26401 29687 26435
rect 30021 26401 30055 26435
rect 30849 26401 30883 26435
rect 1593 26333 1627 26367
rect 2329 26333 2363 26367
rect 4813 26333 4847 26367
rect 8861 26333 8895 26367
rect 11805 26333 11839 26367
rect 16957 26333 16991 26367
rect 20637 26333 20671 26367
rect 22477 26333 22511 26367
rect 22569 26333 22603 26367
rect 25237 26333 25271 26367
rect 27997 26333 28031 26367
rect 28089 26333 28123 26367
rect 29745 26333 29779 26367
rect 29837 26333 29871 26367
rect 30757 26333 30791 26367
rect 2789 26265 2823 26299
rect 9781 26265 9815 26299
rect 10425 26265 10459 26299
rect 12265 26265 12299 26299
rect 12817 26265 12851 26299
rect 14197 26265 14231 26299
rect 15945 26265 15979 26299
rect 19809 26265 19843 26299
rect 24593 26265 24627 26299
rect 27077 26265 27111 26299
rect 30205 26265 30239 26299
rect 8125 26197 8159 26231
rect 9321 26197 9355 26231
rect 15117 26197 15151 26231
rect 19625 26197 19659 26231
rect 21005 26197 21039 26231
rect 25881 26197 25915 26231
rect 1409 25993 1443 26027
rect 5181 25993 5215 26027
rect 6837 25993 6871 26027
rect 8217 25993 8251 26027
rect 14197 25993 14231 26027
rect 15025 25993 15059 26027
rect 16129 25993 16163 26027
rect 17877 25993 17911 26027
rect 19717 25993 19751 26027
rect 21557 25993 21591 26027
rect 22477 25993 22511 26027
rect 22661 25993 22695 26027
rect 27721 25993 27755 26027
rect 11621 25925 11655 25959
rect 23213 25925 23247 25959
rect 28181 25925 28215 25959
rect 7297 25857 7331 25891
rect 9045 25857 9079 25891
rect 18245 25857 18279 25891
rect 18337 25857 18371 25891
rect 21097 25857 21131 25891
rect 25421 25857 25455 25891
rect 26801 25857 26835 25891
rect 26893 25857 26927 25891
rect 2522 25789 2556 25823
rect 2789 25789 2823 25823
rect 3801 25789 3835 25823
rect 7021 25789 7055 25823
rect 7205 25789 7239 25823
rect 7389 25789 7423 25823
rect 7573 25789 7607 25823
rect 8033 25789 8067 25823
rect 9312 25789 9346 25823
rect 12734 25789 12768 25823
rect 13001 25789 13035 25823
rect 14657 25789 14691 25823
rect 18061 25789 18095 25823
rect 18429 25789 18463 25823
rect 18613 25789 18647 25823
rect 22109 25789 22143 25823
rect 23121 25789 23155 25823
rect 24593 25789 24627 25823
rect 24685 25789 24719 25823
rect 25513 25789 25547 25823
rect 25605 25789 25639 25823
rect 26617 25789 26651 25823
rect 26985 25789 27019 25823
rect 27169 25789 27203 25823
rect 27905 25789 27939 25823
rect 27997 25789 28031 25823
rect 28273 25789 28307 25823
rect 28917 25789 28951 25823
rect 31042 25789 31076 25823
rect 31309 25789 31343 25823
rect 4068 25721 4102 25755
rect 15025 25721 15059 25755
rect 17417 25721 17451 25755
rect 20830 25721 20864 25755
rect 22477 25721 22511 25755
rect 28825 25721 28859 25755
rect 5641 25653 5675 25687
rect 6377 25653 6411 25687
rect 10425 25653 10459 25687
rect 11069 25653 11103 25687
rect 13461 25653 13495 25687
rect 15209 25653 15243 25687
rect 23857 25653 23891 25687
rect 24409 25653 24443 25687
rect 25973 25653 26007 25687
rect 26433 25653 26467 25687
rect 29929 25653 29963 25687
rect 1593 25449 1627 25483
rect 3709 25449 3743 25483
rect 6837 25449 6871 25483
rect 13369 25449 13403 25483
rect 16865 25449 16899 25483
rect 18889 25449 18923 25483
rect 23029 25449 23063 25483
rect 24501 25449 24535 25483
rect 26223 25449 26257 25483
rect 31309 25449 31343 25483
rect 9505 25381 9539 25415
rect 9689 25381 9723 25415
rect 10701 25381 10735 25415
rect 13185 25381 13219 25415
rect 13829 25381 13863 25415
rect 17776 25381 17810 25415
rect 25228 25381 25262 25415
rect 26433 25381 26467 25415
rect 30573 25381 30607 25415
rect 1409 25313 1443 25347
rect 6837 25313 6871 25347
rect 8033 25313 8067 25347
rect 8309 25313 8343 25347
rect 8769 25313 8803 25347
rect 8953 25313 8987 25347
rect 10885 25313 10919 25347
rect 12817 25313 12851 25347
rect 14013 25313 14047 25347
rect 14197 25313 14231 25347
rect 14381 25313 14415 25347
rect 14565 25313 14599 25347
rect 15025 25313 15059 25347
rect 15393 25313 15427 25347
rect 15853 25313 15887 25347
rect 16681 25313 16715 25347
rect 17509 25313 17543 25347
rect 20462 25313 20496 25347
rect 21833 25313 21867 25347
rect 22017 25313 22051 25347
rect 22385 25313 22419 25347
rect 23029 25313 23063 25347
rect 23121 25313 23155 25347
rect 23388 25313 23422 25347
rect 24961 25313 24995 25347
rect 25605 25313 25639 25347
rect 26985 25313 27019 25347
rect 27261 25313 27295 25347
rect 27353 25313 27387 25347
rect 29285 25313 29319 25347
rect 29469 25313 29503 25347
rect 29561 25313 29595 25347
rect 29837 25313 29871 25347
rect 30481 25313 30515 25347
rect 31125 25313 31159 25347
rect 2329 25245 2363 25279
rect 2421 25245 2455 25279
rect 2697 25245 2731 25279
rect 12081 25245 12115 25279
rect 12357 25245 12391 25279
rect 14289 25245 14323 25279
rect 20729 25245 20763 25279
rect 27997 25245 28031 25279
rect 28273 25245 28307 25279
rect 29653 25245 29687 25279
rect 5181 25177 5215 25211
rect 8953 25177 8987 25211
rect 15945 25177 15979 25211
rect 19349 25177 19383 25211
rect 26065 25177 26099 25211
rect 2329 25109 2363 25143
rect 4629 25109 4663 25143
rect 5733 25109 5767 25143
rect 13185 25109 13219 25143
rect 21189 25109 21223 25143
rect 22293 25109 22327 25143
rect 25237 25109 25271 25143
rect 26249 25109 26283 25143
rect 27077 25109 27111 25143
rect 27537 25109 27571 25143
rect 30021 25109 30055 25143
rect 16129 24905 16163 24939
rect 23765 24905 23799 24939
rect 24409 24905 24443 24939
rect 23213 24837 23247 24871
rect 2789 24769 2823 24803
rect 4997 24769 5031 24803
rect 7113 24769 7147 24803
rect 8125 24769 8159 24803
rect 9689 24769 9723 24803
rect 11069 24769 11103 24803
rect 12633 24769 12667 24803
rect 19717 24769 19751 24803
rect 20085 24769 20119 24803
rect 20637 24769 20671 24803
rect 22661 24769 22695 24803
rect 25145 24769 25179 24803
rect 25421 24769 25455 24803
rect 25513 24769 25547 24803
rect 26249 24769 26283 24803
rect 26525 24769 26559 24803
rect 26709 24769 26743 24803
rect 27905 24769 27939 24803
rect 27997 24769 28031 24803
rect 30941 24769 30975 24803
rect 3801 24701 3835 24735
rect 3985 24701 4019 24735
rect 4077 24701 4111 24735
rect 4169 24701 4203 24735
rect 4353 24701 4387 24735
rect 6837 24701 6871 24735
rect 8309 24701 8343 24735
rect 8953 24701 8987 24735
rect 9781 24701 9815 24735
rect 10793 24701 10827 24735
rect 10977 24701 11011 24735
rect 11161 24701 11195 24735
rect 11345 24701 11379 24735
rect 12357 24701 12391 24735
rect 12541 24701 12575 24735
rect 12725 24701 12759 24735
rect 12909 24701 12943 24735
rect 14105 24701 14139 24735
rect 18705 24701 18739 24735
rect 19349 24701 19383 24735
rect 19533 24701 19567 24735
rect 19625 24701 19659 24735
rect 19901 24701 19935 24735
rect 20729 24701 20763 24735
rect 22394 24701 22428 24735
rect 23305 24701 23339 24735
rect 24593 24701 24627 24735
rect 25053 24701 25087 24735
rect 25329 24701 25363 24735
rect 25605 24701 25639 24735
rect 25789 24701 25823 24735
rect 26433 24701 26467 24735
rect 26617 24701 26651 24735
rect 26893 24701 26927 24735
rect 27629 24701 27663 24735
rect 27813 24701 27847 24735
rect 28181 24701 28215 24735
rect 28917 24701 28951 24735
rect 29009 24701 29043 24735
rect 30674 24701 30708 24735
rect 2522 24633 2556 24667
rect 5242 24633 5276 24667
rect 14372 24633 14406 24667
rect 16037 24633 16071 24667
rect 17049 24633 17083 24667
rect 1409 24565 1443 24599
rect 4537 24565 4571 24599
rect 6377 24565 6411 24599
rect 9045 24565 9079 24599
rect 10333 24565 10367 24599
rect 11529 24565 11563 24599
rect 13093 24565 13127 24599
rect 15485 24565 15519 24599
rect 21281 24565 21315 24599
rect 25053 24565 25087 24599
rect 28365 24565 28399 24599
rect 29561 24565 29595 24599
rect 2605 24361 2639 24395
rect 5089 24361 5123 24395
rect 10793 24361 10827 24395
rect 16037 24361 16071 24395
rect 18705 24361 18739 24395
rect 21281 24361 21315 24395
rect 21925 24361 21959 24395
rect 23949 24361 23983 24395
rect 27353 24361 27387 24395
rect 28181 24361 28215 24395
rect 28825 24361 28859 24395
rect 29929 24361 29963 24395
rect 30573 24361 30607 24395
rect 15393 24293 15427 24327
rect 26985 24293 27019 24327
rect 27169 24293 27203 24327
rect 29377 24293 29411 24327
rect 1869 24225 1903 24259
rect 2053 24225 2087 24259
rect 2421 24225 2455 24259
rect 5273 24225 5307 24259
rect 5457 24225 5491 24259
rect 5641 24225 5675 24259
rect 5825 24225 5859 24259
rect 7685 24225 7719 24259
rect 7941 24225 7975 24259
rect 8953 24225 8987 24259
rect 9045 24225 9079 24259
rect 9137 24225 9171 24259
rect 9321 24225 9355 24259
rect 9781 24225 9815 24259
rect 9965 24225 9999 24259
rect 10885 24225 10919 24259
rect 11529 24225 11563 24259
rect 13001 24225 13035 24259
rect 13185 24225 13219 24259
rect 13737 24225 13771 24259
rect 14381 24225 14415 24259
rect 17233 24225 17267 24259
rect 17969 24225 18003 24259
rect 18153 24225 18187 24259
rect 18245 24225 18279 24259
rect 18521 24225 18555 24259
rect 19441 24225 19475 24259
rect 19809 24225 19843 24259
rect 20545 24225 20579 24259
rect 20729 24225 20763 24259
rect 20913 24225 20947 24259
rect 21097 24225 21131 24259
rect 22385 24225 22419 24259
rect 22569 24225 22603 24259
rect 22937 24225 22971 24259
rect 24869 24225 24903 24259
rect 26249 24225 26283 24259
rect 26433 24225 26467 24259
rect 28273 24225 28307 24259
rect 28917 24225 28951 24259
rect 31125 24225 31159 24259
rect 2145 24157 2179 24191
rect 2237 24157 2271 24191
rect 3893 24157 3927 24191
rect 4169 24157 4203 24191
rect 5549 24157 5583 24191
rect 8677 24157 8711 24191
rect 14657 24157 14691 24191
rect 15577 24157 15611 24191
rect 17509 24157 17543 24191
rect 18337 24157 18371 24191
rect 19257 24157 19291 24191
rect 20830 24157 20864 24191
rect 22661 24157 22695 24191
rect 22753 24157 22787 24191
rect 23121 24157 23155 24191
rect 25513 24157 25547 24191
rect 13645 24089 13679 24123
rect 19717 24089 19751 24123
rect 23581 24089 23615 24123
rect 6561 24021 6595 24055
rect 9965 24021 9999 24055
rect 11759 24021 11793 24055
rect 23949 24021 23983 24055
rect 24133 24021 24167 24055
rect 26065 24021 26099 24055
rect 26341 24021 26375 24055
rect 31309 24021 31343 24055
rect 3801 23817 3835 23851
rect 8125 23817 8159 23851
rect 12817 23817 12851 23851
rect 13001 23817 13035 23851
rect 13461 23817 13495 23851
rect 16129 23817 16163 23851
rect 18705 23817 18739 23851
rect 19441 23817 19475 23851
rect 19625 23817 19659 23851
rect 23489 23817 23523 23851
rect 24869 23817 24903 23851
rect 27445 23817 27479 23851
rect 12449 23749 12483 23783
rect 17049 23749 17083 23783
rect 21557 23749 21591 23783
rect 25789 23749 25823 23783
rect 7665 23681 7699 23715
rect 7757 23681 7791 23715
rect 14841 23681 14875 23715
rect 19993 23681 20027 23715
rect 24409 23681 24443 23715
rect 1869 23613 1903 23647
rect 4914 23613 4948 23647
rect 5181 23613 5215 23647
rect 6101 23613 6135 23647
rect 6377 23613 6411 23647
rect 7389 23613 7423 23647
rect 7573 23613 7607 23647
rect 7941 23613 7975 23647
rect 9229 23613 9263 23647
rect 9321 23613 9355 23647
rect 9413 23613 9447 23647
rect 9597 23613 9631 23647
rect 11722 23613 11756 23647
rect 11989 23613 12023 23647
rect 14657 23613 14691 23647
rect 14939 23613 14973 23647
rect 15037 23613 15071 23647
rect 15209 23613 15243 23647
rect 15945 23613 15979 23647
rect 16037 23613 16071 23647
rect 16221 23613 16255 23647
rect 17969 23613 18003 23647
rect 18153 23613 18187 23647
rect 18245 23613 18279 23647
rect 18337 23613 18371 23647
rect 18521 23613 18555 23647
rect 20729 23613 20763 23647
rect 22937 23613 22971 23647
rect 23581 23613 23615 23647
rect 24593 23613 24627 23647
rect 24961 23613 24995 23647
rect 26249 23613 26283 23647
rect 26433 23613 26467 23647
rect 28181 23613 28215 23647
rect 28365 23613 28399 23647
rect 28460 23613 28494 23647
rect 28549 23613 28583 23647
rect 28733 23613 28767 23647
rect 30941 23613 30975 23647
rect 10149 23545 10183 23579
rect 16773 23545 16807 23579
rect 20545 23545 20579 23579
rect 22670 23545 22704 23579
rect 25421 23545 25455 23579
rect 25605 23545 25639 23579
rect 27077 23545 27111 23579
rect 27261 23545 27295 23579
rect 28917 23545 28951 23579
rect 30674 23545 30708 23579
rect 1961 23477 1995 23511
rect 2789 23477 2823 23511
rect 8953 23477 8987 23511
rect 10609 23477 10643 23511
rect 12817 23477 12851 23511
rect 14473 23477 14507 23511
rect 19625 23477 19659 23511
rect 26617 23477 26651 23511
rect 29561 23477 29595 23511
rect 3249 23273 3283 23307
rect 3893 23273 3927 23307
rect 7665 23273 7699 23307
rect 18889 23273 18923 23307
rect 19993 23273 20027 23307
rect 22569 23273 22603 23307
rect 24961 23273 24995 23307
rect 26433 23273 26467 23307
rect 30297 23273 30331 23307
rect 31309 23273 31343 23307
rect 17601 23205 17635 23239
rect 29101 23205 29135 23239
rect 29745 23205 29779 23239
rect 2136 23137 2170 23171
rect 4353 23137 4387 23171
rect 4609 23137 4643 23171
rect 6377 23137 6411 23171
rect 6561 23137 6595 23171
rect 6745 23137 6779 23171
rect 6929 23137 6963 23171
rect 7757 23137 7791 23171
rect 8309 23137 8343 23171
rect 9321 23137 9355 23171
rect 9965 23137 9999 23171
rect 11529 23137 11563 23171
rect 12633 23137 12667 23171
rect 12909 23137 12943 23171
rect 13553 23137 13587 23171
rect 13820 23137 13854 23171
rect 15393 23137 15427 23171
rect 15577 23137 15611 23171
rect 15761 23137 15795 23171
rect 15945 23137 15979 23171
rect 17049 23137 17083 23171
rect 19901 23137 19935 23171
rect 20545 23137 20579 23171
rect 20729 23137 20763 23171
rect 20821 23137 20855 23171
rect 20913 23137 20947 23171
rect 21097 23137 21131 23171
rect 21281 23137 21315 23171
rect 21833 23137 21867 23171
rect 22017 23137 22051 23171
rect 22201 23137 22235 23171
rect 22385 23137 22419 23171
rect 23848 23137 23882 23171
rect 25881 23137 25915 23171
rect 27537 23137 27571 23171
rect 27629 23137 27663 23171
rect 27905 23137 27939 23171
rect 28457 23137 28491 23171
rect 28549 23137 28583 23171
rect 29009 23137 29043 23171
rect 31125 23137 31159 23171
rect 1869 23069 1903 23103
rect 6653 23069 6687 23103
rect 8401 23069 8435 23103
rect 8585 23069 8619 23103
rect 9597 23069 9631 23103
rect 10333 23069 10367 23103
rect 11621 23069 11655 23103
rect 15669 23069 15703 23103
rect 22109 23069 22143 23103
rect 23581 23069 23615 23103
rect 26157 23069 26191 23103
rect 8493 23001 8527 23035
rect 9781 23001 9815 23035
rect 27813 23001 27847 23035
rect 5733 22933 5767 22967
rect 7113 22933 7147 22967
rect 14933 22933 14967 22967
rect 16129 22933 16163 22967
rect 16957 22933 16991 22967
rect 23029 22933 23063 22967
rect 26065 22933 26099 22967
rect 27353 22933 27387 22967
rect 2605 22729 2639 22763
rect 5917 22729 5951 22763
rect 8309 22729 8343 22763
rect 10057 22729 10091 22763
rect 19625 22729 19659 22763
rect 23121 22729 23155 22763
rect 23857 22729 23891 22763
rect 24409 22729 24443 22763
rect 26525 22729 26559 22763
rect 29561 22661 29595 22695
rect 2237 22593 2271 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 8401 22593 8435 22627
rect 9505 22593 9539 22627
rect 9597 22593 9631 22627
rect 10885 22593 10919 22627
rect 14749 22593 14783 22627
rect 21005 22593 21039 22627
rect 21741 22593 21775 22627
rect 26985 22593 27019 22627
rect 28457 22593 28491 22627
rect 28549 22593 28583 22627
rect 30941 22593 30975 22627
rect 1857 22515 1891 22549
rect 2057 22525 2091 22559
rect 2154 22525 2188 22559
rect 2421 22525 2455 22559
rect 3985 22525 4019 22559
rect 4629 22525 4663 22559
rect 6837 22525 6871 22559
rect 7021 22525 7055 22559
rect 7389 22525 7423 22559
rect 8125 22525 8159 22559
rect 8217 22525 8251 22559
rect 9689 22525 9723 22559
rect 10609 22525 10643 22559
rect 10793 22525 10827 22559
rect 10977 22525 11011 22559
rect 11161 22525 11195 22559
rect 11805 22525 11839 22559
rect 14473 22525 14507 22559
rect 15761 22525 15795 22559
rect 16028 22525 16062 22559
rect 17601 22525 17635 22559
rect 17969 22525 18003 22559
rect 18429 22525 18463 22559
rect 25789 22525 25823 22559
rect 26709 22525 26743 22559
rect 26893 22525 26927 22559
rect 27077 22525 27111 22559
rect 27261 22525 27295 22559
rect 28181 22525 28215 22559
rect 28365 22525 28399 22559
rect 28733 22525 28767 22559
rect 3249 22457 3283 22491
rect 11345 22457 11379 22491
rect 12050 22457 12084 22491
rect 18705 22457 18739 22491
rect 20738 22457 20772 22491
rect 21986 22457 22020 22491
rect 25522 22457 25556 22491
rect 28917 22457 28951 22491
rect 30674 22457 30708 22491
rect 3893 22389 3927 22423
rect 7573 22389 7607 22423
rect 13185 22389 13219 22423
rect 17141 22389 17175 22423
rect 21005 22185 21039 22219
rect 23489 22185 23523 22219
rect 25145 22185 25179 22219
rect 26433 22185 26467 22219
rect 27077 22185 27111 22219
rect 22201 22117 22235 22151
rect 26065 22117 26099 22151
rect 26249 22117 26283 22151
rect 1409 22049 1443 22083
rect 1676 22049 1710 22083
rect 3249 22049 3283 22083
rect 3433 22049 3467 22083
rect 3617 22049 3651 22083
rect 3801 22049 3835 22083
rect 3985 22049 4019 22083
rect 5558 22049 5592 22083
rect 5825 22049 5859 22083
rect 6828 22049 6862 22083
rect 9045 22049 9079 22083
rect 9229 22049 9263 22083
rect 9597 22049 9631 22083
rect 10241 22049 10275 22083
rect 10425 22049 10459 22083
rect 10793 22049 10827 22083
rect 10977 22049 11011 22083
rect 11785 22049 11819 22083
rect 13369 22049 13403 22083
rect 13461 22049 13495 22083
rect 14657 22049 14691 22083
rect 15945 22049 15979 22083
rect 16773 22049 16807 22083
rect 16957 22049 16991 22083
rect 17049 22049 17083 22083
rect 17325 22049 17359 22083
rect 17509 22049 17543 22083
rect 18429 22049 18463 22083
rect 18613 22049 18647 22083
rect 18981 22049 19015 22083
rect 19892 22049 19926 22083
rect 24409 22049 24443 22083
rect 24593 22049 24627 22083
rect 24961 22049 24995 22083
rect 26985 22049 27019 22083
rect 28089 22049 28123 22083
rect 28273 22047 28307 22081
rect 28457 22049 28491 22083
rect 28641 22049 28675 22083
rect 29285 22049 29319 22083
rect 29377 22049 29411 22083
rect 30481 22049 30515 22083
rect 31309 22049 31343 22083
rect 3709 21981 3743 22015
rect 6561 21981 6595 22015
rect 8861 21981 8895 22015
rect 9413 21981 9447 22015
rect 10517 21981 10551 22015
rect 10609 21981 10643 22015
rect 11529 21981 11563 22015
rect 15669 21981 15703 22015
rect 17141 21981 17175 22015
rect 18705 21981 18739 22015
rect 18797 21981 18831 22015
rect 19625 21981 19659 22015
rect 24685 21981 24719 22015
rect 24777 21981 24811 22015
rect 28365 21981 28399 22015
rect 14565 21913 14599 21947
rect 30665 21913 30699 21947
rect 2789 21845 2823 21879
rect 4445 21845 4479 21879
rect 7941 21845 7975 21879
rect 12909 21845 12943 21879
rect 19165 21845 19199 21879
rect 28825 21845 28859 21879
rect 29929 21845 29963 21879
rect 31125 21845 31159 21879
rect 1593 21641 1627 21675
rect 4721 21641 4755 21675
rect 5273 21641 5307 21675
rect 9229 21641 9263 21675
rect 14473 21641 14507 21675
rect 17785 21641 17819 21675
rect 18429 21641 18463 21675
rect 19441 21641 19475 21675
rect 21281 21641 21315 21675
rect 22293 21641 22327 21675
rect 23121 21641 23155 21675
rect 24409 21641 24443 21675
rect 9413 21573 9447 21607
rect 23765 21573 23799 21607
rect 31125 21573 31159 21607
rect 1961 21505 1995 21539
rect 5641 21505 5675 21539
rect 5733 21505 5767 21539
rect 7021 21505 7055 21539
rect 9965 21505 9999 21539
rect 14933 21505 14967 21539
rect 19809 21505 19843 21539
rect 19901 21505 19935 21539
rect 24777 21505 24811 21539
rect 25973 21505 26007 21539
rect 27169 21505 27203 21539
rect 27261 21505 27295 21539
rect 28365 21505 28399 21539
rect 30481 21505 30515 21539
rect 1777 21437 1811 21471
rect 2053 21437 2087 21471
rect 2145 21437 2179 21471
rect 2329 21437 2363 21471
rect 5457 21437 5491 21471
rect 5825 21437 5859 21471
rect 6009 21437 6043 21471
rect 7288 21437 7322 21471
rect 10241 21437 10275 21471
rect 11253 21437 11287 21471
rect 11529 21437 11563 21471
rect 13001 21437 13035 21471
rect 13185 21437 13219 21471
rect 13553 21437 13587 21471
rect 14657 21437 14691 21471
rect 14841 21437 14875 21471
rect 15021 21437 15055 21471
rect 15209 21439 15243 21473
rect 15761 21437 15795 21471
rect 17877 21437 17911 21471
rect 19625 21437 19659 21471
rect 19993 21437 20027 21471
rect 20177 21415 20211 21449
rect 23213 21437 23247 21471
rect 23673 21437 23707 21471
rect 24593 21437 24627 21471
rect 24869 21437 24903 21471
rect 24961 21437 24995 21471
rect 25145 21437 25179 21471
rect 25605 21437 25639 21471
rect 25789 21431 25823 21465
rect 25881 21437 25915 21471
rect 26157 21437 26191 21471
rect 26985 21437 27019 21471
rect 27353 21437 27387 21471
rect 27537 21437 27571 21471
rect 28181 21437 28215 21471
rect 28457 21437 28491 21471
rect 28549 21437 28583 21471
rect 28733 21437 28767 21471
rect 30573 21437 30607 21471
rect 31033 21437 31067 21471
rect 31309 21437 31343 21471
rect 9045 21369 9079 21403
rect 9261 21369 9295 21403
rect 13461 21369 13495 21403
rect 16028 21369 16062 21403
rect 18521 21369 18555 21403
rect 30297 21369 30331 21403
rect 3157 21301 3191 21335
rect 4261 21301 4295 21335
rect 6561 21301 6595 21335
rect 8401 21301 8435 21335
rect 17141 21301 17175 21335
rect 20729 21301 20763 21335
rect 26341 21301 26375 21335
rect 26801 21301 26835 21335
rect 27997 21301 28031 21335
rect 29561 21301 29595 21335
rect 30573 21301 30607 21335
rect 31033 21301 31067 21335
rect 5641 21097 5675 21131
rect 8953 21097 8987 21131
rect 9597 21097 9631 21131
rect 12909 21097 12943 21131
rect 16773 21097 16807 21131
rect 28641 21097 28675 21131
rect 30757 21097 30791 21131
rect 3617 21029 3651 21063
rect 3817 21029 3851 21063
rect 5733 21029 5767 21063
rect 10885 21029 10919 21063
rect 22017 21029 22051 21063
rect 22109 21029 22143 21063
rect 29754 21029 29788 21063
rect 1409 20961 1443 20995
rect 2237 20961 2271 20995
rect 2881 20961 2915 20995
rect 4629 20961 4663 20995
rect 7205 20961 7239 20995
rect 8217 20961 8251 20995
rect 8401 20961 8435 20995
rect 9689 20961 9723 20995
rect 10801 20961 10835 20995
rect 11529 20961 11563 20995
rect 11713 20961 11747 20995
rect 11805 20961 11839 20995
rect 12081 20961 12115 20995
rect 13093 20961 13127 20995
rect 13277 20961 13311 20995
rect 13461 20961 13495 20995
rect 13645 20961 13679 20995
rect 14289 20961 14323 20995
rect 14473 20961 14507 20995
rect 14565 20961 14599 20995
rect 14657 20961 14691 20995
rect 14841 20961 14875 20995
rect 16681 20961 16715 20995
rect 17969 20961 18003 20995
rect 18981 20961 19015 20995
rect 22385 20961 22419 20995
rect 23213 20961 23247 20995
rect 23469 20961 23503 20995
rect 25881 20961 25915 20995
rect 27905 20961 27939 20995
rect 31033 20961 31067 20995
rect 31217 20961 31251 20995
rect 3157 20893 3191 20927
rect 6469 20893 6503 20927
rect 6929 20893 6963 20927
rect 11897 20893 11931 20927
rect 13369 20893 13403 20927
rect 15853 20893 15887 20927
rect 16129 20893 16163 20927
rect 18245 20893 18279 20927
rect 18705 20893 18739 20927
rect 19993 20893 20027 20927
rect 20269 20893 20303 20927
rect 22477 20893 22511 20927
rect 25605 20893 25639 20927
rect 28181 20893 28215 20927
rect 30021 20893 30055 20927
rect 30941 20893 30975 20927
rect 31125 20893 31159 20927
rect 1593 20825 1627 20859
rect 3065 20825 3099 20859
rect 2329 20757 2363 20791
rect 2973 20757 3007 20791
rect 3801 20757 3835 20791
rect 3985 20757 4019 20791
rect 4537 20757 4571 20791
rect 10333 20757 10367 20791
rect 12265 20757 12299 20791
rect 14105 20757 14139 20791
rect 24593 20757 24627 20791
rect 25145 20757 25179 20791
rect 13185 20553 13219 20587
rect 13369 20553 13403 20587
rect 16681 20553 16715 20587
rect 22477 20553 22511 20587
rect 23121 20553 23155 20587
rect 25513 20553 25547 20587
rect 28733 20553 28767 20587
rect 30941 20553 30975 20587
rect 3157 20485 3191 20519
rect 5273 20485 5307 20519
rect 2973 20417 3007 20451
rect 4445 20417 4479 20451
rect 8217 20417 8251 20451
rect 11897 20417 11931 20451
rect 16221 20417 16255 20451
rect 19533 20417 19567 20451
rect 20821 20417 20855 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 23572 20417 23606 20451
rect 30481 20417 30515 20451
rect 30665 20417 30699 20451
rect 2329 20349 2363 20383
rect 2513 20349 2547 20383
rect 3249 20349 3283 20383
rect 4261 20349 4295 20383
rect 4537 20349 4571 20383
rect 4905 20349 4939 20383
rect 5917 20349 5951 20383
rect 6377 20349 6411 20383
rect 7021 20349 7055 20383
rect 7941 20349 7975 20383
rect 8033 20349 8067 20383
rect 8953 20349 8987 20383
rect 10977 20349 11011 20383
rect 11621 20349 11655 20383
rect 11805 20349 11839 20383
rect 11985 20349 12019 20383
rect 12173 20349 12207 20383
rect 12817 20349 12851 20383
rect 14105 20349 14139 20383
rect 15945 20349 15979 20383
rect 16129 20349 16163 20383
rect 16313 20349 16347 20383
rect 16497 20349 16531 20383
rect 18245 20349 18279 20383
rect 18521 20349 18555 20383
rect 19257 20349 19291 20383
rect 20545 20349 20579 20383
rect 20729 20349 20763 20383
rect 20913 20349 20947 20383
rect 21097 20349 21131 20383
rect 21741 20349 21775 20383
rect 21925 20349 21959 20383
rect 22293 20349 22327 20383
rect 23305 20349 23339 20383
rect 23489 20349 23523 20383
rect 23673 20349 23707 20383
rect 23857 20349 23891 20383
rect 26893 20349 26927 20383
rect 27353 20349 27387 20383
rect 27620 20349 27654 20383
rect 29745 20349 29779 20383
rect 29837 20349 29871 20383
rect 30573 20349 30607 20383
rect 30757 20349 30791 20383
rect 2973 20281 3007 20315
rect 6469 20281 6503 20315
rect 9045 20281 9079 20315
rect 10732 20281 10766 20315
rect 11437 20281 11471 20315
rect 14372 20281 14406 20315
rect 24685 20281 24719 20315
rect 26626 20281 26660 20315
rect 1777 20213 1811 20247
rect 2421 20213 2455 20247
rect 5825 20213 5859 20247
rect 7113 20213 7147 20247
rect 8217 20213 8251 20247
rect 9597 20213 9631 20247
rect 13185 20213 13219 20247
rect 15485 20213 15519 20247
rect 17141 20213 17175 20247
rect 21281 20213 21315 20247
rect 24961 20213 24995 20247
rect 2973 20009 3007 20043
rect 4261 20009 4295 20043
rect 8217 20009 8251 20043
rect 10793 20009 10827 20043
rect 13461 20009 13495 20043
rect 14105 20009 14139 20043
rect 21281 20009 21315 20043
rect 24593 20009 24627 20043
rect 31217 20009 31251 20043
rect 17908 19941 17942 19975
rect 19349 19941 19383 19975
rect 25728 19941 25762 19975
rect 1501 19873 1535 19907
rect 2329 19873 2363 19907
rect 2513 19873 2547 19907
rect 2605 19873 2639 19907
rect 2697 19873 2731 19907
rect 3433 19873 3467 19907
rect 3617 19873 3651 19907
rect 4169 19873 4203 19907
rect 5273 19873 5307 19907
rect 5362 19873 5396 19907
rect 5457 19873 5491 19907
rect 5641 19873 5675 19907
rect 6377 19873 6411 19907
rect 6561 19873 6595 19907
rect 7573 19873 7607 19907
rect 7757 19873 7791 19907
rect 7849 19873 7883 19907
rect 7941 19873 7975 19907
rect 8677 19873 8711 19907
rect 9413 19873 9447 19907
rect 10425 19873 10459 19907
rect 11989 19873 12023 19907
rect 12173 19873 12207 19907
rect 12725 19873 12759 19907
rect 13369 19873 13403 19907
rect 14749 19873 14783 19907
rect 15393 19873 15427 19907
rect 15577 19873 15611 19907
rect 15669 19873 15703 19907
rect 15945 19873 15979 19907
rect 18613 19873 18647 19907
rect 18797 19873 18831 19907
rect 18981 19873 19015 19907
rect 19165 19873 19199 19907
rect 19901 19873 19935 19907
rect 20168 19873 20202 19907
rect 22201 19873 22235 19907
rect 22468 19873 22502 19907
rect 27537 19873 27571 19907
rect 28457 19873 28491 19907
rect 29009 19873 29043 19907
rect 29837 19873 29871 19907
rect 30665 19873 30699 19907
rect 31309 19873 31343 19907
rect 3801 19805 3835 19839
rect 8953 19805 8987 19839
rect 12909 19805 12943 19839
rect 14841 19805 14875 19839
rect 15761 19805 15795 19839
rect 18153 19805 18187 19839
rect 18889 19805 18923 19839
rect 25973 19805 26007 19839
rect 27813 19805 27847 19839
rect 10977 19737 11011 19771
rect 16129 19737 16163 19771
rect 30481 19737 30515 19771
rect 1777 19669 1811 19703
rect 4997 19669 5031 19703
rect 6561 19669 6595 19703
rect 7021 19669 7055 19703
rect 8769 19669 8803 19703
rect 8861 19669 8895 19703
rect 9505 19669 9539 19703
rect 10793 19669 10827 19703
rect 16773 19669 16807 19703
rect 23581 19669 23615 19703
rect 24133 19669 24167 19703
rect 28365 19669 28399 19703
rect 29193 19669 29227 19703
rect 30021 19669 30055 19703
rect 6929 19465 6963 19499
rect 15853 19465 15887 19499
rect 20177 19465 20211 19499
rect 22385 19465 22419 19499
rect 6745 19397 6779 19431
rect 9689 19397 9723 19431
rect 13461 19397 13495 19431
rect 19349 19397 19383 19431
rect 3893 19329 3927 19363
rect 4077 19329 4111 19363
rect 6285 19329 6319 19363
rect 8033 19329 8067 19363
rect 8401 19329 8435 19363
rect 9505 19329 9539 19363
rect 9781 19329 9815 19363
rect 11253 19329 11287 19363
rect 11345 19329 11379 19363
rect 12449 19329 12483 19363
rect 12541 19329 12575 19363
rect 14933 19329 14967 19363
rect 16773 19329 16807 19363
rect 16865 19329 16899 19363
rect 17233 19329 17267 19363
rect 17693 19329 17727 19363
rect 17969 19329 18003 19363
rect 22017 19329 22051 19363
rect 24685 19329 24719 19363
rect 27353 19329 27387 19363
rect 27445 19329 27479 19363
rect 28549 19329 28583 19363
rect 28641 19329 28675 19363
rect 1869 19261 1903 19295
rect 2501 19261 2535 19295
rect 2676 19258 2710 19292
rect 2776 19261 2810 19295
rect 2881 19261 2915 19295
rect 5457 19261 5491 19295
rect 5641 19261 5675 19295
rect 6009 19261 6043 19295
rect 7665 19261 7699 19295
rect 7757 19261 7791 19295
rect 9229 19261 9263 19295
rect 9873 19261 9907 19295
rect 11069 19261 11103 19295
rect 11437 19261 11471 19295
rect 11621 19261 11655 19295
rect 12173 19261 12207 19295
rect 12357 19261 12391 19295
rect 12725 19261 12759 19295
rect 14749 19261 14783 19295
rect 15025 19261 15059 19295
rect 15113 19261 15147 19295
rect 15301 19261 15335 19295
rect 15945 19261 15979 19295
rect 16497 19261 16531 19295
rect 16681 19261 16715 19295
rect 17049 19261 17083 19295
rect 21290 19261 21324 19295
rect 21557 19261 21591 19295
rect 23121 19261 23155 19295
rect 23305 19261 23339 19295
rect 23765 19261 23799 19295
rect 24409 19261 24443 19295
rect 26249 19261 26283 19295
rect 27077 19261 27111 19295
rect 27261 19261 27295 19295
rect 27629 19261 27663 19295
rect 28273 19261 28307 19295
rect 28457 19261 28491 19295
rect 28825 19261 28859 19295
rect 29561 19261 29595 19295
rect 3157 19193 3191 19227
rect 6897 19193 6931 19227
rect 7113 19193 7147 19227
rect 8217 19193 8251 19227
rect 23213 19193 23247 19227
rect 1961 19125 1995 19159
rect 4169 19125 4203 19159
rect 4537 19125 4571 19159
rect 6285 19125 6319 19159
rect 10885 19125 10919 19159
rect 12909 19125 12943 19159
rect 14565 19125 14599 19159
rect 22385 19125 22419 19159
rect 22569 19125 22603 19159
rect 26157 19125 26191 19159
rect 27813 19125 27847 19159
rect 29009 19125 29043 19159
rect 30849 19125 30883 19159
rect 2789 18921 2823 18955
rect 3801 18921 3835 18955
rect 4445 18921 4479 18955
rect 6837 18921 6871 18955
rect 7665 18921 7699 18955
rect 8493 18921 8527 18955
rect 8953 18921 8987 18955
rect 13829 18921 13863 18955
rect 15669 18921 15703 18955
rect 19717 18921 19751 18955
rect 20913 18921 20947 18955
rect 21925 18921 21959 18955
rect 22569 18921 22603 18955
rect 30941 18921 30975 18955
rect 6745 18853 6779 18887
rect 9680 18853 9714 18887
rect 12716 18853 12750 18887
rect 28834 18853 28868 18887
rect 29806 18853 29840 18887
rect 1501 18785 1535 18819
rect 1685 18785 1719 18819
rect 2053 18785 2087 18819
rect 2697 18785 2731 18819
rect 2881 18785 2915 18819
rect 3893 18785 3927 18819
rect 4353 18785 4387 18819
rect 4537 18785 4571 18819
rect 5273 18785 5307 18819
rect 5365 18785 5399 18819
rect 5478 18785 5512 18819
rect 5641 18785 5675 18819
rect 7573 18785 7607 18819
rect 7757 18785 7791 18819
rect 8585 18785 8619 18819
rect 11621 18785 11655 18819
rect 14556 18785 14590 18819
rect 16681 18785 16715 18819
rect 16865 18785 16899 18819
rect 17049 18785 17083 18819
rect 17785 18785 17819 18819
rect 17885 18775 17919 18809
rect 18337 18785 18371 18819
rect 18604 18785 18638 18819
rect 20177 18785 20211 18819
rect 20361 18785 20395 18819
rect 20729 18785 20763 18819
rect 22017 18785 22051 18819
rect 22753 18785 22787 18819
rect 23397 18785 23431 18819
rect 23581 18785 23615 18819
rect 23673 18785 23707 18819
rect 23949 18785 23983 18819
rect 24869 18785 24903 18819
rect 25973 18785 26007 18819
rect 29101 18785 29135 18819
rect 29561 18785 29595 18819
rect 1777 18717 1811 18751
rect 1869 18717 1903 18751
rect 6929 18717 6963 18751
rect 8401 18717 8435 18751
rect 9413 18717 9447 18751
rect 12449 18717 12483 18751
rect 14289 18717 14323 18751
rect 20453 18717 20487 18751
rect 20545 18717 20579 18751
rect 23765 18717 23799 18751
rect 24593 18717 24627 18751
rect 2237 18581 2271 18615
rect 4997 18581 5031 18615
rect 6377 18581 6411 18615
rect 10793 18581 10827 18615
rect 16773 18581 16807 18615
rect 24133 18581 24167 18615
rect 27169 18581 27203 18615
rect 27721 18581 27755 18615
rect 8125 18377 8159 18411
rect 11805 18377 11839 18411
rect 14105 18377 14139 18411
rect 14841 18377 14875 18411
rect 15945 18377 15979 18411
rect 16957 18377 16991 18411
rect 17141 18377 17175 18411
rect 17693 18377 17727 18411
rect 8769 18309 8803 18343
rect 13369 18309 13403 18343
rect 15577 18309 15611 18343
rect 22017 18309 22051 18343
rect 4997 18241 5031 18275
rect 6929 18241 6963 18275
rect 2522 18173 2556 18207
rect 2789 18173 2823 18207
rect 5181 18173 5215 18207
rect 5273 18173 5307 18207
rect 6101 18173 6135 18207
rect 7021 18173 7055 18207
rect 7481 18173 7515 18207
rect 7665 18173 7699 18207
rect 7757 18173 7791 18207
rect 7849 18173 7883 18207
rect 9873 18241 9907 18275
rect 16589 18241 16623 18275
rect 18613 18241 18647 18275
rect 19625 18241 19659 18275
rect 24409 18241 24443 18275
rect 8953 18173 8987 18207
rect 9137 18173 9171 18207
rect 13553 18173 13587 18207
rect 18153 18173 18187 18207
rect 18337 18173 18371 18207
rect 19257 18173 19291 18207
rect 19441 18173 19475 18207
rect 19533 18173 19567 18207
rect 19809 18173 19843 18207
rect 20453 18173 20487 18207
rect 21189 18173 21223 18207
rect 23121 18173 23155 18207
rect 25329 18173 25363 18207
rect 27537 18173 27571 18207
rect 29929 18173 29963 18207
rect 8769 18105 8803 18139
rect 10517 18105 10551 18139
rect 14749 18105 14783 18139
rect 18705 18105 18739 18139
rect 21741 18105 21775 18139
rect 23765 18105 23799 18139
rect 27804 18105 27838 18139
rect 30196 18105 30230 18139
rect 1409 18037 1443 18071
rect 3985 18037 4019 18071
rect 4445 18037 4479 18071
rect 4997 18037 5031 18071
rect 6009 18037 6043 18071
rect 9045 18037 9079 18071
rect 12725 18037 12759 18071
rect 15945 18037 15979 18071
rect 16129 18037 16163 18071
rect 16957 18037 16991 18071
rect 19993 18037 20027 18071
rect 20545 18037 20579 18071
rect 22937 18037 22971 18071
rect 23673 18037 23707 18071
rect 26617 18037 26651 18071
rect 28917 18037 28951 18071
rect 31309 18037 31343 18071
rect 3985 17833 4019 17867
rect 8233 17833 8267 17867
rect 8401 17833 8435 17867
rect 13737 17833 13771 17867
rect 27721 17833 27755 17867
rect 31309 17833 31343 17867
rect 2145 17765 2179 17799
rect 2850 17765 2884 17799
rect 4629 17765 4663 17799
rect 8033 17765 8067 17799
rect 9229 17765 9263 17799
rect 9597 17765 9631 17799
rect 15945 17765 15979 17799
rect 17785 17765 17819 17799
rect 18245 17765 18279 17799
rect 19993 17765 20027 17799
rect 24317 17765 24351 17799
rect 25320 17765 25354 17799
rect 28609 17765 28643 17799
rect 28825 17765 28859 17799
rect 1409 17697 1443 17731
rect 1593 17697 1627 17731
rect 1685 17697 1719 17731
rect 1961 17697 1995 17731
rect 2605 17697 2639 17731
rect 5457 17697 5491 17731
rect 6929 17697 6963 17731
rect 10333 17697 10367 17731
rect 10701 17697 10735 17731
rect 10885 17697 10919 17731
rect 11529 17697 11563 17731
rect 12357 17697 12391 17731
rect 12624 17697 12658 17731
rect 14197 17697 14231 17731
rect 17049 17697 17083 17731
rect 17233 17697 17267 17731
rect 17325 17697 17359 17731
rect 17601 17697 17635 17731
rect 20453 17697 20487 17731
rect 20637 17697 20671 17731
rect 20729 17697 20763 17731
rect 21005 17697 21039 17731
rect 22293 17697 22327 17731
rect 22560 17697 22594 17731
rect 24225 17697 24259 17731
rect 26985 17697 27019 17731
rect 27169 17697 27203 17731
rect 27537 17697 27571 17731
rect 29285 17697 29319 17731
rect 30196 17697 30230 17731
rect 1777 17629 1811 17663
rect 5181 17629 5215 17663
rect 10517 17629 10551 17663
rect 10609 17629 10643 17663
rect 17417 17629 17451 17663
rect 20821 17629 20855 17663
rect 25053 17629 25087 17663
rect 27261 17629 27295 17663
rect 27353 17629 27387 17663
rect 29929 17629 29963 17663
rect 4445 17561 4479 17595
rect 6745 17561 6779 17595
rect 7573 17561 7607 17595
rect 5273 17493 5307 17527
rect 5365 17493 5399 17527
rect 8217 17493 8251 17527
rect 10149 17493 10183 17527
rect 11621 17493 11655 17527
rect 21189 17493 21223 17527
rect 23673 17493 23707 17527
rect 26433 17493 26467 17527
rect 28457 17493 28491 17527
rect 28641 17493 28675 17527
rect 29377 17493 29411 17527
rect 2145 17289 2179 17323
rect 7481 17289 7515 17323
rect 9413 17289 9447 17323
rect 13093 17289 13127 17323
rect 18521 17289 18555 17323
rect 30297 17289 30331 17323
rect 1593 17221 1627 17255
rect 14289 17221 14323 17255
rect 18705 17221 18739 17255
rect 24409 17221 24443 17255
rect 30849 17221 30883 17255
rect 5457 17153 5491 17187
rect 6101 17153 6135 17187
rect 6285 17153 6319 17187
rect 10241 17153 10275 17187
rect 10333 17153 10367 17187
rect 11437 17153 11471 17187
rect 11529 17153 11563 17187
rect 12633 17153 12667 17187
rect 18153 17153 18187 17187
rect 23397 17153 23431 17187
rect 27537 17153 27571 17187
rect 28181 17153 28215 17187
rect 31033 17153 31067 17187
rect 2789 17085 2823 17119
rect 4629 17085 4663 17119
rect 5733 17085 5767 17119
rect 6561 17085 6595 17119
rect 7389 17085 7423 17119
rect 9965 17085 9999 17119
rect 10149 17085 10183 17119
rect 10517 17085 10551 17119
rect 11161 17085 11195 17119
rect 11345 17085 11379 17119
rect 11713 17085 11747 17119
rect 12357 17085 12391 17119
rect 12541 17085 12575 17119
rect 12725 17085 12759 17119
rect 12909 17085 12943 17119
rect 14105 17085 14139 17119
rect 14289 17085 14323 17119
rect 15117 17085 15151 17119
rect 15301 17085 15335 17119
rect 15577 17085 15611 17119
rect 16221 17085 16255 17119
rect 17141 17085 17175 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 17509 17085 17543 17119
rect 17693 17085 17727 17119
rect 19441 17085 19475 17119
rect 19625 17085 19659 17119
rect 20177 17085 20211 17119
rect 20821 17085 20855 17119
rect 23121 17085 23155 17119
rect 23305 17085 23339 17119
rect 23489 17085 23523 17119
rect 23673 17085 23707 17119
rect 25789 17085 25823 17119
rect 26249 17085 26283 17119
rect 26525 17085 26559 17119
rect 28457 17085 28491 17119
rect 29561 17085 29595 17119
rect 29745 17087 29779 17121
rect 29837 17085 29871 17119
rect 29975 17085 30009 17119
rect 30113 17085 30147 17119
rect 30757 17085 30791 17119
rect 2237 17017 2271 17051
rect 8401 17017 8435 17051
rect 10701 17017 10735 17051
rect 14657 17017 14691 17051
rect 15669 17017 15703 17051
rect 18521 17017 18555 17051
rect 20361 17017 20395 17051
rect 21088 17017 21122 17051
rect 23857 17017 23891 17051
rect 25522 17017 25556 17051
rect 2973 16949 3007 16983
rect 4169 16949 4203 16983
rect 4721 16949 4755 16983
rect 11897 16949 11931 16983
rect 16405 16949 16439 16983
rect 16957 16949 16991 16983
rect 22201 16949 22235 16983
rect 30757 16949 30791 16983
rect 1409 16745 1443 16779
rect 3341 16745 3375 16779
rect 6469 16745 6503 16779
rect 10701 16745 10735 16779
rect 14013 16745 14047 16779
rect 14657 16745 14691 16779
rect 18061 16745 18095 16779
rect 21189 16745 21223 16779
rect 22661 16745 22695 16779
rect 23765 16745 23799 16779
rect 26985 16745 27019 16779
rect 30297 16745 30331 16779
rect 31125 16745 31159 16779
rect 5457 16677 5491 16711
rect 10517 16677 10551 16711
rect 27721 16677 27755 16711
rect 1961 16609 1995 16643
rect 2145 16609 2179 16643
rect 2237 16609 2271 16643
rect 2513 16609 2547 16643
rect 3157 16609 3191 16643
rect 4169 16609 4203 16643
rect 4721 16609 4755 16643
rect 4813 16609 4847 16643
rect 7582 16609 7616 16643
rect 8953 16609 8987 16643
rect 9413 16609 9447 16643
rect 11529 16609 11563 16643
rect 13277 16609 13311 16643
rect 13461 16609 13495 16643
rect 13829 16609 13863 16643
rect 14841 16609 14875 16643
rect 15393 16609 15427 16643
rect 15577 16609 15611 16643
rect 15945 16609 15979 16643
rect 16681 16609 16715 16643
rect 16948 16609 16982 16643
rect 18521 16609 18555 16643
rect 18705 16609 18739 16643
rect 18889 16609 18923 16643
rect 19073 16609 19107 16643
rect 19809 16609 19843 16643
rect 20065 16609 20099 16643
rect 22017 16609 22051 16643
rect 22201 16609 22235 16643
rect 22845 16609 22879 16643
rect 23121 16609 23155 16643
rect 23305 16609 23339 16643
rect 24593 16609 24627 16643
rect 25605 16609 25639 16643
rect 25881 16609 25915 16643
rect 28733 16609 28767 16643
rect 28917 16609 28951 16643
rect 29561 16609 29595 16643
rect 29745 16609 29779 16643
rect 30113 16609 30147 16643
rect 31309 16609 31343 16643
rect 2329 16541 2363 16575
rect 7849 16541 7883 16575
rect 11805 16541 11839 16575
rect 13553 16541 13587 16575
rect 13645 16541 13679 16575
rect 15669 16541 15703 16575
rect 15761 16541 15795 16575
rect 18797 16541 18831 16575
rect 21833 16541 21867 16575
rect 23029 16541 23063 16575
rect 24317 16541 24351 16575
rect 27905 16541 27939 16575
rect 28641 16541 28675 16575
rect 29101 16541 29135 16575
rect 29837 16541 29871 16575
rect 29929 16541 29963 16575
rect 3985 16473 4019 16507
rect 5641 16473 5675 16507
rect 9597 16473 9631 16507
rect 10149 16473 10183 16507
rect 19257 16473 19291 16507
rect 22937 16473 22971 16507
rect 2697 16405 2731 16439
rect 8861 16405 8895 16439
rect 10517 16405 10551 16439
rect 16129 16405 16163 16439
rect 3065 16201 3099 16235
rect 4353 16201 4387 16235
rect 6929 16201 6963 16235
rect 14473 16201 14507 16235
rect 20913 16201 20947 16235
rect 21833 16201 21867 16235
rect 24685 16201 24719 16235
rect 28457 16201 28491 16235
rect 29009 16201 29043 16235
rect 30113 16201 30147 16235
rect 2237 16065 2271 16099
rect 2513 16065 2547 16099
rect 4905 16065 4939 16099
rect 5089 16065 5123 16099
rect 5641 16065 5675 16099
rect 6561 16065 6595 16099
rect 7941 16065 7975 16099
rect 8309 16065 8343 16099
rect 10425 16065 10459 16099
rect 11253 16065 11287 16099
rect 15853 16065 15887 16099
rect 16313 16065 16347 16099
rect 17785 16065 17819 16099
rect 25237 16065 25271 16099
rect 4261 15997 4295 16031
rect 5181 15997 5215 16031
rect 6193 15997 6227 16031
rect 6377 15997 6411 16031
rect 6469 15997 6503 16031
rect 6745 15997 6779 16031
rect 7665 15997 7699 16031
rect 7757 15997 7791 16031
rect 8401 15997 8435 16031
rect 9045 15997 9079 16031
rect 9321 15997 9355 16031
rect 9689 15997 9723 16031
rect 10057 15997 10091 16031
rect 10977 15997 11011 16031
rect 11161 15997 11195 16031
rect 11345 15997 11379 16031
rect 11529 15997 11563 16031
rect 12173 15997 12207 16031
rect 16497 15997 16531 16031
rect 16773 15997 16807 16031
rect 17509 15997 17543 16031
rect 17693 15997 17727 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 19625 15997 19659 16031
rect 22017 15997 22051 16031
rect 23857 15997 23891 16031
rect 24593 15997 24627 16031
rect 27077 15997 27111 16031
rect 30665 15997 30699 16031
rect 3157 15929 3191 15963
rect 11713 15929 11747 15963
rect 12418 15929 12452 15963
rect 15586 15929 15620 15963
rect 16865 15929 16899 15963
rect 23612 15929 23646 15963
rect 25504 15929 25538 15963
rect 27344 15929 27378 15963
rect 30021 15929 30055 15963
rect 4905 15861 4939 15895
rect 13553 15861 13587 15895
rect 18245 15861 18279 15895
rect 22477 15861 22511 15895
rect 26617 15861 26651 15895
rect 30757 15861 30791 15895
rect 1593 15657 1627 15691
rect 4813 15657 4847 15691
rect 7021 15657 7055 15691
rect 8861 15657 8895 15691
rect 10701 15657 10735 15691
rect 15393 15657 15427 15691
rect 15945 15657 15979 15691
rect 22109 15657 22143 15691
rect 23581 15657 23615 15691
rect 25789 15657 25823 15691
rect 27721 15657 27755 15691
rect 31049 15657 31083 15691
rect 6193 15589 6227 15623
rect 6653 15589 6687 15623
rect 6869 15589 6903 15623
rect 9588 15589 9622 15623
rect 11796 15589 11830 15623
rect 13737 15589 13771 15623
rect 22277 15589 22311 15623
rect 22477 15589 22511 15623
rect 26341 15589 26375 15623
rect 28181 15589 28215 15623
rect 30849 15589 30883 15623
rect 1409 15521 1443 15555
rect 2237 15521 2271 15555
rect 2504 15521 2538 15555
rect 4445 15521 4479 15555
rect 5273 15521 5307 15555
rect 4261 15453 4295 15487
rect 4353 15453 4387 15487
rect 5549 15453 5583 15487
rect 3617 15385 3651 15419
rect 7757 15521 7791 15555
rect 7849 15521 7883 15555
rect 7941 15521 7975 15555
rect 8125 15521 8159 15555
rect 8585 15521 8619 15555
rect 11529 15521 11563 15555
rect 13369 15521 13403 15555
rect 14657 15521 14691 15555
rect 14841 15521 14875 15555
rect 14933 15521 14967 15555
rect 15209 15521 15243 15555
rect 15853 15521 15887 15555
rect 16773 15521 16807 15555
rect 17509 15521 17543 15555
rect 18153 15521 18187 15555
rect 18705 15521 18739 15555
rect 18889 15521 18923 15555
rect 18981 15521 19015 15555
rect 19257 15521 19291 15555
rect 19441 15521 19475 15555
rect 20269 15521 20303 15555
rect 20637 15521 20671 15555
rect 21189 15521 21223 15555
rect 23121 15521 23155 15555
rect 23213 15521 23247 15555
rect 23397 15521 23431 15555
rect 24501 15521 24535 15555
rect 26985 15521 27019 15555
rect 27169 15521 27203 15555
rect 27353 15521 27387 15555
rect 27537 15521 27571 15555
rect 28365 15521 28399 15555
rect 29285 15521 29319 15555
rect 8861 15453 8895 15487
rect 9321 15453 9355 15487
rect 15025 15453 15059 15487
rect 17417 15453 17451 15487
rect 19073 15453 19107 15487
rect 24777 15453 24811 15487
rect 27261 15453 27295 15487
rect 29561 15453 29595 15487
rect 13921 15385 13955 15419
rect 17969 15385 18003 15419
rect 20269 15385 20303 15419
rect 5365 15317 5399 15351
rect 5457 15317 5491 15351
rect 6193 15317 6227 15351
rect 6837 15317 6871 15351
rect 7481 15317 7515 15351
rect 8677 15317 8711 15351
rect 12909 15317 12943 15351
rect 13737 15317 13771 15351
rect 22293 15317 22327 15351
rect 31033 15317 31067 15351
rect 31217 15317 31251 15351
rect 1593 15113 1627 15147
rect 4077 15113 4111 15147
rect 8401 15113 8435 15147
rect 9689 15113 9723 15147
rect 12035 15113 12069 15147
rect 13461 15113 13495 15147
rect 15669 15113 15703 15147
rect 18061 15113 18095 15147
rect 18521 15113 18555 15147
rect 18705 15113 18739 15147
rect 20269 15113 20303 15147
rect 20453 15113 20487 15147
rect 23121 15113 23155 15147
rect 23857 15113 23891 15147
rect 24501 15113 24535 15147
rect 25053 15113 25087 15147
rect 25789 15113 25823 15147
rect 27629 15113 27663 15147
rect 28365 15113 28399 15147
rect 29653 15113 29687 15147
rect 7113 15045 7147 15079
rect 7205 15045 7239 15079
rect 13277 15045 13311 15079
rect 16497 15045 16531 15079
rect 2881 14977 2915 15011
rect 5549 14977 5583 15011
rect 6193 14977 6227 15011
rect 7297 14977 7331 15011
rect 8953 14977 8987 15011
rect 2605 14909 2639 14943
rect 4813 14909 4847 14943
rect 5089 14909 5123 14943
rect 5825 14909 5859 14943
rect 7021 14909 7055 14943
rect 7757 14909 7791 14943
rect 7941 14909 7975 14943
rect 8033 14909 8067 14943
rect 8125 14909 8159 14943
rect 9505 14909 9539 14943
rect 10241 14909 10275 14943
rect 10517 14909 10551 14943
rect 11805 14909 11839 14943
rect 3893 14841 3927 14875
rect 13553 14909 13587 14943
rect 16313 14909 16347 14943
rect 17141 14909 17175 14943
rect 14197 14841 14231 14875
rect 17417 14841 17451 14875
rect 19901 15045 19935 15079
rect 28825 15045 28859 15079
rect 21189 14977 21223 15011
rect 18153 14909 18187 14943
rect 19257 14909 19291 14943
rect 19441 14909 19475 14943
rect 23213 14909 23247 14943
rect 23673 14909 23707 14943
rect 23857 14909 23891 14943
rect 24409 14909 24443 14943
rect 24593 14909 24627 14943
rect 25973 14909 26007 14943
rect 26157 14909 26191 14943
rect 26249 14909 26283 14943
rect 26341 14909 26375 14943
rect 26525 14909 26559 14943
rect 28181 14909 28215 14943
rect 29009 14909 29043 14943
rect 31033 14909 31067 14943
rect 20269 14841 20303 14875
rect 21456 14841 21490 14875
rect 30766 14841 30800 14875
rect 4093 14773 4127 14807
rect 4261 14773 4295 14807
rect 13277 14773 13311 14807
rect 14657 14773 14691 14807
rect 18061 14773 18095 14807
rect 18521 14773 18555 14807
rect 19349 14773 19383 14807
rect 22569 14773 22603 14807
rect 27077 14773 27111 14807
rect 3801 14569 3835 14603
rect 7665 14569 7699 14603
rect 8493 14569 8527 14603
rect 8953 14569 8987 14603
rect 10149 14569 10183 14603
rect 10609 14569 10643 14603
rect 12173 14569 12207 14603
rect 15669 14569 15703 14603
rect 19165 14569 19199 14603
rect 21189 14569 21223 14603
rect 24041 14569 24075 14603
rect 27629 14569 27663 14603
rect 30389 14569 30423 14603
rect 31309 14569 31343 14603
rect 4445 14501 4479 14535
rect 17049 14501 17083 14535
rect 18052 14501 18086 14535
rect 2329 14433 2363 14467
rect 3065 14433 3099 14467
rect 3157 14433 3191 14467
rect 3341 14433 3375 14467
rect 3433 14433 3467 14467
rect 3525 14433 3559 14467
rect 4261 14433 4295 14467
rect 4537 14433 4571 14467
rect 4997 14433 5031 14467
rect 5641 14433 5675 14467
rect 5825 14433 5859 14467
rect 6561 14433 6595 14467
rect 6745 14433 6779 14467
rect 6929 14433 6963 14467
rect 7113 14433 7147 14467
rect 7573 14433 7607 14467
rect 7757 14433 7791 14467
rect 8585 14433 8619 14467
rect 9413 14433 9447 14467
rect 9597 14433 9631 14467
rect 13093 14433 13127 14467
rect 13360 14433 13394 14467
rect 14933 14433 14967 14467
rect 15117 14433 15151 14467
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 19809 14433 19843 14467
rect 20065 14433 20099 14467
rect 21993 14433 22027 14467
rect 22661 14433 22695 14467
rect 22928 14433 22962 14467
rect 24501 14433 24535 14467
rect 24685 14433 24719 14467
rect 25053 14433 25087 14467
rect 25697 14433 25731 14467
rect 25881 14433 25915 14467
rect 25973 14433 26007 14467
rect 26249 14433 26283 14467
rect 26985 14433 27019 14467
rect 28457 14433 28491 14467
rect 28641 14433 28675 14467
rect 28733 14433 28767 14467
rect 29009 14433 29043 14467
rect 29653 14433 29687 14467
rect 29837 14433 29871 14467
rect 30205 14433 30239 14467
rect 31125 14433 31159 14467
rect 2605 14365 2639 14399
rect 4813 14365 4847 14399
rect 6837 14365 6871 14399
rect 8401 14365 8435 14399
rect 9505 14365 9539 14399
rect 15209 14365 15243 14399
rect 16681 14365 16715 14399
rect 17785 14365 17819 14399
rect 24777 14365 24811 14399
rect 24869 14365 24903 14399
rect 26065 14365 26099 14399
rect 28825 14365 28859 14399
rect 29929 14365 29963 14399
rect 30021 14365 30055 14399
rect 30849 14365 30883 14399
rect 30941 14365 30975 14399
rect 3065 14297 3099 14331
rect 14473 14297 14507 14331
rect 6377 14229 6411 14263
rect 11621 14229 11655 14263
rect 17049 14229 17083 14263
rect 17233 14229 17267 14263
rect 21925 14229 21959 14263
rect 25237 14229 25271 14263
rect 26433 14229 26467 14263
rect 27077 14229 27111 14263
rect 29193 14229 29227 14263
rect 1501 14025 1535 14059
rect 3157 14025 3191 14059
rect 4445 14025 4479 14059
rect 7205 14025 7239 14059
rect 9045 14025 9079 14059
rect 11437 14025 11471 14059
rect 13553 14025 13587 14059
rect 20913 14025 20947 14059
rect 21373 14025 21407 14059
rect 23397 14025 23431 14059
rect 27169 14025 27203 14059
rect 29561 14025 29595 14059
rect 30757 14025 30791 14059
rect 7757 13957 7791 13991
rect 21649 13957 21683 13991
rect 30849 13957 30883 13991
rect 2329 13889 2363 13923
rect 8309 13889 8343 13923
rect 11989 13889 12023 13923
rect 13185 13889 13219 13923
rect 15393 13889 15427 13923
rect 16865 13889 16899 13923
rect 16957 13889 16991 13923
rect 18245 13889 18279 13923
rect 19533 13889 19567 13923
rect 21741 13889 21775 13923
rect 24685 13889 24719 13923
rect 31033 13889 31067 13923
rect 2145 13821 2179 13855
rect 2421 13821 2455 13855
rect 2513 13821 2547 13855
rect 2697 13821 2731 13855
rect 3801 13821 3835 13855
rect 3985 13821 4019 13855
rect 4077 13821 4111 13855
rect 4189 13821 4223 13855
rect 5825 13821 5859 13855
rect 6092 13821 6126 13855
rect 7665 13821 7699 13855
rect 8953 13821 8987 13855
rect 9597 13821 9631 13855
rect 12817 13821 12851 13855
rect 13001 13821 13035 13855
rect 13093 13821 13127 13855
rect 13369 13821 13403 13855
rect 15669 13821 15703 13855
rect 16589 13823 16623 13857
rect 16761 13815 16795 13849
rect 17141 13821 17175 13855
rect 17325 13821 17359 13855
rect 17785 13821 17819 13855
rect 17969 13821 18003 13855
rect 21557 13821 21591 13855
rect 21833 13821 21867 13855
rect 22017 13821 22051 13855
rect 22477 13821 22511 13855
rect 22661 13821 22695 13855
rect 22845 13821 22879 13855
rect 22937 13821 22971 13855
rect 23581 13821 23615 13855
rect 24409 13821 24443 13855
rect 24593 13821 24627 13855
rect 24777 13821 24811 13855
rect 24961 13821 24995 13855
rect 25789 13821 25823 13855
rect 26056 13821 26090 13855
rect 28089 13821 28123 13855
rect 28273 13821 28307 13855
rect 28365 13821 28399 13855
rect 28457 13821 28491 13855
rect 28641 13821 28675 13855
rect 30113 13821 30147 13855
rect 30757 13821 30791 13855
rect 5273 13753 5307 13787
rect 9864 13753 9898 13787
rect 14197 13753 14231 13787
rect 18337 13753 18371 13787
rect 19800 13753 19834 13787
rect 1961 13685 1995 13719
rect 5181 13685 5215 13719
rect 10977 13685 11011 13719
rect 25145 13685 25179 13719
rect 27905 13685 27939 13719
rect 30297 13685 30331 13719
rect 1409 13481 1443 13515
rect 5181 13481 5215 13515
rect 5825 13481 5859 13515
rect 7849 13481 7883 13515
rect 9781 13481 9815 13515
rect 13553 13481 13587 13515
rect 14749 13481 14783 13515
rect 17877 13481 17911 13515
rect 20269 13481 20303 13515
rect 22401 13481 22435 13515
rect 22569 13481 22603 13515
rect 23581 13481 23615 13515
rect 24041 13481 24075 13515
rect 2544 13413 2578 13447
rect 3249 13413 3283 13447
rect 8769 13413 8803 13447
rect 9321 13413 9355 13447
rect 13461 13413 13495 13447
rect 15862 13413 15896 13447
rect 18990 13413 19024 13447
rect 22201 13413 22235 13447
rect 29478 13413 29512 13447
rect 2789 13345 2823 13379
rect 3433 13345 3467 13379
rect 3801 13345 3835 13379
rect 3997 13355 4031 13389
rect 4629 13345 4663 13379
rect 5089 13345 5123 13379
rect 6561 13345 6595 13379
rect 6745 13345 6779 13379
rect 7113 13345 7147 13379
rect 7941 13345 7975 13379
rect 9965 13345 9999 13379
rect 10333 13345 10367 13379
rect 10517 13345 10551 13379
rect 11785 13345 11819 13379
rect 14289 13345 14323 13379
rect 16129 13345 16163 13379
rect 16865 13345 16899 13379
rect 17049 13345 17083 13379
rect 17138 13345 17172 13379
rect 17245 13347 17279 13381
rect 17417 13345 17451 13379
rect 19257 13345 19291 13379
rect 25154 13345 25188 13379
rect 25421 13345 25455 13379
rect 25881 13345 25915 13379
rect 27169 13345 27203 13379
rect 27261 13345 27295 13379
rect 29745 13345 29779 13379
rect 30573 13345 30607 13379
rect 3617 13277 3651 13311
rect 3709 13277 3743 13311
rect 6837 13277 6871 13311
rect 6929 13277 6963 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 11529 13277 11563 13311
rect 26985 13277 27019 13311
rect 30849 13277 30883 13311
rect 12909 13209 12943 13243
rect 19717 13209 19751 13243
rect 27721 13209 27755 13243
rect 30665 13209 30699 13243
rect 4537 13141 4571 13175
rect 7297 13141 7331 13175
rect 14197 13141 14231 13175
rect 16681 13141 16715 13175
rect 21281 13141 21315 13175
rect 22385 13141 22419 13175
rect 25973 13141 26007 13175
rect 27077 13141 27111 13175
rect 28365 13141 28399 13175
rect 30757 13141 30791 13175
rect 5089 12937 5123 12971
rect 6101 12937 6135 12971
rect 10333 12937 10367 12971
rect 11529 12937 11563 12971
rect 15669 12937 15703 12971
rect 19993 12937 20027 12971
rect 21925 12937 21959 12971
rect 22109 12937 22143 12971
rect 23673 12937 23707 12971
rect 29009 12937 29043 12971
rect 31033 12937 31067 12971
rect 3249 12869 3283 12903
rect 13277 12869 13311 12903
rect 5917 12801 5951 12835
rect 7021 12801 7055 12835
rect 11161 12801 11195 12835
rect 14657 12801 14691 12835
rect 14749 12801 14783 12835
rect 17049 12801 17083 12835
rect 17601 12801 17635 12835
rect 19533 12801 19567 12835
rect 20729 12801 20763 12835
rect 25053 12801 25087 12835
rect 30021 12801 30055 12835
rect 1869 12733 1903 12767
rect 4445 12733 4479 12767
rect 4905 12733 4939 12767
rect 5089 12733 5123 12767
rect 6193 12733 6227 12767
rect 6653 12733 6687 12767
rect 6837 12733 6871 12767
rect 6929 12733 6963 12767
rect 7205 12733 7239 12767
rect 7849 12733 7883 12767
rect 8953 12733 8987 12767
rect 10793 12733 10827 12767
rect 10977 12733 11011 12767
rect 11069 12733 11103 12767
rect 11345 12733 11379 12767
rect 12357 12733 12391 12767
rect 12633 12733 12667 12767
rect 14473 12733 14507 12767
rect 14841 12733 14875 12767
rect 15025 12733 15059 12767
rect 16782 12733 16816 12767
rect 17509 12733 17543 12767
rect 19257 12733 19291 12767
rect 19441 12733 19475 12767
rect 19625 12733 19659 12767
rect 19809 12733 19843 12767
rect 22569 12733 22603 12767
rect 23029 12733 23063 12767
rect 24501 12733 24535 12767
rect 25789 12733 25823 12767
rect 26893 12733 26927 12767
rect 27077 12733 27111 12767
rect 27169 12733 27203 12767
rect 27629 12733 27663 12767
rect 29653 12733 29687 12767
rect 29837 12733 29871 12767
rect 29929 12733 29963 12767
rect 30205 12733 30239 12767
rect 2114 12665 2148 12699
rect 4353 12665 4387 12699
rect 9220 12665 9254 12699
rect 12725 12665 12759 12699
rect 13093 12665 13127 12699
rect 21741 12665 21775 12699
rect 27896 12665 27930 12699
rect 31217 12665 31251 12699
rect 5917 12597 5951 12631
rect 7389 12597 7423 12631
rect 7941 12597 7975 12631
rect 14289 12597 14323 12631
rect 18245 12597 18279 12631
rect 21189 12597 21223 12631
rect 21941 12597 21975 12631
rect 25973 12597 26007 12631
rect 26709 12597 26743 12631
rect 30389 12597 30423 12631
rect 30849 12597 30883 12631
rect 31007 12597 31041 12631
rect 1593 12393 1627 12427
rect 2605 12393 2639 12427
rect 3249 12393 3283 12427
rect 3801 12393 3835 12427
rect 9045 12393 9079 12427
rect 12265 12393 12299 12427
rect 13277 12393 13311 12427
rect 15485 12393 15519 12427
rect 15945 12393 15979 12427
rect 23489 12393 23523 12427
rect 24685 12393 24719 12427
rect 27353 12393 27387 12427
rect 29377 12393 29411 12427
rect 31309 12393 31343 12427
rect 11897 12325 11931 12359
rect 12113 12325 12147 12359
rect 13093 12325 13127 12359
rect 14372 12325 14406 12359
rect 25798 12325 25832 12359
rect 26985 12325 27019 12359
rect 27201 12325 27235 12359
rect 30196 12325 30230 12359
rect 1409 12257 1443 12291
rect 3709 12257 3743 12291
rect 3893 12257 3927 12291
rect 4721 12257 4755 12291
rect 5365 12257 5399 12291
rect 5733 12257 5767 12291
rect 7021 12257 7055 12291
rect 8217 12257 8251 12291
rect 8401 12257 8435 12291
rect 10241 12257 10275 12291
rect 10425 12257 10459 12291
rect 10793 12257 10827 12291
rect 12725 12257 12759 12291
rect 17693 12257 17727 12291
rect 17877 12257 17911 12291
rect 18061 12257 18095 12291
rect 18245 12257 18279 12291
rect 19809 12257 19843 12291
rect 22201 12257 22235 12291
rect 22753 12257 22787 12291
rect 23673 12257 23707 12291
rect 26065 12257 26099 12291
rect 27905 12257 27939 12291
rect 28549 12257 28583 12291
rect 29285 12257 29319 12291
rect 4905 12189 4939 12223
rect 7297 12189 7331 12223
rect 10517 12189 10551 12223
rect 10609 12189 10643 12223
rect 14105 12189 14139 12223
rect 17969 12189 18003 12223
rect 19625 12189 19659 12223
rect 21281 12189 21315 12223
rect 21925 12189 21959 12223
rect 22937 12189 22971 12223
rect 23949 12189 23983 12223
rect 29929 12189 29963 12223
rect 5089 12121 5123 12155
rect 9597 12053 9631 12087
rect 10977 12053 11011 12087
rect 12081 12053 12115 12087
rect 13093 12053 13127 12087
rect 16681 12053 16715 12087
rect 17509 12053 17543 12087
rect 18705 12053 18739 12087
rect 19993 12053 20027 12087
rect 20453 12053 20487 12087
rect 23857 12053 23891 12087
rect 27169 12053 27203 12087
rect 28457 12053 28491 12087
rect 2973 11849 3007 11883
rect 9597 11849 9631 11883
rect 13369 11849 13403 11883
rect 14381 11849 14415 11883
rect 20821 11849 20855 11883
rect 21005 11849 21039 11883
rect 21925 11849 21959 11883
rect 22109 11849 22143 11883
rect 24409 11849 24443 11883
rect 24593 11849 24627 11883
rect 30941 11849 30975 11883
rect 5457 11781 5491 11815
rect 26065 11781 26099 11815
rect 1869 11713 1903 11747
rect 1961 11713 1995 11747
rect 7021 11713 7055 11747
rect 11161 11713 11195 11747
rect 15577 11713 15611 11747
rect 19625 11713 19659 11747
rect 21557 11713 21591 11747
rect 23305 11713 23339 11747
rect 28549 11713 28583 11747
rect 28641 11713 28675 11747
rect 29837 11713 29871 11747
rect 29929 11713 29963 11747
rect 30849 11713 30883 11747
rect 1593 11645 1627 11679
rect 1777 11645 1811 11679
rect 2145 11645 2179 11679
rect 2789 11645 2823 11679
rect 4169 11645 4203 11679
rect 6377 11645 6411 11679
rect 6561 11645 6595 11679
rect 7288 11645 7322 11679
rect 9781 11645 9815 11679
rect 9965 11645 9999 11679
rect 10057 11645 10091 11679
rect 10149 11645 10183 11679
rect 10333 11645 10367 11679
rect 11345 11645 11379 11679
rect 11989 11645 12023 11679
rect 16773 11645 16807 11679
rect 17049 11645 17083 11679
rect 19257 11645 19291 11679
rect 19441 11645 19475 11679
rect 19533 11645 19567 11679
rect 19809 11645 19843 11679
rect 20453 11645 20487 11679
rect 23029 11645 23063 11679
rect 24961 11645 24995 11679
rect 25697 11645 25731 11679
rect 25881 11645 25915 11679
rect 25973 11645 26007 11679
rect 26157 11645 26191 11679
rect 26985 11645 27019 11679
rect 27169 11645 27203 11679
rect 27629 11645 27663 11679
rect 27813 11645 27847 11679
rect 28273 11645 28307 11679
rect 28457 11645 28491 11679
rect 28825 11645 28859 11679
rect 29561 11645 29595 11679
rect 29745 11645 29779 11679
rect 30113 11645 30147 11679
rect 31125 11645 31159 11679
rect 12256 11577 12290 11611
rect 14933 11577 14967 11611
rect 15761 11577 15795 11611
rect 18613 11577 18647 11611
rect 2329 11509 2363 11543
rect 6469 11509 6503 11543
rect 8401 11509 8435 11543
rect 9045 11509 9079 11543
rect 11529 11509 11563 11543
rect 15025 11509 15059 11543
rect 18061 11509 18095 11543
rect 19993 11509 20027 11543
rect 20830 11509 20864 11543
rect 21925 11509 21959 11543
rect 24593 11509 24627 11543
rect 26341 11509 26375 11543
rect 27077 11509 27111 11543
rect 27629 11509 27663 11543
rect 29009 11509 29043 11543
rect 30297 11509 30331 11543
rect 31309 11509 31343 11543
rect 5457 11305 5491 11339
rect 8769 11305 8803 11339
rect 9413 11305 9447 11339
rect 12173 11305 12207 11339
rect 12633 11305 12667 11339
rect 15577 11305 15611 11339
rect 16865 11305 16899 11339
rect 20729 11305 20763 11339
rect 22293 11305 22327 11339
rect 24317 11305 24351 11339
rect 25881 11305 25915 11339
rect 27169 11305 27203 11339
rect 30573 11305 30607 11339
rect 31309 11305 31343 11339
rect 6529 11237 6563 11271
rect 6745 11237 6779 11271
rect 7634 11237 7668 11271
rect 13461 11237 13495 11271
rect 14013 11237 14047 11271
rect 16957 11237 16991 11271
rect 19616 11237 19650 11271
rect 25007 11237 25041 11271
rect 28273 11237 28307 11271
rect 1961 11169 1995 11203
rect 2145 11169 2179 11203
rect 2329 11169 2363 11203
rect 2513 11169 2547 11203
rect 3157 11169 3191 11203
rect 3525 11169 3559 11203
rect 3709 11169 3743 11203
rect 4905 11169 4939 11203
rect 5457 11169 5491 11203
rect 7389 11169 7423 11203
rect 9229 11169 9263 11203
rect 10149 11169 10183 11203
rect 11989 11169 12023 11203
rect 14749 11169 14783 11203
rect 15485 11169 15519 11203
rect 17509 11169 17543 11203
rect 17765 11169 17799 11203
rect 22109 11169 22143 11203
rect 23204 11169 23238 11203
rect 24777 11169 24811 11203
rect 25421 11169 25455 11203
rect 25881 11169 25915 11203
rect 26065 11169 26099 11203
rect 27353 11169 27387 11203
rect 27445 11169 27479 11203
rect 27629 11169 27663 11203
rect 27813 11169 27847 11203
rect 31125 11169 31159 11203
rect 2237 11101 2271 11135
rect 3341 11101 3375 11135
rect 3433 11101 3467 11135
rect 4721 11101 4755 11135
rect 5089 11101 5123 11135
rect 10425 11101 10459 11135
rect 14197 11101 14231 11135
rect 19349 11101 19383 11135
rect 22937 11101 22971 11135
rect 27537 11101 27571 11135
rect 1777 11033 1811 11067
rect 6377 11033 6411 11067
rect 2973 10965 3007 10999
rect 6561 10965 6595 10999
rect 14841 10965 14875 10999
rect 18889 10965 18923 10999
rect 25053 10965 25087 10999
rect 29561 10965 29595 10999
rect 3985 10761 4019 10795
rect 5641 10761 5675 10795
rect 10609 10761 10643 10795
rect 19441 10761 19475 10795
rect 19625 10761 19659 10795
rect 21465 10761 21499 10795
rect 24501 10761 24535 10795
rect 28549 10761 28583 10795
rect 30941 10761 30975 10795
rect 2973 10625 3007 10659
rect 3249 10625 3283 10659
rect 4077 10625 4111 10659
rect 4537 10625 4571 10659
rect 5641 10625 5675 10659
rect 6009 10625 6043 10659
rect 6101 10625 6135 10659
rect 8033 10625 8067 10659
rect 18337 10625 18371 10659
rect 20085 10625 20119 10659
rect 27261 10625 27295 10659
rect 1961 10557 1995 10591
rect 3801 10557 3835 10591
rect 3893 10557 3927 10591
rect 4793 10557 4827 10591
rect 4905 10557 4939 10591
rect 5018 10557 5052 10591
rect 5181 10557 5215 10591
rect 5733 10557 5767 10591
rect 5917 10557 5951 10591
rect 6285 10557 6319 10591
rect 7113 10557 7147 10591
rect 7849 10557 7883 10591
rect 8125 10557 8159 10591
rect 8217 10557 8251 10591
rect 8401 10557 8435 10591
rect 9505 10557 9539 10591
rect 9781 10557 9815 10591
rect 11722 10557 11756 10591
rect 11989 10557 12023 10591
rect 12449 10557 12483 10591
rect 12633 10557 12667 10591
rect 13553 10557 13587 10591
rect 14105 10557 14139 10591
rect 16129 10557 16163 10591
rect 17969 10557 18003 10591
rect 18153 10557 18187 10591
rect 18245 10557 18279 10591
rect 18521 10557 18555 10591
rect 22293 10557 22327 10591
rect 22477 10557 22511 10591
rect 22569 10557 22603 10591
rect 23121 10557 23155 10591
rect 23305 10557 23339 10591
rect 25145 10557 25179 10591
rect 26617 10557 26651 10591
rect 26801 10557 26835 10591
rect 27537 10557 27571 10591
rect 29561 10557 29595 10591
rect 29817 10557 29851 10591
rect 1869 10489 1903 10523
rect 14372 10489 14406 10523
rect 16396 10489 16430 10523
rect 19257 10489 19291 10523
rect 19473 10489 19507 10523
rect 20352 10489 20386 10523
rect 24961 10489 24995 10523
rect 25789 10489 25823 10523
rect 25973 10489 26007 10523
rect 6469 10421 6503 10455
rect 7021 10421 7055 10455
rect 7665 10421 7699 10455
rect 12541 10421 12575 10455
rect 13461 10421 13495 10455
rect 15485 10421 15519 10455
rect 17509 10421 17543 10455
rect 18705 10421 18739 10455
rect 22109 10421 22143 10455
rect 23489 10421 23523 10455
rect 25329 10421 25363 10455
rect 26157 10421 26191 10455
rect 26709 10421 26743 10455
rect 2421 10217 2455 10251
rect 5457 10217 5491 10251
rect 7757 10217 7791 10251
rect 8493 10217 8527 10251
rect 10333 10217 10367 10251
rect 13001 10217 13035 10251
rect 14289 10217 14323 10251
rect 19441 10217 19475 10251
rect 20269 10217 20303 10251
rect 23213 10217 23247 10251
rect 30941 10217 30975 10251
rect 3534 10149 3568 10183
rect 6622 10149 6656 10183
rect 9198 10149 9232 10183
rect 12357 10149 12391 10183
rect 24869 10149 24903 10183
rect 29828 10149 29862 10183
rect 4537 10081 4571 10115
rect 5365 10081 5399 10115
rect 6377 10081 6411 10115
rect 10793 10081 10827 10115
rect 11805 10081 11839 10115
rect 13553 10081 13587 10115
rect 13737 10081 13771 10115
rect 13829 10081 13863 10115
rect 14105 10081 14139 10115
rect 15005 10081 15039 10115
rect 18061 10081 18095 10115
rect 18328 10081 18362 10115
rect 20085 10081 20119 10115
rect 20729 10081 20763 10115
rect 22017 10081 22051 10115
rect 22293 10081 22327 10115
rect 22477 10081 22511 10115
rect 23397 10081 23431 10115
rect 24041 10081 24075 10115
rect 24133 10081 24167 10115
rect 24685 10081 24719 10115
rect 25513 10081 25547 10115
rect 25881 10081 25915 10115
rect 28098 10081 28132 10115
rect 3801 10013 3835 10047
rect 5273 10013 5307 10047
rect 8953 10013 8987 10047
rect 12541 10013 12575 10047
rect 13921 10013 13955 10047
rect 14749 10013 14783 10047
rect 17233 10013 17267 10047
rect 17509 10013 17543 10047
rect 22201 10013 22235 10047
rect 28365 10013 28399 10047
rect 29561 10013 29595 10047
rect 22109 9945 22143 9979
rect 26985 9945 27019 9979
rect 1961 9877 1995 9911
rect 4445 9877 4479 9911
rect 5825 9877 5859 9911
rect 10885 9877 10919 9911
rect 11713 9877 11747 9911
rect 16129 9877 16163 9911
rect 20821 9877 20855 9911
rect 21833 9877 21867 9911
rect 25053 9877 25087 9911
rect 25605 9877 25639 9911
rect 26065 9877 26099 9911
rect 28825 9877 28859 9911
rect 14841 9673 14875 9707
rect 22753 9673 22787 9707
rect 23581 9673 23615 9707
rect 4905 9605 4939 9639
rect 5457 9605 5491 9639
rect 7389 9605 7423 9639
rect 10425 9605 10459 9639
rect 12449 9605 12483 9639
rect 16773 9605 16807 9639
rect 17969 9605 18003 9639
rect 20177 9605 20211 9639
rect 22201 9605 22235 9639
rect 30113 9605 30147 9639
rect 13001 9537 13035 9571
rect 15301 9537 15335 9571
rect 24777 9537 24811 9571
rect 26709 9537 26743 9571
rect 2522 9469 2556 9503
rect 2789 9469 2823 9503
rect 4261 9469 4295 9503
rect 4445 9469 4479 9503
rect 4540 9469 4574 9503
rect 4629 9469 4663 9503
rect 6101 9469 6135 9503
rect 8309 9469 8343 9503
rect 9045 9469 9079 9503
rect 9321 9469 9355 9503
rect 11621 9469 11655 9503
rect 14105 9469 14139 9503
rect 15025 9469 15059 9503
rect 15209 9469 15243 9503
rect 15393 9469 15427 9503
rect 15577 9469 15611 9503
rect 16037 9469 16071 9503
rect 16221 9469 16255 9503
rect 16313 9469 16347 9503
rect 16405 9469 16439 9503
rect 16589 9469 16623 9503
rect 19633 9469 19667 9503
rect 20085 9469 20119 9503
rect 20821 9469 20855 9503
rect 21088 9469 21122 9503
rect 22845 9469 22879 9503
rect 24685 9469 24719 9503
rect 25329 9469 25363 9503
rect 25513 9469 25547 9503
rect 26433 9469 26467 9503
rect 26617 9469 26651 9503
rect 26801 9469 26835 9503
rect 26985 9469 27019 9503
rect 29009 9469 29043 9503
rect 31125 9469 31159 9503
rect 6837 9401 6871 9435
rect 11437 9401 11471 9435
rect 12817 9401 12851 9435
rect 14381 9401 14415 9435
rect 17325 9401 17359 9435
rect 18153 9401 18187 9435
rect 25697 9401 25731 9435
rect 27169 9401 27203 9435
rect 28742 9401 28776 9435
rect 1409 9333 1443 9367
rect 6009 9333 6043 9367
rect 6745 9333 6779 9367
rect 11253 9333 11287 9367
rect 12909 9333 12943 9367
rect 17417 9333 17451 9367
rect 19441 9333 19475 9367
rect 27629 9333 27663 9367
rect 29561 9333 29595 9367
rect 31309 9333 31343 9367
rect 1961 9129 1995 9163
rect 2513 9129 2547 9163
rect 3801 9129 3835 9163
rect 5549 9129 5583 9163
rect 24225 9129 24259 9163
rect 29193 9129 29227 9163
rect 10885 9061 10919 9095
rect 11897 9061 11931 9095
rect 18889 9061 18923 9095
rect 23857 9061 23891 9095
rect 24073 9061 24107 9095
rect 28641 9061 28675 9095
rect 30297 9061 30331 9095
rect 1869 8993 1903 9027
rect 4445 8993 4479 9027
rect 4629 8993 4663 9027
rect 4813 8993 4847 9027
rect 4997 8993 5031 9027
rect 5457 8993 5491 9027
rect 5641 8993 5675 9027
rect 6377 8993 6411 9027
rect 6561 8993 6595 9027
rect 6929 8993 6963 9027
rect 7665 8993 7699 9027
rect 7932 8993 7966 9027
rect 9505 8993 9539 9027
rect 10149 8993 10183 9027
rect 10977 8993 11011 9027
rect 11713 8993 11747 9027
rect 12357 8993 12391 9027
rect 12633 8993 12667 9027
rect 12725 8993 12759 9027
rect 12817 8993 12851 9027
rect 13737 8993 13771 9027
rect 14197 8993 14231 9027
rect 16681 8993 16715 9027
rect 17693 8993 17727 9027
rect 21997 8993 22031 9027
rect 22661 8993 22695 9027
rect 22845 8993 22879 9027
rect 23213 8993 23247 9027
rect 25881 8993 25915 9027
rect 26157 8993 26191 9027
rect 26249 8993 26283 9027
rect 26433 8993 26467 9027
rect 27353 8993 27387 9027
rect 27537 8993 27571 9027
rect 27905 8993 27939 9027
rect 28549 8993 28583 9027
rect 4721 8925 4755 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 12541 8925 12575 8959
rect 17785 8925 17819 8959
rect 22201 8925 22235 8959
rect 22937 8925 22971 8959
rect 23029 8925 23063 8959
rect 26065 8925 26099 8959
rect 27629 8925 27663 8959
rect 27721 8925 27755 8959
rect 9045 8857 9079 8891
rect 9597 8857 9631 8891
rect 21281 8857 21315 8891
rect 28089 8857 28123 8891
rect 3157 8789 3191 8823
rect 4261 8789 4295 8823
rect 7113 8789 7147 8823
rect 10241 8789 10275 8823
rect 11529 8789 11563 8823
rect 13001 8789 13035 8823
rect 13645 8789 13679 8823
rect 15669 8789 15703 8823
rect 16773 8789 16807 8823
rect 17877 8789 17911 8823
rect 18061 8789 18095 8823
rect 20177 8789 20211 8823
rect 21833 8789 21867 8823
rect 23397 8789 23431 8823
rect 24041 8789 24075 8823
rect 24685 8789 24719 8823
rect 25697 8789 25731 8823
rect 29745 8789 29779 8823
rect 30849 8789 30883 8823
rect 5365 8585 5399 8619
rect 8401 8585 8435 8619
rect 10609 8585 10643 8619
rect 11805 8585 11839 8619
rect 12909 8585 12943 8619
rect 13461 8585 13495 8619
rect 14105 8585 14139 8619
rect 21373 8585 21407 8619
rect 24777 8585 24811 8619
rect 27353 8585 27387 8619
rect 28457 8585 28491 8619
rect 29561 8585 29595 8619
rect 2329 8517 2363 8551
rect 6469 8517 6503 8551
rect 18153 8517 18187 8551
rect 18429 8517 18463 8551
rect 23765 8517 23799 8551
rect 27905 8517 27939 8551
rect 30665 8517 30699 8551
rect 2513 8449 2547 8483
rect 11345 8449 11379 8483
rect 12541 8449 12575 8483
rect 12633 8449 12667 8483
rect 18061 8449 18095 8483
rect 19993 8449 20027 8483
rect 25421 8449 25455 8483
rect 26065 8449 26099 8483
rect 31217 8449 31251 8483
rect 1777 8381 1811 8415
rect 2237 8381 2271 8415
rect 2973 8381 3007 8415
rect 3157 8381 3191 8415
rect 3985 8381 4019 8415
rect 4252 8381 4286 8415
rect 7582 8381 7616 8415
rect 7849 8381 7883 8415
rect 9229 8381 9263 8415
rect 11069 8381 11103 8415
rect 11253 8381 11287 8415
rect 11437 8381 11471 8415
rect 11621 8381 11655 8415
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 12725 8381 12759 8415
rect 13369 8381 13403 8415
rect 15485 8381 15519 8415
rect 16313 8381 16347 8415
rect 16405 8381 16439 8415
rect 17785 8381 17819 8415
rect 17969 8381 18003 8415
rect 18245 8381 18279 8415
rect 19349 8381 19383 8415
rect 22385 8381 22419 8415
rect 25973 8381 26007 8415
rect 26157 8381 26191 8415
rect 26617 8381 26651 8415
rect 26801 8381 26835 8415
rect 26893 8381 26927 8415
rect 26985 8381 27019 8415
rect 27169 8381 27203 8415
rect 27813 8381 27847 8415
rect 1685 8313 1719 8347
rect 2513 8313 2547 8347
rect 9496 8313 9530 8347
rect 15218 8313 15252 8347
rect 17141 8313 17175 8347
rect 17325 8313 17359 8347
rect 20238 8313 20272 8347
rect 22652 8313 22686 8347
rect 25145 8313 25179 8347
rect 25237 8313 25271 8347
rect 30205 8313 30239 8347
rect 3065 8245 3099 8279
rect 5917 8245 5951 8279
rect 16957 8245 16991 8279
rect 19533 8245 19567 8279
rect 8309 8041 8343 8075
rect 9597 8041 9631 8075
rect 11529 8041 11563 8075
rect 22753 8041 22787 8075
rect 24593 8041 24627 8075
rect 25789 8041 25823 8075
rect 28273 8041 28307 8075
rect 30665 8041 30699 8075
rect 31217 8041 31251 8075
rect 12725 7973 12759 8007
rect 12909 7973 12943 8007
rect 13553 7973 13587 8007
rect 18337 7973 18371 8007
rect 19432 7973 19466 8007
rect 21097 7973 21131 8007
rect 23480 7973 23514 8007
rect 29386 7973 29420 8007
rect 2033 7905 2067 7939
rect 2145 7905 2179 7939
rect 2237 7908 2271 7942
rect 2421 7905 2455 7939
rect 3249 7905 3283 7939
rect 3893 7905 3927 7939
rect 5457 7905 5491 7939
rect 5641 7905 5675 7939
rect 6929 7905 6963 7939
rect 7481 7905 7515 7939
rect 8401 7905 8435 7939
rect 8861 7905 8895 7939
rect 9045 7905 9079 7939
rect 9413 7905 9447 7939
rect 10149 7905 10183 7939
rect 10425 7905 10459 7939
rect 10534 7905 10568 7939
rect 11713 7905 11747 7939
rect 11805 7905 11839 7939
rect 12081 7905 12115 7939
rect 13369 7905 13403 7939
rect 13737 7905 13771 7939
rect 15402 7905 15436 7939
rect 16681 7905 16715 7939
rect 16865 7905 16899 7939
rect 16957 7905 16991 7939
rect 17233 7905 17267 7939
rect 18245 7905 18279 7939
rect 22017 7905 22051 7939
rect 22201 7905 22235 7939
rect 22580 7905 22614 7939
rect 25421 7905 25455 7939
rect 25605 7905 25639 7939
rect 26249 7905 26283 7939
rect 27077 7905 27111 7939
rect 27261 7905 27295 7939
rect 27353 7905 27387 7939
rect 27629 7905 27663 7939
rect 30113 7905 30147 7939
rect 3525 7837 3559 7871
rect 4261 7837 4295 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 15669 7837 15703 7871
rect 17049 7837 17083 7871
rect 18061 7837 18095 7871
rect 19165 7837 19199 7871
rect 22293 7837 22327 7871
rect 22385 7837 22419 7871
rect 23213 7837 23247 7871
rect 26341 7837 26375 7871
rect 27445 7837 27479 7871
rect 29653 7837 29687 7871
rect 3709 7769 3743 7803
rect 6837 7769 6871 7803
rect 14289 7769 14323 7803
rect 20545 7769 20579 7803
rect 1777 7701 1811 7735
rect 4997 7701 5031 7735
rect 5641 7701 5675 7735
rect 7573 7701 7607 7735
rect 10241 7701 10275 7735
rect 10701 7701 10735 7735
rect 11989 7701 12023 7735
rect 12541 7701 12575 7735
rect 17417 7701 17451 7735
rect 18705 7701 18739 7735
rect 27813 7701 27847 7735
rect 1777 7497 1811 7531
rect 3985 7497 4019 7531
rect 4721 7497 4755 7531
rect 6837 7497 6871 7531
rect 8953 7497 8987 7531
rect 12265 7497 12299 7531
rect 14289 7497 14323 7531
rect 14473 7497 14507 7531
rect 14933 7497 14967 7531
rect 16129 7497 16163 7531
rect 16773 7497 16807 7531
rect 17233 7497 17267 7531
rect 19625 7497 19659 7531
rect 22753 7497 22787 7531
rect 24777 7497 24811 7531
rect 29561 7497 29595 7531
rect 30113 7497 30147 7531
rect 3157 7429 3191 7463
rect 3801 7429 3835 7463
rect 6101 7429 6135 7463
rect 1685 7361 1719 7395
rect 1869 7361 1903 7395
rect 2513 7361 2547 7395
rect 3249 7361 3283 7395
rect 5365 7361 5399 7395
rect 10977 7361 11011 7395
rect 11345 7361 11379 7395
rect 14197 7361 14231 7395
rect 15301 7361 15335 7395
rect 17785 7429 17819 7463
rect 18061 7429 18095 7463
rect 23305 7429 23339 7463
rect 25513 7429 25547 7463
rect 16313 7361 16347 7395
rect 18153 7361 18187 7395
rect 20361 7361 20395 7395
rect 26341 7361 26375 7395
rect 26617 7361 26651 7395
rect 1961 7293 1995 7327
rect 2605 7293 2639 7327
rect 2881 7293 2915 7327
rect 4629 7293 4663 7327
rect 5273 7293 5307 7327
rect 5549 7293 5583 7327
rect 5641 7293 5675 7327
rect 7941 7293 7975 7327
rect 9137 7293 9171 7327
rect 9321 7293 9355 7327
rect 9413 7293 9447 7327
rect 9505 7293 9539 7327
rect 9689 7293 9723 7327
rect 10609 7293 10643 7327
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 11161 7293 11195 7327
rect 11989 7293 12023 7327
rect 12357 7293 12391 7327
rect 12817 7293 12851 7327
rect 14105 7293 14139 7327
rect 15117 7293 15151 7327
rect 15393 7293 15427 7327
rect 15485 7293 15519 7327
rect 15669 7293 15703 7327
rect 16129 7293 16163 7327
rect 16221 7293 16255 7327
rect 16497 7293 16531 7327
rect 16589 7293 16623 7327
rect 17969 7293 18003 7327
rect 18245 7293 18279 7327
rect 18430 7293 18464 7327
rect 19257 7293 19291 7327
rect 19441 7293 19475 7327
rect 20085 7293 20119 7327
rect 21373 7293 21407 7327
rect 24777 7293 24811 7327
rect 25421 7293 25455 7327
rect 25605 7293 25639 7327
rect 25697 7293 25731 7327
rect 25881 7293 25915 7327
rect 28742 7293 28776 7327
rect 29009 7293 29043 7327
rect 31125 7293 31159 7327
rect 3969 7225 4003 7259
rect 4169 7225 4203 7259
rect 6883 7259 6917 7293
rect 6653 7225 6687 7259
rect 13001 7225 13035 7259
rect 21640 7225 21674 7259
rect 5273 7157 5307 7191
rect 5365 7157 5399 7191
rect 7021 7157 7055 7191
rect 8033 7157 8067 7191
rect 11805 7157 11839 7191
rect 13185 7157 13219 7191
rect 23765 7157 23799 7191
rect 25237 7157 25271 7191
rect 27629 7157 27663 7191
rect 31309 7157 31343 7191
rect 3525 6953 3559 6987
rect 5181 6953 5215 6987
rect 9505 6953 9539 6987
rect 17233 6953 17267 6987
rect 20085 6953 20119 6987
rect 22017 6953 22051 6987
rect 31309 6953 31343 6987
rect 3157 6885 3191 6919
rect 1685 6817 1719 6851
rect 1848 6817 1882 6851
rect 1961 6817 1995 6851
rect 2099 6817 2133 6851
rect 4445 6817 4479 6851
rect 4537 6817 4571 6851
rect 5457 6817 5491 6851
rect 5549 6817 5583 6851
rect 5641 6817 5675 6851
rect 5837 6817 5871 6851
rect 7297 6817 7331 6851
rect 10618 6817 10652 6851
rect 10885 6817 10919 6851
rect 11713 6817 11747 6851
rect 11897 6817 11931 6851
rect 12081 6817 12115 6851
rect 12265 6817 12299 6851
rect 12449 6817 12483 6851
rect 14022 6817 14056 6851
rect 15025 6817 15059 6851
rect 15209 6817 15243 6851
rect 15393 6817 15427 6851
rect 15577 6817 15611 6851
rect 15761 6817 15795 6851
rect 16865 6817 16899 6851
rect 17049 6817 17083 6851
rect 18061 6817 18095 6851
rect 18245 6817 18279 6851
rect 19349 6817 19383 6851
rect 19533 6817 19567 6851
rect 19993 6817 20027 6851
rect 20177 6817 20211 6851
rect 20637 6817 20671 6851
rect 22201 6817 22235 6851
rect 22477 6817 22511 6851
rect 22569 6817 22603 6851
rect 22753 6817 22787 6851
rect 23673 6817 23707 6851
rect 24685 6817 24719 6851
rect 25145 6817 25179 6851
rect 25329 6817 25363 6851
rect 25605 6817 25639 6851
rect 25789 6817 25823 6851
rect 26249 6817 26283 6851
rect 27169 6817 27203 6851
rect 27353 6817 27387 6851
rect 27721 6817 27755 6851
rect 29009 6817 29043 6851
rect 30573 6817 30607 6851
rect 31125 6817 31159 6851
rect 2329 6749 2363 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 4721 6749 4755 6783
rect 11989 6749 12023 6783
rect 14289 6749 14323 6783
rect 15485 6749 15519 6783
rect 18429 6749 18463 6783
rect 22385 6749 22419 6783
rect 24593 6749 24627 6783
rect 25513 6749 25547 6783
rect 26341 6749 26375 6783
rect 27445 6749 27479 6783
rect 27537 6749 27571 6783
rect 6377 6681 6411 6715
rect 8585 6681 8619 6715
rect 24317 6681 24351 6715
rect 25421 6681 25455 6715
rect 30021 6681 30055 6715
rect 4629 6613 4663 6647
rect 12909 6613 12943 6647
rect 20729 6613 20763 6647
rect 23765 6613 23799 6647
rect 24685 6613 24719 6647
rect 27905 6613 27939 6647
rect 28365 6613 28399 6647
rect 29469 6613 29503 6647
rect 2973 6409 3007 6443
rect 3985 6409 4019 6443
rect 11437 6409 11471 6443
rect 13277 6409 13311 6443
rect 14105 6409 14139 6443
rect 15945 6409 15979 6443
rect 16589 6409 16623 6443
rect 17509 6409 17543 6443
rect 18705 6409 18739 6443
rect 27077 6409 27111 6443
rect 29561 6409 29595 6443
rect 30113 6409 30147 6443
rect 30941 6409 30975 6443
rect 2053 6341 2087 6375
rect 5917 6341 5951 6375
rect 7113 6341 7147 6375
rect 8401 6341 8435 6375
rect 20729 6341 20763 6375
rect 5365 6273 5399 6307
rect 6929 6273 6963 6307
rect 7665 6273 7699 6307
rect 10517 6273 10551 6307
rect 14565 6273 14599 6307
rect 19901 6273 19935 6307
rect 22109 6273 22143 6307
rect 22845 6273 22879 6307
rect 23765 6273 23799 6307
rect 24409 6273 24443 6307
rect 26525 6273 26559 6307
rect 4077 6205 4111 6239
rect 4537 6205 4571 6239
rect 4721 6205 4755 6239
rect 5549 6205 5583 6239
rect 6653 6205 6687 6239
rect 7297 6205 7331 6239
rect 8953 6205 8987 6239
rect 9137 6205 9171 6239
rect 9223 6205 9257 6239
rect 9321 6205 9355 6239
rect 9516 6205 9550 6239
rect 9689 6205 9723 6239
rect 10149 6205 10183 6239
rect 10333 6205 10367 6239
rect 10425 6205 10459 6239
rect 10701 6205 10735 6239
rect 12449 6205 12483 6239
rect 12725 6205 12759 6239
rect 13185 6205 13219 6239
rect 14289 6205 14323 6239
rect 14473 6205 14507 6239
rect 14657 6205 14691 6239
rect 14841 6205 14875 6239
rect 16037 6205 16071 6239
rect 16681 6205 16715 6239
rect 17141 6205 17175 6239
rect 17969 6205 18003 6239
rect 19533 6205 19567 6239
rect 19717 6205 19751 6239
rect 19809 6205 19843 6239
rect 20085 6205 20119 6239
rect 21833 6205 21867 6239
rect 22569 6205 22603 6239
rect 22753 6205 22787 6239
rect 22937 6205 22971 6239
rect 23121 6205 23155 6239
rect 24685 6205 24719 6239
rect 26249 6205 26283 6239
rect 26341 6205 26375 6239
rect 26617 6205 26651 6239
rect 27629 6205 27663 6239
rect 27896 6205 27930 6239
rect 1869 6137 1903 6171
rect 2881 6137 2915 6171
rect 17325 6137 17359 6171
rect 18061 6137 18095 6171
rect 4629 6069 4663 6103
rect 5457 6069 5491 6103
rect 10885 6069 10919 6103
rect 15301 6069 15335 6103
rect 20269 6069 20303 6103
rect 23305 6069 23339 6103
rect 26065 6069 26099 6103
rect 29009 6069 29043 6103
rect 1593 5865 1627 5899
rect 2881 5865 2915 5899
rect 3433 5865 3467 5899
rect 5181 5865 5215 5899
rect 7205 5865 7239 5899
rect 9137 5865 9171 5899
rect 10977 5865 11011 5899
rect 16773 5865 16807 5899
rect 19073 5865 19107 5899
rect 22109 5865 22143 5899
rect 22661 5865 22695 5899
rect 24501 5865 24535 5899
rect 25697 5865 25731 5899
rect 27721 5865 27755 5899
rect 28365 5865 28399 5899
rect 29009 5865 29043 5899
rect 30573 5865 30607 5899
rect 31125 5865 31159 5899
rect 2237 5797 2271 5831
rect 8024 5797 8058 5831
rect 16957 5797 16991 5831
rect 23774 5797 23808 5831
rect 1501 5729 1535 5763
rect 1685 5729 1719 5763
rect 2329 5729 2363 5763
rect 2973 5729 3007 5763
rect 4169 5729 4203 5763
rect 4445 5729 4479 5763
rect 4537 5729 4571 5763
rect 4721 5729 4755 5763
rect 5457 5729 5491 5763
rect 5562 5729 5596 5763
rect 5662 5732 5696 5766
rect 5825 5729 5859 5763
rect 6377 5729 6411 5763
rect 6653 5729 6687 5763
rect 7113 5729 7147 5763
rect 7757 5729 7791 5763
rect 9597 5729 9631 5763
rect 9689 5729 9723 5763
rect 10241 5729 10275 5763
rect 10425 5729 10459 5763
rect 10609 5729 10643 5763
rect 10793 5729 10827 5763
rect 11621 5729 11655 5763
rect 14022 5729 14056 5763
rect 15209 5729 15243 5763
rect 15485 5729 15519 5763
rect 15577 5729 15611 5763
rect 15761 5729 15795 5763
rect 17141 5729 17175 5763
rect 17785 5729 17819 5763
rect 18153 5729 18187 5763
rect 20186 5729 20220 5763
rect 21097 5729 21131 5763
rect 24041 5729 24075 5763
rect 24685 5729 24719 5763
rect 24961 5729 24995 5763
rect 25053 5729 25087 5763
rect 25237 5729 25271 5763
rect 25881 5729 25915 5763
rect 26065 5729 26099 5763
rect 26261 5727 26295 5761
rect 26433 5729 26467 5763
rect 27169 5729 27203 5763
rect 27629 5729 27663 5763
rect 28457 5729 28491 5763
rect 4353 5661 4387 5695
rect 6745 5661 6779 5695
rect 10517 5661 10551 5695
rect 11897 5661 11931 5695
rect 14289 5661 14323 5695
rect 15393 5661 15427 5695
rect 20453 5661 20487 5695
rect 24869 5661 24903 5695
rect 26163 5661 26197 5695
rect 27077 5661 27111 5695
rect 17601 5593 17635 5627
rect 29469 5593 29503 5627
rect 30021 5593 30055 5627
rect 3985 5525 4019 5559
rect 12909 5525 12943 5559
rect 15025 5525 15059 5559
rect 17785 5525 17819 5559
rect 21005 5525 21039 5559
rect 3065 5321 3099 5355
rect 5181 5321 5215 5355
rect 17233 5321 17267 5355
rect 18705 5321 18739 5355
rect 19257 5321 19291 5355
rect 25605 5321 25639 5355
rect 28181 5321 28215 5355
rect 28733 5321 28767 5355
rect 29653 5321 29687 5355
rect 30665 5321 30699 5355
rect 9137 5253 9171 5287
rect 7481 5185 7515 5219
rect 10241 5185 10275 5219
rect 10977 5185 11011 5219
rect 12909 5185 12943 5219
rect 13001 5185 13035 5219
rect 16773 5185 16807 5219
rect 16865 5185 16899 5219
rect 18239 5185 18273 5219
rect 22109 5185 22143 5219
rect 22569 5185 22603 5219
rect 22845 5185 22879 5219
rect 24777 5185 24811 5219
rect 25973 5185 26007 5219
rect 27270 5185 27304 5219
rect 1685 5117 1719 5151
rect 3801 5117 3835 5151
rect 4068 5117 4102 5151
rect 7941 5117 7975 5151
rect 9229 5117 9263 5151
rect 10517 5117 10551 5151
rect 11253 5117 11287 5151
rect 12633 5117 12667 5151
rect 12817 5117 12851 5151
rect 13185 5117 13219 5151
rect 14381 5117 14415 5151
rect 16497 5117 16531 5151
rect 16681 5117 16715 5151
rect 17049 5117 17083 5151
rect 17969 5117 18003 5151
rect 18153 5117 18187 5151
rect 18383 5117 18417 5151
rect 18521 5117 18555 5151
rect 19257 5117 19291 5151
rect 19349 5117 19383 5151
rect 19625 5117 19659 5151
rect 24593 5117 24627 5151
rect 24869 5117 24903 5151
rect 24961 5117 24995 5151
rect 25145 5117 25179 5151
rect 25789 5117 25823 5151
rect 26065 5117 26099 5151
rect 26157 5117 26191 5151
rect 26341 5117 26375 5151
rect 26985 5117 27019 5151
rect 27169 5117 27203 5151
rect 27353 5117 27387 5151
rect 27537 5117 27571 5151
rect 31125 5117 31159 5151
rect 1930 5049 1964 5083
rect 7214 5049 7248 5083
rect 14648 5049 14682 5083
rect 21842 5049 21876 5083
rect 6101 4981 6135 5015
rect 8125 4981 8159 5015
rect 13369 4981 13403 5015
rect 15761 4981 15795 5015
rect 20729 4981 20763 5015
rect 24409 4981 24443 5015
rect 27721 4981 27755 5015
rect 31309 4981 31343 5015
rect 1961 4777 1995 4811
rect 2605 4777 2639 4811
rect 3065 4777 3099 4811
rect 3709 4777 3743 4811
rect 7113 4777 7147 4811
rect 9045 4777 9079 4811
rect 12265 4777 12299 4811
rect 14381 4777 14415 4811
rect 19441 4777 19475 4811
rect 21833 4777 21867 4811
rect 23029 4777 23063 4811
rect 27077 4777 27111 4811
rect 27629 4777 27663 4811
rect 29929 4777 29963 4811
rect 31033 4777 31067 4811
rect 1869 4709 1903 4743
rect 18153 4709 18187 4743
rect 28742 4709 28776 4743
rect 30481 4709 30515 4743
rect 4629 4641 4663 4675
rect 4813 4641 4847 4675
rect 4997 4641 5031 4675
rect 5181 4641 5215 4675
rect 6377 4641 6411 4675
rect 6561 4641 6595 4675
rect 6745 4641 6779 4675
rect 6929 4641 6963 4675
rect 7665 4641 7699 4675
rect 7932 4641 7966 4675
rect 10609 4641 10643 4675
rect 11529 4641 11563 4675
rect 11713 4641 11747 4675
rect 11897 4641 11931 4675
rect 12081 4641 12115 4675
rect 12909 4641 12943 4675
rect 13093 4641 13127 4675
rect 13277 4641 13311 4675
rect 13461 4641 13495 4675
rect 15494 4641 15528 4675
rect 15761 4641 15795 4675
rect 17509 4641 17543 4675
rect 18705 4641 18739 4675
rect 18889 4641 18923 4675
rect 18981 4641 19015 4675
rect 19257 4641 19291 4675
rect 19901 4641 19935 4675
rect 20168 4641 20202 4675
rect 22017 4641 22051 4675
rect 22385 4641 22419 4675
rect 22569 4641 22603 4675
rect 24153 4641 24187 4675
rect 24409 4641 24443 4675
rect 24869 4641 24903 4675
rect 26157 4641 26191 4675
rect 27169 4641 27203 4675
rect 29009 4641 29043 4675
rect 4905 4573 4939 4607
rect 5733 4573 5767 4607
rect 6653 4573 6687 4607
rect 10333 4573 10367 4607
rect 11805 4573 11839 4607
rect 13185 4573 13219 4607
rect 17233 4573 17267 4607
rect 19073 4573 19107 4607
rect 22201 4573 22235 4607
rect 22293 4573 22327 4607
rect 25145 4573 25179 4607
rect 17969 4505 18003 4539
rect 26249 4505 26283 4539
rect 4445 4437 4479 4471
rect 12725 4437 12759 4471
rect 21281 4437 21315 4471
rect 1685 4233 1719 4267
rect 4445 4233 4479 4267
rect 7021 4233 7055 4267
rect 13461 4233 13495 4267
rect 14197 4233 14231 4267
rect 15485 4233 15519 4267
rect 20637 4233 20671 4267
rect 22477 4233 22511 4267
rect 28089 4233 28123 4267
rect 3801 4097 3835 4131
rect 5825 4097 5859 4131
rect 8309 4097 8343 4131
rect 9137 4097 9171 4131
rect 9505 4097 9539 4131
rect 9597 4097 9631 4131
rect 12541 4097 12575 4131
rect 14657 4097 14691 4131
rect 15853 4097 15887 4131
rect 15945 4097 15979 4131
rect 16681 4097 16715 4131
rect 17141 4097 17175 4131
rect 17969 4097 18003 4131
rect 18061 4097 18095 4131
rect 18429 4097 18463 4131
rect 19533 4097 19567 4131
rect 23765 4097 23799 4131
rect 27537 4097 27571 4131
rect 28549 4097 28583 4131
rect 29653 4097 29687 4131
rect 30205 4097 30239 4131
rect 30941 4097 30975 4131
rect 2329 4029 2363 4063
rect 5558 4029 5592 4063
rect 7757 4029 7791 4063
rect 8401 4029 8435 4063
rect 9321 4029 9355 4063
rect 9689 4029 9723 4063
rect 9873 4029 9907 4063
rect 10517 4029 10551 4063
rect 10977 4029 11011 4063
rect 12265 4029 12299 4063
rect 12449 4029 12483 4063
rect 12633 4029 12667 4063
rect 12817 4029 12851 4063
rect 14105 4029 14139 4063
rect 14381 4029 14415 4063
rect 14473 4029 14507 4063
rect 15669 4029 15703 4063
rect 16037 4029 16071 4063
rect 16221 4029 16255 4063
rect 16865 4029 16899 4063
rect 16957 4029 16991 4063
rect 17233 4029 17267 4063
rect 17693 4029 17727 4063
rect 17877 4029 17911 4063
rect 18245 4029 18279 4063
rect 19073 4029 19107 4063
rect 19257 4029 19291 4063
rect 20545 4029 20579 4063
rect 21189 4029 21223 4063
rect 23673 4029 23707 4063
rect 24593 4029 24627 4063
rect 24869 4029 24903 4063
rect 28273 4029 28307 4063
rect 28365 4029 28399 4063
rect 28641 4029 28675 4063
rect 2881 3961 2915 3995
rect 10425 3961 10459 3995
rect 25881 3961 25915 3995
rect 6561 3893 6595 3927
rect 7665 3893 7699 3927
rect 11207 3893 11241 3927
rect 13001 3893 13035 3927
rect 19073 3893 19107 3927
rect 2881 3689 2915 3723
rect 3893 3689 3927 3723
rect 4445 3689 4479 3723
rect 5733 3689 5767 3723
rect 6469 3689 6503 3723
rect 7941 3689 7975 3723
rect 11529 3689 11563 3723
rect 15669 3689 15703 3723
rect 17693 3689 17727 3723
rect 19441 3689 19475 3723
rect 27169 3689 27203 3723
rect 30573 3689 30607 3723
rect 5089 3621 5123 3655
rect 7481 3621 7515 3655
rect 14534 3621 14568 3655
rect 29653 3621 29687 3655
rect 1869 3553 1903 3587
rect 9065 3553 9099 3587
rect 9321 3553 9355 3587
rect 9965 3553 9999 3587
rect 10241 3553 10275 3587
rect 10333 3553 10367 3587
rect 10517 3553 10551 3587
rect 12081 3553 12115 3587
rect 16681 3553 16715 3587
rect 17877 3553 17911 3587
rect 17969 3553 18003 3587
rect 18245 3553 18279 3587
rect 18889 3553 18923 3587
rect 18981 3553 19015 3587
rect 19441 3553 19475 3587
rect 19533 3553 19567 3587
rect 19717 3553 19751 3587
rect 19809 3553 19843 3587
rect 20085 3553 20119 3587
rect 22385 3553 22419 3587
rect 23857 3553 23891 3587
rect 24593 3553 24627 3587
rect 24961 3553 24995 3587
rect 25145 3553 25179 3587
rect 25605 3553 25639 3587
rect 25789 3553 25823 3587
rect 26157 3553 26191 3587
rect 27077 3553 27111 3587
rect 27721 3553 27755 3587
rect 27977 3553 28011 3587
rect 31125 3553 31159 3587
rect 2145 3485 2179 3519
rect 9781 3485 9815 3519
rect 10149 3485 10183 3519
rect 13829 3485 13863 3519
rect 14289 3485 14323 3519
rect 18153 3485 18187 3519
rect 19901 3485 19935 3519
rect 20269 3485 20303 3519
rect 23581 3485 23615 3519
rect 24777 3485 24811 3519
rect 24869 3485 24903 3519
rect 25881 3485 25915 3519
rect 25973 3485 26007 3519
rect 16773 3349 16807 3383
rect 20729 3349 20763 3383
rect 22293 3349 22327 3383
rect 24409 3349 24443 3383
rect 26341 3349 26375 3383
rect 29101 3349 29135 3383
rect 31309 3349 31343 3383
rect 2697 3145 2731 3179
rect 3157 3145 3191 3179
rect 3801 3145 3835 3179
rect 4353 3145 4387 3179
rect 5549 3145 5583 3179
rect 6101 3145 6135 3179
rect 7297 3145 7331 3179
rect 8401 3145 8435 3179
rect 9321 3145 9355 3179
rect 11621 3145 11655 3179
rect 12173 3145 12207 3179
rect 15945 3145 15979 3179
rect 16773 3145 16807 3179
rect 17417 3145 17451 3179
rect 19349 3145 19383 3179
rect 26525 3145 26559 3179
rect 29653 3145 29687 3179
rect 30113 3145 30147 3179
rect 31033 3145 31067 3179
rect 1501 3077 1535 3111
rect 22201 3077 22235 3111
rect 5089 3009 5123 3043
rect 6837 3009 6871 3043
rect 10149 3009 10183 3043
rect 13553 3009 13587 3043
rect 14565 3009 14599 3043
rect 17969 3009 18003 3043
rect 18429 3009 18463 3043
rect 24777 3009 24811 3043
rect 24869 3009 24903 3043
rect 26065 3009 26099 3043
rect 28641 3009 28675 3043
rect 9413 2941 9447 2975
rect 9873 2941 9907 2975
rect 10057 2941 10091 2975
rect 10241 2941 10275 2975
rect 10436 2941 10470 2975
rect 11713 2941 11747 2975
rect 13286 2941 13320 2975
rect 16865 2941 16899 2975
rect 17325 2941 17359 2975
rect 18153 2941 18187 2975
rect 18337 2941 18371 2975
rect 18521 2941 18555 2975
rect 18705 2941 18739 2975
rect 19257 2941 19291 2975
rect 21465 2941 21499 2975
rect 23397 2941 23431 2975
rect 23673 2941 23707 2975
rect 24593 2941 24627 2975
rect 24961 2941 24995 2975
rect 25145 2941 25179 2975
rect 25789 2941 25823 2975
rect 25973 2941 26007 2975
rect 26157 2941 26191 2975
rect 26341 2941 26375 2975
rect 26985 2941 27019 2975
rect 28457 2941 28491 2975
rect 28724 2941 28758 2975
rect 28825 2941 28859 2975
rect 29009 2941 29043 2975
rect 29561 2941 29595 2975
rect 29837 2941 29871 2975
rect 29929 2941 29963 2975
rect 2145 2873 2179 2907
rect 14832 2873 14866 2907
rect 21198 2873 21232 2907
rect 22017 2873 22051 2907
rect 10609 2805 10643 2839
rect 20085 2805 20119 2839
rect 24409 2805 24443 2839
rect 27215 2805 27249 2839
rect 28273 2805 28307 2839
rect 1593 2601 1627 2635
rect 2697 2601 2731 2635
rect 3249 2601 3283 2635
rect 4169 2601 4203 2635
rect 5641 2601 5675 2635
rect 6377 2601 6411 2635
rect 7389 2601 7423 2635
rect 8401 2601 8435 2635
rect 12725 2601 12759 2635
rect 14197 2601 14231 2635
rect 16681 2601 16715 2635
rect 23213 2601 23247 2635
rect 23765 2601 23799 2635
rect 29561 2601 29595 2635
rect 30389 2601 30423 2635
rect 9536 2533 9570 2567
rect 10241 2533 10275 2567
rect 22100 2533 22134 2567
rect 9781 2465 9815 2499
rect 10425 2465 10459 2499
rect 10793 2465 10827 2499
rect 10977 2465 11011 2499
rect 11529 2465 11563 2499
rect 11713 2465 11747 2499
rect 12081 2465 12115 2499
rect 13645 2465 13679 2499
rect 14105 2465 14139 2499
rect 15016 2465 15050 2499
rect 16865 2465 16899 2499
rect 17049 2465 17083 2499
rect 17141 2465 17175 2499
rect 17233 2465 17267 2499
rect 17413 2465 17447 2499
rect 17877 2465 17911 2499
rect 18061 2465 18095 2499
rect 18245 2465 18279 2499
rect 18429 2465 18463 2499
rect 19073 2465 19107 2499
rect 19257 2465 19291 2499
rect 19349 2465 19383 2499
rect 19441 2465 19475 2499
rect 19625 2465 19659 2499
rect 21833 2465 21867 2499
rect 24889 2465 24923 2499
rect 25145 2465 25179 2499
rect 25605 2465 25639 2499
rect 26985 2465 27019 2499
rect 27261 2465 27295 2499
rect 28273 2465 28307 2499
rect 28457 2465 28491 2499
rect 28549 2465 28583 2499
rect 28825 2465 28859 2499
rect 29469 2465 29503 2499
rect 10609 2397 10643 2431
rect 10701 2397 10735 2431
rect 11805 2397 11839 2431
rect 11897 2397 11931 2431
rect 14749 2397 14783 2431
rect 18153 2397 18187 2431
rect 21005 2397 21039 2431
rect 21281 2397 21315 2431
rect 25881 2397 25915 2431
rect 28641 2397 28675 2431
rect 16129 2329 16163 2363
rect 30849 2329 30883 2363
rect 12265 2261 12299 2295
rect 13553 2261 13587 2295
rect 18613 2261 18647 2295
rect 19809 2261 19843 2295
rect 29009 2261 29043 2295
rect 1501 2057 1535 2091
rect 2513 2057 2547 2091
rect 3157 2057 3191 2091
rect 3801 2057 3835 2091
rect 6009 2057 6043 2091
rect 9597 2057 9631 2091
rect 12725 2057 12759 2091
rect 13277 2057 13311 2091
rect 16773 2057 16807 2091
rect 19625 2057 19659 2091
rect 22845 2057 22879 2091
rect 23305 2057 23339 2091
rect 24409 2057 24443 2091
rect 26341 2057 26375 2091
rect 28457 2057 28491 2091
rect 29009 2057 29043 2091
rect 2053 1989 2087 2023
rect 6837 1989 6871 2023
rect 7389 1989 7423 2023
rect 8401 1989 8435 2023
rect 9045 1989 9079 2023
rect 10609 1989 10643 2023
rect 15669 1989 15703 2023
rect 14105 1921 14139 1955
rect 25789 1921 25823 1955
rect 11989 1853 12023 1887
rect 14381 1853 14415 1887
rect 16681 1853 16715 1887
rect 18449 1853 18483 1887
rect 18705 1853 18739 1887
rect 21005 1853 21039 1887
rect 21465 1853 21499 1887
rect 25533 1853 25567 1887
rect 26249 1853 26283 1887
rect 27077 1853 27111 1887
rect 11744 1785 11778 1819
rect 20738 1785 20772 1819
rect 21732 1785 21766 1819
rect 27344 1785 27378 1819
rect 29561 1785 29595 1819
rect 30113 1785 30147 1819
rect 10149 1717 10183 1751
rect 17325 1717 17359 1751
rect 30941 1717 30975 1751
rect 8033 1513 8067 1547
rect 8585 1513 8619 1547
rect 9137 1513 9171 1547
rect 9597 1513 9631 1547
rect 12725 1513 12759 1547
rect 14565 1513 14599 1547
rect 16773 1513 16807 1547
rect 18889 1513 18923 1547
rect 21833 1513 21867 1547
rect 24501 1513 24535 1547
rect 29009 1513 29043 1547
rect 29469 1513 29503 1547
rect 30021 1513 30055 1547
rect 10710 1445 10744 1479
rect 20002 1445 20036 1479
rect 1869 1377 1903 1411
rect 10977 1377 11011 1411
rect 13452 1377 13486 1411
rect 15577 1377 15611 1411
rect 15945 1377 15979 1411
rect 16129 1377 16163 1411
rect 17886 1377 17920 1411
rect 22937 1377 22971 1411
rect 23305 1377 23339 1411
rect 23489 1377 23523 1411
rect 24409 1377 24443 1411
rect 26166 1377 26200 1411
rect 26433 1377 26467 1411
rect 28190 1377 28224 1411
rect 31125 1377 31159 1411
rect 2789 1309 2823 1343
rect 13185 1309 13219 1343
rect 15393 1309 15427 1343
rect 15761 1309 15795 1343
rect 15853 1309 15887 1343
rect 18153 1309 18187 1343
rect 20269 1309 20303 1343
rect 22753 1309 22787 1343
rect 23121 1309 23155 1343
rect 23213 1309 23247 1343
rect 28457 1309 28491 1343
rect 2145 1241 2179 1275
rect 11621 1241 11655 1275
rect 12081 1173 12115 1207
rect 20729 1173 20763 1207
rect 25053 1173 25087 1207
rect 27077 1173 27111 1207
rect 31309 1173 31343 1207
rect 1593 969 1627 1003
rect 8401 969 8435 1003
rect 10425 969 10459 1003
rect 15301 969 15335 1003
rect 16037 969 16071 1003
rect 17509 969 17543 1003
rect 18061 969 18095 1003
rect 18613 969 18647 1003
rect 19441 969 19475 1003
rect 20729 969 20763 1003
rect 21833 969 21867 1003
rect 22385 969 22419 1003
rect 27629 969 27663 1003
rect 28089 969 28123 1003
rect 28733 969 28767 1003
rect 7849 901 7883 935
rect 11805 901 11839 935
rect 14105 901 14139 935
rect 21189 901 21223 935
rect 23029 901 23063 935
rect 23489 901 23523 935
rect 25513 901 25547 935
rect 29561 901 29595 935
rect 13185 833 13219 867
rect 17049 833 17083 867
rect 17141 833 17175 867
rect 25973 833 26007 867
rect 27077 833 27111 867
rect 9413 765 9447 799
rect 12918 765 12952 799
rect 14289 765 14323 799
rect 15945 765 15979 799
rect 16773 765 16807 799
rect 16957 765 16991 799
rect 17325 765 17359 799
rect 19625 765 19659 799
rect 24777 765 24811 799
rect 24961 765 24995 799
rect 25697 765 25731 799
rect 25835 765 25869 799
rect 26061 765 26095 799
rect 26249 765 26283 799
rect 7297 697 7331 731
rect 30113 697 30147 731
rect 9505 629 9539 663
rect 10977 629 11011 663
rect 20177 629 20211 663
<< metal1 >>
rect 1104 48442 32016 48464
rect 1104 48390 11253 48442
rect 11305 48390 11317 48442
rect 11369 48390 11381 48442
rect 11433 48390 11445 48442
rect 11497 48390 11509 48442
rect 11561 48390 21557 48442
rect 21609 48390 21621 48442
rect 21673 48390 21685 48442
rect 21737 48390 21749 48442
rect 21801 48390 21813 48442
rect 21865 48390 32016 48442
rect 1104 48368 32016 48390
rect 1397 48195 1455 48201
rect 1397 48161 1409 48195
rect 1443 48161 1455 48195
rect 1397 48155 1455 48161
rect 0 47988 800 48002
rect 1412 47988 1440 48155
rect 8478 48152 8484 48204
rect 8536 48192 8542 48204
rect 9125 48195 9183 48201
rect 9125 48192 9137 48195
rect 8536 48164 9137 48192
rect 8536 48152 8542 48164
rect 9125 48161 9137 48164
rect 9171 48161 9183 48195
rect 15838 48192 15844 48204
rect 15799 48164 15844 48192
rect 9125 48155 9183 48161
rect 15838 48152 15844 48164
rect 15896 48152 15902 48204
rect 24762 48152 24768 48204
rect 24820 48192 24826 48204
rect 25133 48195 25191 48201
rect 25133 48192 25145 48195
rect 24820 48164 25145 48192
rect 24820 48152 24826 48164
rect 25133 48161 25145 48164
rect 25179 48161 25191 48195
rect 25133 48155 25191 48161
rect 31113 48195 31171 48201
rect 31113 48161 31125 48195
rect 31159 48192 31171 48195
rect 31294 48192 31300 48204
rect 31159 48164 31300 48192
rect 31159 48161 31171 48164
rect 31113 48155 31171 48161
rect 31294 48152 31300 48164
rect 31352 48152 31358 48204
rect 8294 48016 8300 48068
rect 8352 48056 8358 48068
rect 8941 48059 8999 48065
rect 8941 48056 8953 48059
rect 8352 48028 8953 48056
rect 8352 48016 8358 48028
rect 8941 48025 8953 48028
rect 8987 48025 8999 48059
rect 8941 48019 8999 48025
rect 14918 48016 14924 48068
rect 14976 48056 14982 48068
rect 15381 48059 15439 48065
rect 15381 48056 15393 48059
rect 14976 48028 15393 48056
rect 14976 48016 14982 48028
rect 15381 48025 15393 48028
rect 15427 48056 15439 48059
rect 15427 48028 18184 48056
rect 15427 48025 15439 48028
rect 15381 48019 15439 48025
rect 0 47960 1440 47988
rect 1581 47991 1639 47997
rect 0 47946 800 47960
rect 1044 47784 1072 47960
rect 1581 47957 1593 47991
rect 1627 47988 1639 47991
rect 5718 47988 5724 48000
rect 1627 47960 5724 47988
rect 1627 47957 1639 47960
rect 1581 47951 1639 47957
rect 5718 47948 5724 47960
rect 5776 47948 5782 48000
rect 11606 47948 11612 48000
rect 11664 47988 11670 48000
rect 11701 47991 11759 47997
rect 11701 47988 11713 47991
rect 11664 47960 11713 47988
rect 11664 47948 11670 47960
rect 11701 47957 11713 47960
rect 11747 47957 11759 47991
rect 15930 47988 15936 48000
rect 15891 47960 15936 47988
rect 11701 47951 11759 47957
rect 15930 47948 15936 47960
rect 15988 47948 15994 48000
rect 16758 47948 16764 48000
rect 16816 47988 16822 48000
rect 18156 47997 18184 48028
rect 24854 48016 24860 48068
rect 24912 48056 24918 48068
rect 24949 48059 25007 48065
rect 24949 48056 24961 48059
rect 24912 48028 24961 48056
rect 24912 48016 24918 48028
rect 24949 48025 24961 48028
rect 24995 48025 25007 48059
rect 24949 48019 25007 48025
rect 16945 47991 17003 47997
rect 16945 47988 16957 47991
rect 16816 47960 16957 47988
rect 16816 47948 16822 47960
rect 16945 47957 16957 47960
rect 16991 47957 17003 47991
rect 16945 47951 17003 47957
rect 18141 47991 18199 47997
rect 18141 47957 18153 47991
rect 18187 47988 18199 47991
rect 19521 47991 19579 47997
rect 19521 47988 19533 47991
rect 18187 47960 19533 47988
rect 18187 47957 18199 47960
rect 18141 47951 18199 47957
rect 19521 47957 19533 47960
rect 19567 47988 19579 47991
rect 20070 47988 20076 48000
rect 19567 47960 20076 47988
rect 19567 47957 19579 47960
rect 19521 47951 19579 47957
rect 20070 47948 20076 47960
rect 20128 47948 20134 48000
rect 31297 47991 31355 47997
rect 31297 47957 31309 47991
rect 31343 47988 31355 47991
rect 32320 47988 33120 48002
rect 31343 47960 33120 47988
rect 31343 47957 31355 47960
rect 31297 47951 31355 47957
rect 32320 47946 33120 47960
rect 1104 47898 32016 47920
rect 1104 47846 6102 47898
rect 6154 47846 6166 47898
rect 6218 47846 6230 47898
rect 6282 47846 6294 47898
rect 6346 47846 6358 47898
rect 6410 47846 16405 47898
rect 16457 47846 16469 47898
rect 16521 47846 16533 47898
rect 16585 47846 16597 47898
rect 16649 47846 16661 47898
rect 16713 47846 26709 47898
rect 26761 47846 26773 47898
rect 26825 47846 26837 47898
rect 26889 47846 26901 47898
rect 26953 47846 26965 47898
rect 27017 47846 32016 47898
rect 1104 47824 32016 47846
rect 1397 47787 1455 47793
rect 1397 47784 1409 47787
rect 1044 47756 1409 47784
rect 1397 47753 1409 47756
rect 1443 47753 1455 47787
rect 1397 47747 1455 47753
rect 14185 47787 14243 47793
rect 14185 47753 14197 47787
rect 14231 47784 14243 47787
rect 18322 47784 18328 47796
rect 14231 47756 18328 47784
rect 14231 47753 14243 47756
rect 14185 47747 14243 47753
rect 18322 47744 18328 47756
rect 18380 47744 18386 47796
rect 11606 47676 11612 47728
rect 11664 47716 11670 47728
rect 14918 47716 14924 47728
rect 11664 47688 14924 47716
rect 11664 47676 11670 47688
rect 14918 47676 14924 47688
rect 14976 47676 14982 47728
rect 12894 47608 12900 47660
rect 12952 47648 12958 47660
rect 13265 47651 13323 47657
rect 13265 47648 13277 47651
rect 12952 47620 13277 47648
rect 12952 47608 12958 47620
rect 13265 47617 13277 47620
rect 13311 47617 13323 47651
rect 13265 47611 13323 47617
rect 8297 47583 8355 47589
rect 8297 47549 8309 47583
rect 8343 47580 8355 47583
rect 10410 47580 10416 47592
rect 8343 47552 10416 47580
rect 8343 47549 8355 47552
rect 8297 47543 8355 47549
rect 10410 47540 10416 47552
rect 10468 47580 10474 47592
rect 10505 47583 10563 47589
rect 10505 47580 10517 47583
rect 10468 47552 10517 47580
rect 10468 47540 10474 47552
rect 10505 47549 10517 47552
rect 10551 47549 10563 47583
rect 10505 47543 10563 47549
rect 12989 47583 13047 47589
rect 12989 47549 13001 47583
rect 13035 47549 13047 47583
rect 12989 47543 13047 47549
rect 8018 47512 8024 47524
rect 8076 47521 8082 47524
rect 7988 47484 8024 47512
rect 8018 47472 8024 47484
rect 8076 47475 8088 47521
rect 10772 47515 10830 47521
rect 10772 47481 10784 47515
rect 10818 47512 10830 47515
rect 10962 47512 10968 47524
rect 10818 47484 10968 47512
rect 10818 47481 10830 47484
rect 10772 47475 10830 47481
rect 8076 47472 8082 47475
rect 10962 47472 10968 47484
rect 11020 47472 11026 47524
rect 6914 47444 6920 47456
rect 6875 47416 6920 47444
rect 6914 47404 6920 47416
rect 6972 47404 6978 47456
rect 10870 47404 10876 47456
rect 10928 47444 10934 47456
rect 11885 47447 11943 47453
rect 11885 47444 11897 47447
rect 10928 47416 11897 47444
rect 10928 47404 10934 47416
rect 11885 47413 11897 47416
rect 11931 47413 11943 47447
rect 12802 47444 12808 47456
rect 12763 47416 12808 47444
rect 11885 47407 11943 47413
rect 12802 47404 12808 47416
rect 12860 47404 12866 47456
rect 13004 47444 13032 47543
rect 13078 47540 13084 47592
rect 13136 47580 13142 47592
rect 13173 47583 13231 47589
rect 13173 47580 13185 47583
rect 13136 47552 13185 47580
rect 13136 47540 13142 47552
rect 13173 47549 13185 47552
rect 13219 47549 13231 47583
rect 13173 47543 13231 47549
rect 13357 47583 13415 47589
rect 13357 47549 13369 47583
rect 13403 47549 13415 47583
rect 13357 47543 13415 47549
rect 13541 47583 13599 47589
rect 13541 47549 13553 47583
rect 13587 47580 13599 47583
rect 13722 47580 13728 47592
rect 13587 47552 13728 47580
rect 13587 47549 13599 47552
rect 13541 47543 13599 47549
rect 13372 47512 13400 47543
rect 13722 47540 13728 47552
rect 13780 47540 13786 47592
rect 14366 47540 14372 47592
rect 14424 47580 14430 47592
rect 15381 47583 15439 47589
rect 15381 47580 15393 47583
rect 14424 47552 15393 47580
rect 14424 47540 14430 47552
rect 15381 47549 15393 47552
rect 15427 47549 15439 47583
rect 15381 47543 15439 47549
rect 17313 47583 17371 47589
rect 17313 47549 17325 47583
rect 17359 47580 17371 47583
rect 18046 47580 18052 47592
rect 17359 47552 18052 47580
rect 17359 47549 17371 47552
rect 17313 47543 17371 47549
rect 18046 47540 18052 47552
rect 18104 47540 18110 47592
rect 21085 47583 21143 47589
rect 21085 47549 21097 47583
rect 21131 47580 21143 47583
rect 21821 47583 21879 47589
rect 21821 47580 21833 47583
rect 21131 47552 21833 47580
rect 21131 47549 21143 47552
rect 21085 47543 21143 47549
rect 21821 47549 21833 47552
rect 21867 47580 21879 47583
rect 21910 47580 21916 47592
rect 21867 47552 21916 47580
rect 21867 47549 21879 47552
rect 21821 47543 21879 47549
rect 21910 47540 21916 47552
rect 21968 47540 21974 47592
rect 13814 47512 13820 47524
rect 13372 47484 13820 47512
rect 13814 47472 13820 47484
rect 13872 47472 13878 47524
rect 15648 47515 15706 47521
rect 15648 47481 15660 47515
rect 15694 47512 15706 47515
rect 15746 47512 15752 47524
rect 15694 47484 15752 47512
rect 15694 47481 15706 47484
rect 15648 47475 15706 47481
rect 15746 47472 15752 47484
rect 15804 47472 15810 47524
rect 17580 47515 17638 47521
rect 17580 47481 17592 47515
rect 17626 47512 17638 47515
rect 17862 47512 17868 47524
rect 17626 47484 17868 47512
rect 17626 47481 17638 47484
rect 17580 47475 17638 47481
rect 17862 47472 17868 47484
rect 17920 47472 17926 47524
rect 20840 47515 20898 47521
rect 20840 47481 20852 47515
rect 20886 47512 20898 47515
rect 20990 47512 20996 47524
rect 20886 47484 20996 47512
rect 20886 47481 20898 47484
rect 20840 47475 20898 47481
rect 20990 47472 20996 47484
rect 21048 47472 21054 47524
rect 22088 47515 22146 47521
rect 22088 47481 22100 47515
rect 22134 47512 22146 47515
rect 22554 47512 22560 47524
rect 22134 47484 22560 47512
rect 22134 47481 22146 47484
rect 22088 47475 22146 47481
rect 22554 47472 22560 47484
rect 22612 47472 22618 47524
rect 13538 47444 13544 47456
rect 13004 47416 13544 47444
rect 13538 47404 13544 47416
rect 13596 47404 13602 47456
rect 16114 47404 16120 47456
rect 16172 47444 16178 47456
rect 16761 47447 16819 47453
rect 16761 47444 16773 47447
rect 16172 47416 16773 47444
rect 16172 47404 16178 47416
rect 16761 47413 16773 47416
rect 16807 47413 16819 47447
rect 16761 47407 16819 47413
rect 17678 47404 17684 47456
rect 17736 47444 17742 47456
rect 18693 47447 18751 47453
rect 18693 47444 18705 47447
rect 17736 47416 18705 47444
rect 17736 47404 17742 47416
rect 18693 47413 18705 47416
rect 18739 47413 18751 47447
rect 19702 47444 19708 47456
rect 19663 47416 19708 47444
rect 18693 47407 18751 47413
rect 19702 47404 19708 47416
rect 19760 47404 19766 47456
rect 22370 47404 22376 47456
rect 22428 47444 22434 47456
rect 23201 47447 23259 47453
rect 23201 47444 23213 47447
rect 22428 47416 23213 47444
rect 22428 47404 22434 47416
rect 23201 47413 23213 47416
rect 23247 47444 23259 47447
rect 24486 47444 24492 47456
rect 23247 47416 24492 47444
rect 23247 47413 23259 47416
rect 23201 47407 23259 47413
rect 24486 47404 24492 47416
rect 24544 47404 24550 47456
rect 1104 47354 32016 47376
rect 1104 47302 11253 47354
rect 11305 47302 11317 47354
rect 11369 47302 11381 47354
rect 11433 47302 11445 47354
rect 11497 47302 11509 47354
rect 11561 47302 21557 47354
rect 21609 47302 21621 47354
rect 21673 47302 21685 47354
rect 21737 47302 21749 47354
rect 21801 47302 21813 47354
rect 21865 47302 32016 47354
rect 1104 47280 32016 47302
rect 15378 47240 15384 47252
rect 15291 47212 15384 47240
rect 15378 47200 15384 47212
rect 15436 47240 15442 47252
rect 15838 47240 15844 47252
rect 15436 47212 15844 47240
rect 15436 47200 15442 47212
rect 15838 47200 15844 47212
rect 15896 47200 15902 47252
rect 22554 47240 22560 47252
rect 22515 47212 22560 47240
rect 22554 47200 22560 47212
rect 22612 47200 22618 47252
rect 24762 47240 24768 47252
rect 24723 47212 24768 47240
rect 24762 47200 24768 47212
rect 24820 47200 24826 47252
rect 31294 47240 31300 47252
rect 31255 47212 31300 47240
rect 31294 47200 31300 47212
rect 31352 47200 31358 47252
rect 10410 47172 10416 47184
rect 7760 47144 10416 47172
rect 7760 47116 7788 47144
rect 7742 47104 7748 47116
rect 7655 47076 7748 47104
rect 7742 47064 7748 47076
rect 7800 47064 7806 47116
rect 7834 47064 7840 47116
rect 7892 47104 7898 47116
rect 9600 47113 9628 47144
rect 10410 47132 10416 47144
rect 10468 47132 10474 47184
rect 12428 47175 12486 47181
rect 12428 47141 12440 47175
rect 12474 47172 12486 47175
rect 12802 47172 12808 47184
rect 12474 47144 12808 47172
rect 12474 47141 12486 47144
rect 12428 47135 12486 47141
rect 12802 47132 12808 47144
rect 12860 47132 12866 47184
rect 20714 47172 20720 47184
rect 18708 47144 20720 47172
rect 9858 47113 9864 47116
rect 8001 47107 8059 47113
rect 8001 47104 8013 47107
rect 7892 47076 8013 47104
rect 7892 47064 7898 47076
rect 8001 47073 8013 47076
rect 8047 47073 8059 47107
rect 8001 47067 8059 47073
rect 9585 47107 9643 47113
rect 9585 47073 9597 47107
rect 9631 47073 9643 47107
rect 9585 47067 9643 47073
rect 9852 47067 9864 47113
rect 9916 47104 9922 47116
rect 9916 47076 9952 47104
rect 9858 47064 9864 47067
rect 9916 47064 9922 47076
rect 13354 47064 13360 47116
rect 13412 47104 13418 47116
rect 14257 47107 14315 47113
rect 14257 47104 14269 47107
rect 13412 47076 14269 47104
rect 13412 47064 13418 47076
rect 14257 47073 14269 47076
rect 14303 47073 14315 47107
rect 16114 47104 16120 47116
rect 16075 47076 16120 47104
rect 14257 47067 14315 47073
rect 16114 47064 16120 47076
rect 16172 47064 16178 47116
rect 17402 47064 17408 47116
rect 17460 47104 17466 47116
rect 17782 47107 17840 47113
rect 17782 47104 17794 47107
rect 17460 47076 17794 47104
rect 17460 47064 17466 47076
rect 17782 47073 17794 47076
rect 17828 47073 17840 47107
rect 18046 47104 18052 47116
rect 17959 47076 18052 47104
rect 17782 47067 17840 47073
rect 18046 47064 18052 47076
rect 18104 47104 18110 47116
rect 18708 47113 18736 47144
rect 20714 47132 20720 47144
rect 20772 47132 20778 47184
rect 23652 47175 23710 47181
rect 23652 47141 23664 47175
rect 23698 47172 23710 47175
rect 23842 47172 23848 47184
rect 23698 47144 23848 47172
rect 23698 47141 23710 47144
rect 23652 47135 23710 47141
rect 23842 47132 23848 47144
rect 23900 47172 23906 47184
rect 25225 47175 25283 47181
rect 25225 47172 25237 47175
rect 23900 47144 25237 47172
rect 23900 47132 23906 47144
rect 25225 47141 25237 47144
rect 25271 47141 25283 47175
rect 25225 47135 25283 47141
rect 18693 47107 18751 47113
rect 18693 47104 18705 47107
rect 18104 47076 18705 47104
rect 18104 47064 18110 47076
rect 18693 47073 18705 47076
rect 18739 47073 18751 47107
rect 18693 47067 18751 47073
rect 18782 47064 18788 47116
rect 18840 47104 18846 47116
rect 18949 47107 19007 47113
rect 18949 47104 18961 47107
rect 18840 47076 18961 47104
rect 18840 47064 18846 47076
rect 18949 47073 18961 47076
rect 18995 47073 19007 47107
rect 18949 47067 19007 47073
rect 19702 47064 19708 47116
rect 19760 47104 19766 47116
rect 20162 47104 20168 47116
rect 19760 47076 20168 47104
rect 19760 47064 19766 47076
rect 20162 47064 20168 47076
rect 20220 47104 20226 47116
rect 21085 47107 21143 47113
rect 21085 47104 21097 47107
rect 20220 47076 21097 47104
rect 20220 47064 20226 47076
rect 21085 47073 21097 47076
rect 21131 47073 21143 47107
rect 21085 47067 21143 47073
rect 21450 47064 21456 47116
rect 21508 47104 21514 47116
rect 21821 47107 21879 47113
rect 21821 47104 21833 47107
rect 21508 47076 21833 47104
rect 21508 47064 21514 47076
rect 21821 47073 21833 47076
rect 21867 47073 21879 47107
rect 22002 47104 22008 47116
rect 21963 47076 22008 47104
rect 21821 47067 21879 47073
rect 22002 47064 22008 47076
rect 22060 47064 22066 47116
rect 22370 47104 22376 47116
rect 22331 47076 22376 47104
rect 22370 47064 22376 47076
rect 22428 47064 22434 47116
rect 30650 47064 30656 47116
rect 30708 47104 30714 47116
rect 31113 47107 31171 47113
rect 31113 47104 31125 47107
rect 30708 47076 31125 47104
rect 30708 47064 30714 47076
rect 31113 47073 31125 47076
rect 31159 47073 31171 47107
rect 31113 47067 31171 47073
rect 12158 47036 12164 47048
rect 12119 47008 12164 47036
rect 12158 46996 12164 47008
rect 12216 46996 12222 47048
rect 14001 47039 14059 47045
rect 14001 47005 14013 47039
rect 14047 47005 14059 47039
rect 14001 46999 14059 47005
rect 11606 46968 11612 46980
rect 11567 46940 11612 46968
rect 11606 46928 11612 46940
rect 11664 46928 11670 46980
rect 9125 46903 9183 46909
rect 9125 46869 9137 46903
rect 9171 46900 9183 46903
rect 9214 46900 9220 46912
rect 9171 46872 9220 46900
rect 9171 46869 9183 46872
rect 9125 46863 9183 46869
rect 9214 46860 9220 46872
rect 9272 46860 9278 46912
rect 10870 46860 10876 46912
rect 10928 46900 10934 46912
rect 10965 46903 11023 46909
rect 10965 46900 10977 46903
rect 10928 46872 10977 46900
rect 10928 46860 10934 46872
rect 10965 46869 10977 46872
rect 11011 46869 11023 46903
rect 13538 46900 13544 46912
rect 13499 46872 13544 46900
rect 10965 46863 11023 46869
rect 13538 46860 13544 46872
rect 13596 46860 13602 46912
rect 14016 46900 14044 46999
rect 21266 46996 21272 47048
rect 21324 47036 21330 47048
rect 22097 47039 22155 47045
rect 22097 47036 22109 47039
rect 21324 47008 22109 47036
rect 21324 46996 21330 47008
rect 22097 47005 22109 47008
rect 22143 47005 22155 47039
rect 22097 46999 22155 47005
rect 22189 47039 22247 47045
rect 22189 47005 22201 47039
rect 22235 47036 22247 47039
rect 22554 47036 22560 47048
rect 22235 47008 22560 47036
rect 22235 47005 22247 47008
rect 22189 46999 22247 47005
rect 22554 46996 22560 47008
rect 22612 46996 22618 47048
rect 23385 47039 23443 47045
rect 23385 47005 23397 47039
rect 23431 47005 23443 47039
rect 23385 46999 23443 47005
rect 16022 46968 16028 46980
rect 15983 46940 16028 46968
rect 16022 46928 16028 46940
rect 16080 46928 16086 46980
rect 20622 46968 20628 46980
rect 20583 46940 20628 46968
rect 20622 46928 20628 46940
rect 20680 46928 20686 46980
rect 21177 46971 21235 46977
rect 21177 46937 21189 46971
rect 21223 46968 21235 46971
rect 21358 46968 21364 46980
rect 21223 46940 21364 46968
rect 21223 46937 21235 46940
rect 21177 46931 21235 46937
rect 21358 46928 21364 46940
rect 21416 46928 21422 46980
rect 21910 46928 21916 46980
rect 21968 46968 21974 46980
rect 23400 46968 23428 46999
rect 21968 46940 23428 46968
rect 21968 46928 21974 46940
rect 14366 46900 14372 46912
rect 14016 46872 14372 46900
rect 14366 46860 14372 46872
rect 14424 46860 14430 46912
rect 16669 46903 16727 46909
rect 16669 46869 16681 46903
rect 16715 46900 16727 46903
rect 17310 46900 17316 46912
rect 16715 46872 17316 46900
rect 16715 46869 16727 46872
rect 16669 46863 16727 46869
rect 17310 46860 17316 46872
rect 17368 46860 17374 46912
rect 18966 46860 18972 46912
rect 19024 46900 19030 46912
rect 20073 46903 20131 46909
rect 20073 46900 20085 46903
rect 19024 46872 20085 46900
rect 19024 46860 19030 46872
rect 20073 46869 20085 46872
rect 20119 46900 20131 46903
rect 21082 46900 21088 46912
rect 20119 46872 21088 46900
rect 20119 46869 20131 46872
rect 20073 46863 20131 46869
rect 21082 46860 21088 46872
rect 21140 46860 21146 46912
rect 30650 46900 30656 46912
rect 30611 46872 30656 46900
rect 30650 46860 30656 46872
rect 30708 46860 30714 46912
rect 1104 46810 32016 46832
rect 1104 46758 6102 46810
rect 6154 46758 6166 46810
rect 6218 46758 6230 46810
rect 6282 46758 6294 46810
rect 6346 46758 6358 46810
rect 6410 46758 16405 46810
rect 16457 46758 16469 46810
rect 16521 46758 16533 46810
rect 16585 46758 16597 46810
rect 16649 46758 16661 46810
rect 16713 46758 26709 46810
rect 26761 46758 26773 46810
rect 26825 46758 26837 46810
rect 26889 46758 26901 46810
rect 26953 46758 26965 46810
rect 27017 46758 32016 46810
rect 1104 46736 32016 46758
rect 7834 46656 7840 46708
rect 7892 46696 7898 46708
rect 8389 46699 8447 46705
rect 8389 46696 8401 46699
rect 7892 46668 8401 46696
rect 7892 46656 7898 46668
rect 8389 46665 8401 46668
rect 8435 46665 8447 46699
rect 8389 46659 8447 46665
rect 13541 46699 13599 46705
rect 13541 46665 13553 46699
rect 13587 46696 13599 46699
rect 13814 46696 13820 46708
rect 13587 46668 13820 46696
rect 13587 46665 13599 46668
rect 13541 46659 13599 46665
rect 13814 46656 13820 46668
rect 13872 46656 13878 46708
rect 17862 46696 17868 46708
rect 17823 46668 17868 46696
rect 17862 46656 17868 46668
rect 17920 46656 17926 46708
rect 18322 46696 18328 46708
rect 18283 46668 18328 46696
rect 18322 46656 18328 46668
rect 18380 46656 18386 46708
rect 8036 46600 9536 46628
rect 6914 46520 6920 46572
rect 6972 46560 6978 46572
rect 8036 46569 8064 46600
rect 9508 46572 9536 46600
rect 23750 46588 23756 46640
rect 23808 46628 23814 46640
rect 23808 46600 24808 46628
rect 23808 46588 23814 46600
rect 8021 46563 8079 46569
rect 6972 46532 7880 46560
rect 6972 46520 6978 46532
rect 7852 46504 7880 46532
rect 8021 46529 8033 46563
rect 8067 46529 8079 46563
rect 9214 46560 9220 46572
rect 8021 46523 8079 46529
rect 8220 46532 9220 46560
rect 7282 46452 7288 46504
rect 7340 46492 7346 46504
rect 7653 46495 7711 46501
rect 7653 46492 7665 46495
rect 7340 46464 7665 46492
rect 7340 46452 7346 46464
rect 7653 46461 7665 46464
rect 7699 46461 7711 46495
rect 7834 46492 7840 46504
rect 7747 46464 7840 46492
rect 7653 46455 7711 46461
rect 7834 46452 7840 46464
rect 7892 46452 7898 46504
rect 8220 46501 8248 46532
rect 9214 46520 9220 46532
rect 9272 46520 9278 46572
rect 9490 46560 9496 46572
rect 9403 46532 9496 46560
rect 9490 46520 9496 46532
rect 9548 46520 9554 46572
rect 13538 46520 13544 46572
rect 13596 46560 13602 46572
rect 13596 46532 14504 46560
rect 13596 46520 13602 46532
rect 7929 46495 7987 46501
rect 7929 46461 7941 46495
rect 7975 46461 7987 46495
rect 7929 46455 7987 46461
rect 8205 46495 8263 46501
rect 8205 46461 8217 46495
rect 8251 46461 8263 46495
rect 8205 46455 8263 46461
rect 7558 46384 7564 46436
rect 7616 46424 7622 46436
rect 7944 46424 7972 46455
rect 9030 46452 9036 46504
rect 9088 46492 9094 46504
rect 9125 46495 9183 46501
rect 9125 46492 9137 46495
rect 9088 46464 9137 46492
rect 9088 46452 9094 46464
rect 9125 46461 9137 46464
rect 9171 46461 9183 46495
rect 9125 46455 9183 46461
rect 9309 46495 9367 46501
rect 9309 46461 9321 46495
rect 9355 46461 9367 46495
rect 9309 46455 9367 46461
rect 7616 46396 7972 46424
rect 9324 46424 9352 46455
rect 9398 46452 9404 46504
rect 9456 46492 9462 46504
rect 9674 46492 9680 46504
rect 9456 46464 9501 46492
rect 9635 46464 9680 46492
rect 9456 46452 9462 46464
rect 9674 46452 9680 46464
rect 9732 46452 9738 46504
rect 10321 46495 10379 46501
rect 10321 46461 10333 46495
rect 10367 46492 10379 46495
rect 10410 46492 10416 46504
rect 10367 46464 10416 46492
rect 10367 46461 10379 46464
rect 10321 46455 10379 46461
rect 10410 46452 10416 46464
rect 10468 46492 10474 46504
rect 12158 46492 12164 46504
rect 10468 46464 12164 46492
rect 10468 46452 10474 46464
rect 12158 46452 12164 46464
rect 12216 46452 12222 46504
rect 12802 46452 12808 46504
rect 12860 46492 12866 46504
rect 13556 46492 13584 46520
rect 14366 46492 14372 46504
rect 12860 46464 13584 46492
rect 14327 46464 14372 46492
rect 12860 46452 12866 46464
rect 14366 46452 14372 46464
rect 14424 46452 14430 46504
rect 14476 46492 14504 46532
rect 21910 46520 21916 46572
rect 21968 46560 21974 46572
rect 22465 46563 22523 46569
rect 22465 46560 22477 46563
rect 21968 46532 22477 46560
rect 21968 46520 21974 46532
rect 22465 46529 22477 46532
rect 22511 46529 22523 46563
rect 22465 46523 22523 46529
rect 23474 46520 23480 46572
rect 23532 46560 23538 46572
rect 24667 46563 24725 46569
rect 24667 46560 24679 46563
rect 23532 46532 24679 46560
rect 23532 46520 23538 46532
rect 24667 46529 24679 46532
rect 24713 46529 24725 46563
rect 24667 46523 24725 46529
rect 16209 46495 16267 46501
rect 16209 46492 16221 46495
rect 14476 46464 16221 46492
rect 16209 46461 16221 46464
rect 16255 46461 16267 46495
rect 16209 46455 16267 46461
rect 16666 46452 16672 46504
rect 16724 46492 16730 46504
rect 17126 46492 17132 46504
rect 16724 46464 17132 46492
rect 16724 46452 16730 46464
rect 17126 46452 17132 46464
rect 17184 46452 17190 46504
rect 17310 46492 17316 46504
rect 17271 46464 17316 46492
rect 17310 46452 17316 46464
rect 17368 46452 17374 46504
rect 17405 46495 17463 46501
rect 17405 46461 17417 46495
rect 17451 46461 17463 46495
rect 17405 46455 17463 46461
rect 17497 46495 17555 46501
rect 17497 46461 17509 46495
rect 17543 46461 17555 46495
rect 17678 46492 17684 46504
rect 17639 46464 17684 46492
rect 17497 46455 17555 46461
rect 9766 46424 9772 46436
rect 9324 46396 9772 46424
rect 7616 46384 7622 46396
rect 9766 46384 9772 46396
rect 9824 46384 9830 46436
rect 9861 46427 9919 46433
rect 9861 46393 9873 46427
rect 9907 46424 9919 46427
rect 10566 46427 10624 46433
rect 10566 46424 10578 46427
rect 9907 46396 10578 46424
rect 9907 46393 9919 46396
rect 9861 46387 9919 46393
rect 10566 46393 10578 46396
rect 10612 46393 10624 46427
rect 10566 46387 10624 46393
rect 12428 46427 12486 46433
rect 12428 46393 12440 46427
rect 12474 46424 12486 46427
rect 14090 46424 14096 46436
rect 12474 46396 14096 46424
rect 12474 46393 12486 46396
rect 12428 46387 12486 46393
rect 14090 46384 14096 46396
rect 14148 46384 14154 46436
rect 14642 46433 14648 46436
rect 14636 46387 14648 46433
rect 14700 46424 14706 46436
rect 14700 46396 14736 46424
rect 14642 46384 14648 46387
rect 14700 46384 14706 46396
rect 11698 46356 11704 46368
rect 11659 46328 11704 46356
rect 11698 46316 11704 46328
rect 11756 46316 11762 46368
rect 12618 46316 12624 46368
rect 12676 46356 12682 46368
rect 13722 46356 13728 46368
rect 12676 46328 13728 46356
rect 12676 46316 12682 46328
rect 13722 46316 13728 46328
rect 13780 46316 13786 46368
rect 15102 46316 15108 46368
rect 15160 46356 15166 46368
rect 15749 46359 15807 46365
rect 15749 46356 15761 46359
rect 15160 46328 15761 46356
rect 15160 46316 15166 46328
rect 15749 46325 15761 46328
rect 15795 46325 15807 46359
rect 16298 46356 16304 46368
rect 16259 46328 16304 46356
rect 15749 46319 15807 46325
rect 16298 46316 16304 46328
rect 16356 46316 16362 46368
rect 17420 46356 17448 46455
rect 17512 46424 17540 46455
rect 17678 46452 17684 46464
rect 17736 46452 17742 46504
rect 18322 46452 18328 46504
rect 18380 46492 18386 46504
rect 24210 46492 24216 46504
rect 18380 46464 24216 46492
rect 18380 46452 18386 46464
rect 24210 46452 24216 46464
rect 24268 46452 24274 46504
rect 24397 46495 24455 46501
rect 24397 46461 24409 46495
rect 24443 46461 24455 46495
rect 24397 46455 24455 46461
rect 17586 46424 17592 46436
rect 17512 46396 17592 46424
rect 17586 46384 17592 46396
rect 17644 46384 17650 46436
rect 19610 46384 19616 46436
rect 19668 46424 19674 46436
rect 20070 46424 20076 46436
rect 19668 46396 20076 46424
rect 19668 46384 19674 46396
rect 20070 46384 20076 46396
rect 20128 46424 20134 46436
rect 20257 46427 20315 46433
rect 20257 46424 20269 46427
rect 20128 46396 20269 46424
rect 20128 46384 20134 46396
rect 20257 46393 20269 46396
rect 20303 46393 20315 46427
rect 20257 46387 20315 46393
rect 20806 46384 20812 46436
rect 20864 46424 20870 46436
rect 22710 46427 22768 46433
rect 22710 46424 22722 46427
rect 20864 46396 22722 46424
rect 20864 46384 20870 46396
rect 22710 46393 22722 46396
rect 22756 46393 22768 46427
rect 22710 46387 22768 46393
rect 23106 46384 23112 46436
rect 23164 46424 23170 46436
rect 24412 46424 24440 46455
rect 24486 46452 24492 46504
rect 24544 46494 24550 46504
rect 24780 46501 24808 46600
rect 24581 46495 24639 46501
rect 24581 46494 24593 46495
rect 24544 46466 24593 46494
rect 24544 46452 24550 46466
rect 24581 46461 24593 46466
rect 24627 46461 24639 46495
rect 24581 46455 24639 46461
rect 24765 46495 24823 46501
rect 24765 46461 24777 46495
rect 24811 46461 24823 46495
rect 24949 46495 25007 46501
rect 24949 46492 24961 46495
rect 24765 46455 24823 46461
rect 24872 46464 24961 46492
rect 23164 46396 24440 46424
rect 23164 46384 23170 46396
rect 17494 46356 17500 46368
rect 17420 46328 17500 46356
rect 17494 46316 17500 46328
rect 17552 46316 17558 46368
rect 19797 46359 19855 46365
rect 19797 46325 19809 46359
rect 19843 46356 19855 46359
rect 19978 46356 19984 46368
rect 19843 46328 19984 46356
rect 19843 46325 19855 46328
rect 19797 46319 19855 46325
rect 19978 46316 19984 46328
rect 20036 46316 20042 46368
rect 20714 46316 20720 46368
rect 20772 46356 20778 46368
rect 21545 46359 21603 46365
rect 21545 46356 21557 46359
rect 20772 46328 21557 46356
rect 20772 46316 20778 46328
rect 21545 46325 21557 46328
rect 21591 46356 21603 46359
rect 21910 46356 21916 46368
rect 21591 46328 21916 46356
rect 21591 46325 21603 46328
rect 21545 46319 21603 46325
rect 21910 46316 21916 46328
rect 21968 46316 21974 46368
rect 22002 46316 22008 46368
rect 22060 46356 22066 46368
rect 23658 46356 23664 46368
rect 22060 46328 23664 46356
rect 22060 46316 22066 46328
rect 23658 46316 23664 46328
rect 23716 46356 23722 46368
rect 23845 46359 23903 46365
rect 23845 46356 23857 46359
rect 23716 46328 23857 46356
rect 23716 46316 23722 46328
rect 23845 46325 23857 46328
rect 23891 46325 23903 46359
rect 23845 46319 23903 46325
rect 24302 46316 24308 46368
rect 24360 46356 24366 46368
rect 24872 46356 24900 46464
rect 24949 46461 24961 46464
rect 24995 46492 25007 46495
rect 25593 46495 25651 46501
rect 25593 46492 25605 46495
rect 24995 46464 25605 46492
rect 24995 46461 25007 46464
rect 24949 46455 25007 46461
rect 25593 46461 25605 46464
rect 25639 46461 25651 46495
rect 25593 46455 25651 46461
rect 25130 46356 25136 46368
rect 24360 46328 24900 46356
rect 25091 46328 25136 46356
rect 24360 46316 24366 46328
rect 25130 46316 25136 46328
rect 25188 46316 25194 46368
rect 25682 46356 25688 46368
rect 25643 46328 25688 46356
rect 25682 46316 25688 46328
rect 25740 46316 25746 46368
rect 1104 46266 32016 46288
rect 1104 46214 11253 46266
rect 11305 46214 11317 46266
rect 11369 46214 11381 46266
rect 11433 46214 11445 46266
rect 11497 46214 11509 46266
rect 11561 46214 21557 46266
rect 21609 46214 21621 46266
rect 21673 46214 21685 46266
rect 21737 46214 21749 46266
rect 21801 46214 21813 46266
rect 21865 46214 32016 46266
rect 1104 46192 32016 46214
rect 9398 46152 9404 46164
rect 9324 46124 9404 46152
rect 7742 46084 7748 46096
rect 6380 46056 7748 46084
rect 1394 46025 1400 46028
rect 1385 46019 1400 46025
rect 1385 46016 1397 46019
rect 1044 45988 1397 46016
rect 0 45948 800 45962
rect 1044 45948 1072 45988
rect 1385 45985 1397 45988
rect 1385 45979 1400 45985
rect 1394 45976 1400 45979
rect 1452 45976 1458 46028
rect 6380 46025 6408 46056
rect 7742 46044 7748 46056
rect 7800 46044 7806 46096
rect 6365 46019 6423 46025
rect 6365 45985 6377 46019
rect 6411 45985 6423 46019
rect 6365 45979 6423 45985
rect 6632 46019 6690 46025
rect 6632 45985 6644 46019
rect 6678 46016 6690 46019
rect 7190 46016 7196 46028
rect 6678 45988 7196 46016
rect 6678 45985 6690 45988
rect 6632 45979 6690 45985
rect 7190 45976 7196 45988
rect 7248 45976 7254 46028
rect 8389 46019 8447 46025
rect 8389 45985 8401 46019
rect 8435 45985 8447 46019
rect 9030 46016 9036 46028
rect 8943 45988 9036 46016
rect 8389 45979 8447 45985
rect 0 45920 1072 45948
rect 0 45906 800 45920
rect 7466 45840 7472 45892
rect 7524 45880 7530 45892
rect 7745 45883 7803 45889
rect 7745 45880 7757 45883
rect 7524 45852 7757 45880
rect 7524 45840 7530 45852
rect 7745 45849 7757 45852
rect 7791 45880 7803 45883
rect 8404 45880 8432 45979
rect 9030 45976 9036 45988
rect 9088 45976 9094 46028
rect 9214 46016 9220 46028
rect 9175 45988 9220 46016
rect 9214 45976 9220 45988
rect 9272 45976 9278 46028
rect 9048 45948 9076 45976
rect 9324 45957 9352 46124
rect 9398 46112 9404 46124
rect 9456 46112 9462 46164
rect 9769 46155 9827 46161
rect 9769 46121 9781 46155
rect 9815 46152 9827 46155
rect 9858 46152 9864 46164
rect 9815 46124 9864 46152
rect 9815 46121 9827 46124
rect 9769 46115 9827 46121
rect 9858 46112 9864 46124
rect 9916 46112 9922 46164
rect 10962 46152 10968 46164
rect 10923 46124 10968 46152
rect 10962 46112 10968 46124
rect 11020 46112 11026 46164
rect 13354 46152 13360 46164
rect 13315 46124 13360 46152
rect 13354 46112 13360 46124
rect 13412 46112 13418 46164
rect 14553 46155 14611 46161
rect 14553 46121 14565 46155
rect 14599 46152 14611 46155
rect 14642 46152 14648 46164
rect 14599 46124 14648 46152
rect 14599 46121 14611 46124
rect 14553 46115 14611 46121
rect 14642 46112 14648 46124
rect 14700 46112 14706 46164
rect 15746 46152 15752 46164
rect 15707 46124 15752 46152
rect 15746 46112 15752 46124
rect 15804 46112 15810 46164
rect 17402 46152 17408 46164
rect 17363 46124 17408 46152
rect 17402 46112 17408 46124
rect 17460 46112 17466 46164
rect 18782 46152 18788 46164
rect 18743 46124 18788 46152
rect 18782 46112 18788 46124
rect 18840 46112 18846 46164
rect 20717 46155 20775 46161
rect 20717 46121 20729 46155
rect 20763 46152 20775 46155
rect 20806 46152 20812 46164
rect 20763 46124 20812 46152
rect 20763 46121 20775 46124
rect 20717 46115 20775 46121
rect 20806 46112 20812 46124
rect 20864 46112 20870 46164
rect 22002 46152 22008 46164
rect 21928 46124 22008 46152
rect 9674 46044 9680 46096
rect 9732 46084 9738 46096
rect 15378 46084 15384 46096
rect 9732 46056 11560 46084
rect 9732 46044 9738 46056
rect 9401 46019 9459 46025
rect 9401 45985 9413 46019
rect 9447 46016 9459 46019
rect 9490 46016 9496 46028
rect 9447 45988 9496 46016
rect 9447 45985 9459 45988
rect 9401 45979 9459 45985
rect 9490 45976 9496 45988
rect 9548 45976 9554 46028
rect 9585 46019 9643 46025
rect 9585 45985 9597 46019
rect 9631 46016 9643 46019
rect 9766 46016 9772 46028
rect 9631 45988 9772 46016
rect 9631 45985 9643 45988
rect 9585 45979 9643 45985
rect 9766 45976 9772 45988
rect 9824 45976 9830 46028
rect 10226 46016 10232 46028
rect 10187 45988 10232 46016
rect 10226 45976 10232 45988
rect 10284 45976 10290 46028
rect 10428 46025 10456 46056
rect 10413 46019 10471 46025
rect 10413 45985 10425 46019
rect 10459 45985 10471 46019
rect 10778 46016 10784 46028
rect 10739 45988 10784 46016
rect 10413 45979 10471 45985
rect 10778 45976 10784 45988
rect 10836 45976 10842 46028
rect 11532 46016 11560 46056
rect 13188 46056 15384 46084
rect 11698 46025 11704 46028
rect 11677 46019 11704 46025
rect 11677 46016 11689 46019
rect 11532 45988 11689 46016
rect 11677 45985 11689 45988
rect 11677 45979 11704 45985
rect 11698 45976 11704 45979
rect 11756 45976 11762 46028
rect 12618 46016 12624 46028
rect 12579 45988 12624 46016
rect 12618 45976 12624 45988
rect 12676 45976 12682 46028
rect 12802 46016 12808 46028
rect 12763 45988 12808 46016
rect 12802 45976 12808 45988
rect 12860 45976 12866 46028
rect 13188 46025 13216 46056
rect 13173 46019 13231 46025
rect 13173 45985 13185 46019
rect 13219 45985 13231 46019
rect 13173 45979 13231 45985
rect 13722 45976 13728 46028
rect 13780 46016 13786 46028
rect 14016 46025 14044 46056
rect 15378 46044 15384 46056
rect 15436 46044 15442 46096
rect 16114 46044 16120 46096
rect 16172 46084 16178 46096
rect 17494 46084 17500 46096
rect 16172 46056 16896 46084
rect 16172 46044 16178 46056
rect 13817 46019 13875 46025
rect 13817 46016 13829 46019
rect 13780 45988 13829 46016
rect 13780 45976 13786 45988
rect 13817 45985 13829 45988
rect 13863 45985 13875 46019
rect 13817 45979 13875 45985
rect 14001 46019 14059 46025
rect 14001 45985 14013 46019
rect 14047 45985 14059 46019
rect 14001 45979 14059 45985
rect 14369 46019 14427 46025
rect 14369 45985 14381 46019
rect 14415 45985 14427 46019
rect 14369 45979 14427 45985
rect 9309 45951 9367 45957
rect 9048 45920 9168 45948
rect 7791 45852 8432 45880
rect 7791 45849 7803 45852
rect 7745 45843 7803 45849
rect 1581 45815 1639 45821
rect 1581 45781 1593 45815
rect 1627 45812 1639 45815
rect 4982 45812 4988 45824
rect 1627 45784 4988 45812
rect 1627 45781 1639 45784
rect 1581 45775 1639 45781
rect 4982 45772 4988 45784
rect 5040 45772 5046 45824
rect 8386 45772 8392 45824
rect 8444 45812 8450 45824
rect 8481 45815 8539 45821
rect 8481 45812 8493 45815
rect 8444 45784 8493 45812
rect 8444 45772 8450 45784
rect 8481 45781 8493 45784
rect 8527 45781 8539 45815
rect 9140 45812 9168 45920
rect 9309 45917 9321 45951
rect 9355 45948 9367 45951
rect 10502 45948 10508 45960
rect 9355 45920 10508 45948
rect 9355 45917 9367 45920
rect 9309 45911 9367 45917
rect 10502 45908 10508 45920
rect 10560 45908 10566 45960
rect 10594 45908 10600 45960
rect 10652 45948 10658 45960
rect 12894 45948 12900 45960
rect 10652 45920 10697 45948
rect 12855 45920 12900 45948
rect 10652 45908 10658 45920
rect 12894 45908 12900 45920
rect 12952 45908 12958 45960
rect 12986 45908 12992 45960
rect 13044 45948 13050 45960
rect 14093 45951 14151 45957
rect 14093 45948 14105 45951
rect 13044 45920 13089 45948
rect 13832 45920 14105 45948
rect 13044 45908 13050 45920
rect 9766 45840 9772 45892
rect 9824 45880 9830 45892
rect 10870 45880 10876 45892
rect 9824 45852 10876 45880
rect 9824 45840 9830 45852
rect 10870 45840 10876 45852
rect 10928 45840 10934 45892
rect 10226 45812 10232 45824
rect 9140 45784 10232 45812
rect 8481 45775 8539 45781
rect 10226 45772 10232 45784
rect 10284 45772 10290 45824
rect 10962 45772 10968 45824
rect 11020 45812 11026 45824
rect 11609 45815 11667 45821
rect 11609 45812 11621 45815
rect 11020 45784 11621 45812
rect 11020 45772 11026 45784
rect 11609 45781 11621 45784
rect 11655 45781 11667 45815
rect 13004 45812 13032 45908
rect 13078 45840 13084 45892
rect 13136 45880 13142 45892
rect 13722 45880 13728 45892
rect 13136 45852 13728 45880
rect 13136 45840 13142 45852
rect 13722 45840 13728 45852
rect 13780 45880 13786 45892
rect 13832 45880 13860 45920
rect 14093 45917 14105 45920
rect 14139 45917 14151 45951
rect 14093 45911 14151 45917
rect 14182 45908 14188 45960
rect 14240 45948 14246 45960
rect 14384 45948 14412 45979
rect 14826 45976 14832 46028
rect 14884 46016 14890 46028
rect 15013 46019 15071 46025
rect 15013 46016 15025 46019
rect 14884 45988 15025 46016
rect 14884 45976 14890 45988
rect 15013 45985 15025 45988
rect 15059 45985 15071 46019
rect 15013 45979 15071 45985
rect 15102 45976 15108 46028
rect 15160 46016 15166 46028
rect 15197 46019 15255 46025
rect 15197 46016 15209 46019
rect 15160 45988 15209 46016
rect 15160 45976 15166 45988
rect 15197 45985 15209 45988
rect 15243 45985 15255 46019
rect 15197 45979 15255 45985
rect 15565 46019 15623 46025
rect 15565 45985 15577 46019
rect 15611 46016 15623 46019
rect 16132 46016 16160 46044
rect 16666 46016 16672 46028
rect 15611 45988 16160 46016
rect 16627 45988 16672 46016
rect 15611 45985 15623 45988
rect 15565 45979 15623 45985
rect 16666 45976 16672 45988
rect 16724 45976 16730 46028
rect 16868 46025 16896 46056
rect 16960 46056 17500 46084
rect 16960 46025 16988 46056
rect 17494 46044 17500 46056
rect 17552 46044 17558 46096
rect 21928 46084 21956 46124
rect 22002 46112 22008 46124
rect 22060 46112 22066 46164
rect 22278 46084 22284 46096
rect 19444 46056 20300 46084
rect 16853 46019 16911 46025
rect 16853 45985 16865 46019
rect 16899 45985 16911 46019
rect 16853 45979 16911 45985
rect 16945 46019 17003 46025
rect 16945 45985 16957 46019
rect 16991 45985 17003 46019
rect 16945 45979 17003 45985
rect 17221 46019 17279 46025
rect 17221 45985 17233 46019
rect 17267 46016 17279 46019
rect 17310 46016 17316 46028
rect 17267 45988 17316 46016
rect 17267 45985 17279 45988
rect 17221 45979 17279 45985
rect 17310 45976 17316 45988
rect 17368 46016 17374 46028
rect 17865 46019 17923 46025
rect 17865 46016 17877 46019
rect 17368 45988 17877 46016
rect 17368 45976 17374 45988
rect 17865 45985 17877 45988
rect 17911 45985 17923 46019
rect 18966 46016 18972 46028
rect 18927 45988 18972 46016
rect 17865 45979 17923 45985
rect 18966 45976 18972 45988
rect 19024 45976 19030 46028
rect 19334 46016 19340 46028
rect 19295 45988 19340 46016
rect 19334 45976 19340 45988
rect 19392 45976 19398 46028
rect 15120 45948 15148 45976
rect 15286 45948 15292 45960
rect 14240 45920 14285 45948
rect 14384 45920 15148 45948
rect 15247 45920 15292 45948
rect 14240 45908 14246 45920
rect 13780 45852 13860 45880
rect 13780 45840 13786 45852
rect 13906 45840 13912 45892
rect 13964 45880 13970 45892
rect 14384 45880 14412 45920
rect 15286 45908 15292 45920
rect 15344 45908 15350 45960
rect 15381 45951 15439 45957
rect 15381 45917 15393 45951
rect 15427 45948 15439 45951
rect 17037 45951 17095 45957
rect 17037 45948 17049 45951
rect 15427 45920 17049 45948
rect 15427 45917 15439 45920
rect 15381 45911 15439 45917
rect 17037 45917 17049 45920
rect 17083 45948 17095 45951
rect 17586 45948 17592 45960
rect 17083 45920 17592 45948
rect 17083 45917 17095 45920
rect 17037 45911 17095 45917
rect 17586 45908 17592 45920
rect 17644 45908 17650 45960
rect 19153 45951 19211 45957
rect 19153 45917 19165 45951
rect 19199 45917 19211 45951
rect 19153 45911 19211 45917
rect 19245 45951 19303 45957
rect 19245 45917 19257 45951
rect 19291 45948 19303 45951
rect 19444 45948 19472 46056
rect 19521 46019 19579 46025
rect 19521 45985 19533 46019
rect 19567 46016 19579 46019
rect 19981 46019 20039 46025
rect 19981 46016 19993 46019
rect 19567 45988 19993 46016
rect 19567 45985 19579 45988
rect 19521 45979 19579 45985
rect 19981 45985 19993 45988
rect 20027 45985 20039 46019
rect 20162 46016 20168 46028
rect 20123 45988 20168 46016
rect 19981 45979 20039 45985
rect 19291 45920 19472 45948
rect 19996 45948 20024 45979
rect 20162 45976 20168 45988
rect 20220 45976 20226 46028
rect 20272 46025 20300 46056
rect 20548 46056 21956 46084
rect 22020 46056 22284 46084
rect 20548 46025 20576 46056
rect 20257 46019 20315 46025
rect 20257 45985 20269 46019
rect 20303 46016 20315 46019
rect 20533 46019 20591 46025
rect 20303 45988 20484 46016
rect 20303 45985 20315 45988
rect 20257 45979 20315 45985
rect 20346 45948 20352 45960
rect 19996 45920 20116 45948
rect 20307 45920 20352 45948
rect 19291 45917 19303 45920
rect 19245 45911 19303 45917
rect 13964 45852 14412 45880
rect 13964 45840 13970 45852
rect 14182 45812 14188 45824
rect 13004 45784 14188 45812
rect 11609 45775 11667 45781
rect 14182 45772 14188 45784
rect 14240 45772 14246 45824
rect 17957 45815 18015 45821
rect 17957 45781 17969 45815
rect 18003 45812 18015 45815
rect 18046 45812 18052 45824
rect 18003 45784 18052 45812
rect 18003 45781 18015 45784
rect 17957 45775 18015 45781
rect 18046 45772 18052 45784
rect 18104 45772 18110 45824
rect 19168 45812 19196 45911
rect 20088 45880 20116 45920
rect 20346 45908 20352 45920
rect 20404 45908 20410 45960
rect 20456 45948 20484 45988
rect 20533 45985 20545 46019
rect 20579 45985 20591 46019
rect 20533 45979 20591 45985
rect 20806 45976 20812 46028
rect 20864 46016 20870 46028
rect 22020 46025 22048 46056
rect 22278 46044 22284 46056
rect 22336 46044 22342 46096
rect 23192 46087 23250 46093
rect 23192 46053 23204 46087
rect 23238 46084 23250 46087
rect 25130 46084 25136 46096
rect 23238 46056 25136 46084
rect 23238 46053 23250 46056
rect 23192 46047 23250 46053
rect 25130 46044 25136 46056
rect 25188 46044 25194 46096
rect 21177 46019 21235 46025
rect 21177 46016 21189 46019
rect 20864 45988 21189 46016
rect 20864 45976 20870 45988
rect 21177 45985 21189 45988
rect 21223 45985 21235 46019
rect 21177 45979 21235 45985
rect 22005 46019 22063 46025
rect 22005 45985 22017 46019
rect 22051 45985 22063 46019
rect 22005 45979 22063 45985
rect 22094 45976 22100 46028
rect 22152 46016 22158 46028
rect 22370 46016 22376 46028
rect 22152 45988 22197 46016
rect 22331 45988 22376 46016
rect 22152 45976 22158 45988
rect 22370 45976 22376 45988
rect 22428 45976 22434 46028
rect 22833 46019 22891 46025
rect 22833 45985 22845 46019
rect 22879 46016 22891 46019
rect 24026 46016 24032 46028
rect 22879 45988 24032 46016
rect 22879 45985 22891 45988
rect 22833 45979 22891 45985
rect 24026 45976 24032 45988
rect 24084 45976 24090 46028
rect 24118 45976 24124 46028
rect 24176 46016 24182 46028
rect 25878 46019 25936 46025
rect 25878 46016 25890 46019
rect 24176 45988 25890 46016
rect 24176 45976 24182 45988
rect 25878 45985 25890 45988
rect 25924 45985 25936 46019
rect 30650 46016 30656 46028
rect 30563 45988 30656 46016
rect 25878 45979 25936 45985
rect 30650 45976 30656 45988
rect 30708 46016 30714 46028
rect 31113 46019 31171 46025
rect 31113 46016 31125 46019
rect 30708 45988 31125 46016
rect 30708 45976 30714 45988
rect 31113 45985 31125 45988
rect 31159 46016 31171 46019
rect 31570 46016 31576 46028
rect 31159 45988 31576 46016
rect 31159 45985 31171 45988
rect 31113 45979 31171 45985
rect 31570 45976 31576 45988
rect 31628 45976 31634 46028
rect 21266 45948 21272 45960
rect 20456 45920 21272 45948
rect 21266 45908 21272 45920
rect 21324 45948 21330 45960
rect 21542 45948 21548 45960
rect 21324 45920 21548 45948
rect 21324 45908 21330 45920
rect 21542 45908 21548 45920
rect 21600 45908 21606 45960
rect 21910 45908 21916 45960
rect 21968 45948 21974 45960
rect 22925 45951 22983 45957
rect 22925 45948 22937 45951
rect 21968 45920 22937 45948
rect 21968 45908 21974 45920
rect 22925 45917 22937 45920
rect 22971 45917 22983 45951
rect 26142 45948 26148 45960
rect 26103 45920 26148 45948
rect 22925 45911 22983 45917
rect 26142 45908 26148 45920
rect 26200 45908 26206 45960
rect 32320 45948 33120 45962
rect 31726 45920 33120 45948
rect 21450 45880 21456 45892
rect 20088 45852 21456 45880
rect 21450 45840 21456 45852
rect 21508 45840 21514 45892
rect 22281 45883 22339 45889
rect 22281 45849 22293 45883
rect 22327 45880 22339 45883
rect 22833 45883 22891 45889
rect 22833 45880 22845 45883
rect 22327 45852 22845 45880
rect 22327 45849 22339 45852
rect 22281 45843 22339 45849
rect 22833 45849 22845 45852
rect 22879 45849 22891 45883
rect 22833 45843 22891 45849
rect 24210 45840 24216 45892
rect 24268 45880 24274 45892
rect 31297 45883 31355 45889
rect 24268 45852 25268 45880
rect 24268 45840 24274 45852
rect 20346 45812 20352 45824
rect 19168 45784 20352 45812
rect 20346 45772 20352 45784
rect 20404 45812 20410 45824
rect 20898 45812 20904 45824
rect 20404 45784 20904 45812
rect 20404 45772 20410 45784
rect 20898 45772 20904 45784
rect 20956 45772 20962 45824
rect 21082 45772 21088 45824
rect 21140 45812 21146 45824
rect 21634 45812 21640 45824
rect 21140 45784 21640 45812
rect 21140 45772 21146 45784
rect 21634 45772 21640 45784
rect 21692 45772 21698 45824
rect 21821 45815 21879 45821
rect 21821 45781 21833 45815
rect 21867 45812 21879 45815
rect 21910 45812 21916 45824
rect 21867 45784 21916 45812
rect 21867 45781 21879 45784
rect 21821 45775 21879 45781
rect 21910 45772 21916 45784
rect 21968 45772 21974 45824
rect 24302 45812 24308 45824
rect 24263 45784 24308 45812
rect 24302 45772 24308 45784
rect 24360 45772 24366 45824
rect 24394 45772 24400 45824
rect 24452 45812 24458 45824
rect 24765 45815 24823 45821
rect 24765 45812 24777 45815
rect 24452 45784 24777 45812
rect 24452 45772 24458 45784
rect 24765 45781 24777 45784
rect 24811 45781 24823 45815
rect 25240 45812 25268 45852
rect 31297 45849 31309 45883
rect 31343 45880 31355 45883
rect 31726 45880 31754 45920
rect 32320 45906 33120 45920
rect 31343 45852 31754 45880
rect 31343 45849 31355 45852
rect 31297 45843 31355 45849
rect 26234 45812 26240 45824
rect 25240 45784 26240 45812
rect 24765 45775 24823 45781
rect 26234 45772 26240 45784
rect 26292 45772 26298 45824
rect 1104 45722 32016 45744
rect 1104 45670 6102 45722
rect 6154 45670 6166 45722
rect 6218 45670 6230 45722
rect 6282 45670 6294 45722
rect 6346 45670 6358 45722
rect 6410 45670 16405 45722
rect 16457 45670 16469 45722
rect 16521 45670 16533 45722
rect 16585 45670 16597 45722
rect 16649 45670 16661 45722
rect 16713 45670 26709 45722
rect 26761 45670 26773 45722
rect 26825 45670 26837 45722
rect 26889 45670 26901 45722
rect 26953 45670 26965 45722
rect 27017 45670 32016 45722
rect 1104 45648 32016 45670
rect 1394 45608 1400 45620
rect 1355 45580 1400 45608
rect 1394 45568 1400 45580
rect 1452 45568 1458 45620
rect 9401 45611 9459 45617
rect 9401 45577 9413 45611
rect 9447 45608 9459 45611
rect 9490 45608 9496 45620
rect 9447 45580 9496 45608
rect 9447 45577 9459 45580
rect 9401 45571 9459 45577
rect 9490 45568 9496 45580
rect 9548 45608 9554 45620
rect 10594 45608 10600 45620
rect 9548 45580 10600 45608
rect 9548 45568 9554 45580
rect 10594 45568 10600 45580
rect 10652 45568 10658 45620
rect 13722 45568 13728 45620
rect 13780 45608 13786 45620
rect 15286 45608 15292 45620
rect 13780 45580 15292 45608
rect 13780 45568 13786 45580
rect 8018 45540 8024 45552
rect 7979 45512 8024 45540
rect 8018 45500 8024 45512
rect 8076 45500 8082 45552
rect 9858 45500 9864 45552
rect 9916 45540 9922 45552
rect 11606 45540 11612 45552
rect 9916 45512 11612 45540
rect 9916 45500 9922 45512
rect 11606 45500 11612 45512
rect 11664 45540 11670 45552
rect 14182 45540 14188 45552
rect 11664 45512 14188 45540
rect 11664 45500 11670 45512
rect 14182 45500 14188 45512
rect 14240 45500 14246 45552
rect 14274 45500 14280 45552
rect 14332 45500 14338 45552
rect 7558 45472 7564 45484
rect 7519 45444 7564 45472
rect 7558 45432 7564 45444
rect 7616 45432 7622 45484
rect 12805 45475 12863 45481
rect 12805 45441 12817 45475
rect 12851 45472 12863 45475
rect 12894 45472 12900 45484
rect 12851 45444 12900 45472
rect 12851 45441 12863 45444
rect 12805 45435 12863 45441
rect 12894 45432 12900 45444
rect 12952 45432 12958 45484
rect 14090 45472 14096 45484
rect 14051 45444 14096 45472
rect 14090 45432 14096 45444
rect 14148 45432 14154 45484
rect 14292 45472 14320 45500
rect 14568 45481 14596 45580
rect 15286 45568 15292 45580
rect 15344 45568 15350 45620
rect 19610 45568 19616 45620
rect 19668 45608 19674 45620
rect 26142 45608 26148 45620
rect 19668 45580 24348 45608
rect 19668 45568 19674 45580
rect 16206 45500 16212 45552
rect 16264 45540 16270 45552
rect 16393 45543 16451 45549
rect 16393 45540 16405 45543
rect 16264 45512 16405 45540
rect 16264 45500 16270 45512
rect 16393 45509 16405 45512
rect 16439 45509 16451 45543
rect 16393 45503 16451 45509
rect 20990 45500 20996 45552
rect 21048 45540 21054 45552
rect 21085 45543 21143 45549
rect 21085 45540 21097 45543
rect 21048 45512 21097 45540
rect 21048 45500 21054 45512
rect 21085 45509 21097 45512
rect 21131 45509 21143 45543
rect 21085 45503 21143 45509
rect 21450 45500 21456 45552
rect 21508 45500 21514 45552
rect 22278 45500 22284 45552
rect 22336 45540 22342 45552
rect 22373 45543 22431 45549
rect 22373 45540 22385 45543
rect 22336 45512 22385 45540
rect 22336 45500 22342 45512
rect 22373 45509 22385 45512
rect 22419 45509 22431 45543
rect 22373 45503 22431 45509
rect 23474 45500 23480 45552
rect 23532 45500 23538 45552
rect 14461 45475 14519 45481
rect 14461 45472 14473 45475
rect 14292 45444 14473 45472
rect 14461 45441 14473 45444
rect 14507 45441 14519 45475
rect 14461 45435 14519 45441
rect 14553 45475 14611 45481
rect 14553 45441 14565 45475
rect 14599 45441 14611 45475
rect 14553 45435 14611 45441
rect 15746 45432 15752 45484
rect 15804 45472 15810 45484
rect 15804 45444 16252 45472
rect 15804 45432 15810 45444
rect 6825 45407 6883 45413
rect 6825 45373 6837 45407
rect 6871 45404 6883 45407
rect 6914 45404 6920 45416
rect 6871 45376 6920 45404
rect 6871 45373 6883 45376
rect 6825 45367 6883 45373
rect 6914 45364 6920 45376
rect 6972 45364 6978 45416
rect 7282 45404 7288 45416
rect 7243 45376 7288 45404
rect 7282 45364 7288 45376
rect 7340 45364 7346 45416
rect 7466 45404 7472 45416
rect 7524 45413 7530 45416
rect 7431 45376 7472 45404
rect 7466 45364 7472 45376
rect 7524 45367 7531 45413
rect 7653 45407 7711 45413
rect 7653 45373 7665 45407
rect 7699 45373 7711 45407
rect 7834 45404 7840 45416
rect 7795 45376 7840 45404
rect 7653 45367 7711 45373
rect 7524 45364 7530 45367
rect 7374 45296 7380 45348
rect 7432 45336 7438 45348
rect 7668 45336 7696 45367
rect 7834 45364 7840 45376
rect 7892 45364 7898 45416
rect 9214 45364 9220 45416
rect 9272 45404 9278 45416
rect 10045 45407 10103 45413
rect 10045 45404 10057 45407
rect 9272 45376 10057 45404
rect 9272 45364 9278 45376
rect 10045 45373 10057 45376
rect 10091 45373 10103 45407
rect 10870 45404 10876 45416
rect 10831 45376 10876 45404
rect 10045 45367 10103 45373
rect 10870 45364 10876 45376
rect 10928 45364 10934 45416
rect 11425 45407 11483 45413
rect 11425 45373 11437 45407
rect 11471 45404 11483 45407
rect 11974 45404 11980 45416
rect 11471 45376 11980 45404
rect 11471 45373 11483 45376
rect 11425 45367 11483 45373
rect 11974 45364 11980 45376
rect 12032 45364 12038 45416
rect 12069 45407 12127 45413
rect 12069 45373 12081 45407
rect 12115 45404 12127 45407
rect 12526 45404 12532 45416
rect 12115 45376 12434 45404
rect 12487 45376 12532 45404
rect 12115 45373 12127 45376
rect 12069 45367 12127 45373
rect 9490 45336 9496 45348
rect 7432 45308 7696 45336
rect 9451 45308 9496 45336
rect 7432 45296 7438 45308
rect 9490 45296 9496 45308
rect 9548 45296 9554 45348
rect 12406 45336 12434 45376
rect 12526 45364 12532 45376
rect 12584 45364 12590 45416
rect 13814 45364 13820 45416
rect 13872 45404 13878 45416
rect 14277 45407 14335 45413
rect 14277 45404 14289 45407
rect 13872 45376 14289 45404
rect 13872 45364 13878 45376
rect 14277 45373 14289 45376
rect 14323 45373 14335 45407
rect 14277 45367 14335 45373
rect 13906 45336 13912 45348
rect 12406 45308 13912 45336
rect 13906 45296 13912 45308
rect 13964 45296 13970 45348
rect 14292 45336 14320 45367
rect 14642 45364 14648 45416
rect 14700 45404 14706 45416
rect 14700 45376 14745 45404
rect 14700 45364 14706 45376
rect 14826 45364 14832 45416
rect 14884 45404 14890 45416
rect 16224 45413 16252 45444
rect 20898 45432 20904 45484
rect 20956 45472 20962 45484
rect 21468 45472 21496 45500
rect 23385 45475 23443 45481
rect 20956 45444 21404 45472
rect 21468 45444 21864 45472
rect 20956 45432 20962 45444
rect 15289 45407 15347 45413
rect 14884 45376 14929 45404
rect 14884 45364 14890 45376
rect 15289 45373 15301 45407
rect 15335 45373 15347 45407
rect 15289 45367 15347 45373
rect 16117 45407 16175 45413
rect 16117 45373 16129 45407
rect 16163 45373 16175 45407
rect 16117 45367 16175 45373
rect 16209 45407 16267 45413
rect 16209 45373 16221 45407
rect 16255 45373 16267 45407
rect 16209 45367 16267 45373
rect 16485 45407 16543 45413
rect 16485 45373 16497 45407
rect 16531 45404 16543 45407
rect 17313 45407 17371 45413
rect 16531 45376 17264 45404
rect 16531 45373 16543 45376
rect 16485 45367 16543 45373
rect 15304 45336 15332 45367
rect 14292 45308 15332 45336
rect 16132 45336 16160 45367
rect 16666 45336 16672 45348
rect 16132 45308 16672 45336
rect 16666 45296 16672 45308
rect 16724 45296 16730 45348
rect 6733 45271 6791 45277
rect 6733 45237 6745 45271
rect 6779 45268 6791 45271
rect 8018 45268 8024 45280
rect 6779 45240 8024 45268
rect 6779 45237 6791 45240
rect 6733 45231 6791 45237
rect 8018 45228 8024 45240
rect 8076 45228 8082 45280
rect 9766 45228 9772 45280
rect 9824 45268 9830 45280
rect 10137 45271 10195 45277
rect 10137 45268 10149 45271
rect 9824 45240 10149 45268
rect 9824 45228 9830 45240
rect 10137 45237 10149 45240
rect 10183 45237 10195 45271
rect 10778 45268 10784 45280
rect 10739 45240 10784 45268
rect 10137 45231 10195 45237
rect 10778 45228 10784 45240
rect 10836 45228 10842 45280
rect 11977 45271 12035 45277
rect 11977 45237 11989 45271
rect 12023 45268 12035 45271
rect 15102 45268 15108 45280
rect 12023 45240 15108 45268
rect 12023 45237 12035 45240
rect 11977 45231 12035 45237
rect 15102 45228 15108 45240
rect 15160 45228 15166 45280
rect 15381 45271 15439 45277
rect 15381 45237 15393 45271
rect 15427 45268 15439 45271
rect 15562 45268 15568 45280
rect 15427 45240 15568 45268
rect 15427 45237 15439 45240
rect 15381 45231 15439 45237
rect 15562 45228 15568 45240
rect 15620 45228 15626 45280
rect 15933 45271 15991 45277
rect 15933 45237 15945 45271
rect 15979 45268 15991 45271
rect 16850 45268 16856 45280
rect 15979 45240 16856 45268
rect 15979 45237 15991 45240
rect 15933 45231 15991 45237
rect 16850 45228 16856 45240
rect 16908 45228 16914 45280
rect 17236 45268 17264 45376
rect 17313 45373 17325 45407
rect 17359 45404 17371 45407
rect 20625 45407 20683 45413
rect 20625 45404 20637 45407
rect 17359 45376 20637 45404
rect 17359 45373 17371 45376
rect 17313 45367 17371 45373
rect 20625 45373 20637 45376
rect 20671 45404 20683 45407
rect 20714 45404 20720 45416
rect 20671 45376 20720 45404
rect 20671 45373 20683 45376
rect 20625 45367 20683 45373
rect 20714 45364 20720 45376
rect 20772 45364 20778 45416
rect 21269 45407 21327 45413
rect 21269 45373 21281 45407
rect 21315 45373 21327 45407
rect 21376 45404 21404 45444
rect 21453 45407 21511 45413
rect 21453 45404 21465 45407
rect 21376 45376 21465 45404
rect 21269 45367 21327 45373
rect 21453 45373 21465 45376
rect 21499 45373 21511 45407
rect 21545 45407 21603 45413
rect 21545 45394 21557 45407
rect 21591 45394 21603 45407
rect 21453 45367 21511 45373
rect 17580 45339 17638 45345
rect 17580 45305 17592 45339
rect 17626 45336 17638 45339
rect 17954 45336 17960 45348
rect 17626 45308 17960 45336
rect 17626 45305 17638 45308
rect 17580 45299 17638 45305
rect 17954 45296 17960 45308
rect 18012 45296 18018 45348
rect 20380 45339 20438 45345
rect 20380 45305 20392 45339
rect 20426 45336 20438 45339
rect 21174 45336 21180 45348
rect 20426 45308 21180 45336
rect 20426 45305 20438 45308
rect 20380 45299 20438 45305
rect 21174 45296 21180 45308
rect 21232 45296 21238 45348
rect 18506 45268 18512 45280
rect 17236 45240 18512 45268
rect 18506 45228 18512 45240
rect 18564 45228 18570 45280
rect 18690 45268 18696 45280
rect 18651 45240 18696 45268
rect 18690 45228 18696 45240
rect 18748 45228 18754 45280
rect 19245 45271 19303 45277
rect 19245 45237 19257 45271
rect 19291 45268 19303 45271
rect 19334 45268 19340 45280
rect 19291 45240 19340 45268
rect 19291 45237 19303 45240
rect 19245 45231 19303 45237
rect 19334 45228 19340 45240
rect 19392 45268 19398 45280
rect 19794 45268 19800 45280
rect 19392 45240 19800 45268
rect 19392 45228 19398 45240
rect 19794 45228 19800 45240
rect 19852 45228 19858 45280
rect 20162 45228 20168 45280
rect 20220 45268 20226 45280
rect 21284 45268 21312 45367
rect 20220 45240 21312 45268
rect 21468 45268 21496 45367
rect 21542 45342 21548 45394
rect 21600 45342 21606 45394
rect 21634 45364 21640 45416
rect 21692 45404 21698 45416
rect 21836 45413 21864 45444
rect 23385 45441 23397 45475
rect 23431 45472 23443 45475
rect 23492 45472 23520 45500
rect 23750 45472 23756 45484
rect 23431 45444 23520 45472
rect 23584 45444 23756 45472
rect 23431 45441 23443 45444
rect 23385 45435 23443 45441
rect 21821 45407 21879 45413
rect 21692 45376 21772 45404
rect 21692 45364 21698 45376
rect 21744 45336 21772 45376
rect 21821 45373 21833 45407
rect 21867 45373 21879 45407
rect 21821 45367 21879 45373
rect 22281 45407 22339 45413
rect 22281 45373 22293 45407
rect 22327 45373 22339 45407
rect 23106 45404 23112 45416
rect 23067 45376 23112 45404
rect 22281 45367 22339 45373
rect 22296 45336 22324 45367
rect 23106 45364 23112 45376
rect 23164 45364 23170 45416
rect 23290 45364 23296 45416
rect 23348 45406 23354 45416
rect 23477 45407 23535 45413
rect 23348 45378 23391 45406
rect 23348 45364 23354 45378
rect 23477 45373 23489 45407
rect 23523 45404 23535 45407
rect 23584 45404 23612 45444
rect 23750 45432 23756 45444
rect 23808 45432 23814 45484
rect 23523 45376 23612 45404
rect 23661 45407 23719 45413
rect 23523 45373 23535 45376
rect 23477 45367 23535 45373
rect 23661 45373 23673 45407
rect 23707 45373 23719 45407
rect 24320 45404 24348 45580
rect 24412 45580 26148 45608
rect 24412 45481 24440 45580
rect 26142 45568 26148 45580
rect 26200 45568 26206 45620
rect 26234 45568 26240 45620
rect 26292 45608 26298 45620
rect 26292 45580 26337 45608
rect 26292 45568 26298 45580
rect 24397 45475 24455 45481
rect 24397 45441 24409 45475
rect 24443 45441 24455 45475
rect 24397 45435 24455 45441
rect 26142 45432 26148 45484
rect 26200 45472 26206 45484
rect 27614 45472 27620 45484
rect 26200 45444 27620 45472
rect 26200 45432 26206 45444
rect 27614 45432 27620 45444
rect 27672 45432 27678 45484
rect 26789 45407 26847 45413
rect 26789 45404 26801 45407
rect 24320 45376 26801 45404
rect 23661 45367 23719 45373
rect 26789 45373 26801 45376
rect 26835 45404 26847 45407
rect 27522 45404 27528 45416
rect 26835 45376 27528 45404
rect 26835 45373 26847 45376
rect 26789 45367 26847 45373
rect 21744 45308 22324 45336
rect 23667 45336 23695 45367
rect 27522 45364 27528 45376
rect 27580 45364 27586 45416
rect 23845 45339 23903 45345
rect 23667 45308 23796 45336
rect 22186 45268 22192 45280
rect 21468 45240 22192 45268
rect 20220 45228 20226 45240
rect 22186 45228 22192 45240
rect 22244 45228 22250 45280
rect 23768 45268 23796 45308
rect 23845 45305 23857 45339
rect 23891 45336 23903 45339
rect 24642 45339 24700 45345
rect 24642 45336 24654 45339
rect 23891 45308 24654 45336
rect 23891 45305 23903 45308
rect 23845 45299 23903 45305
rect 24642 45305 24654 45308
rect 24688 45305 24700 45339
rect 24642 45299 24700 45305
rect 23934 45268 23940 45280
rect 23768 45240 23940 45268
rect 23934 45228 23940 45240
rect 23992 45268 23998 45280
rect 25777 45271 25835 45277
rect 25777 45268 25789 45271
rect 23992 45240 25789 45268
rect 23992 45228 23998 45240
rect 25777 45237 25789 45240
rect 25823 45268 25835 45271
rect 26050 45268 26056 45280
rect 25823 45240 26056 45268
rect 25823 45237 25835 45240
rect 25777 45231 25835 45237
rect 26050 45228 26056 45240
rect 26108 45228 26114 45280
rect 1104 45178 32016 45200
rect 1104 45126 11253 45178
rect 11305 45126 11317 45178
rect 11369 45126 11381 45178
rect 11433 45126 11445 45178
rect 11497 45126 11509 45178
rect 11561 45126 21557 45178
rect 21609 45126 21621 45178
rect 21673 45126 21685 45178
rect 21737 45126 21749 45178
rect 21801 45126 21813 45178
rect 21865 45126 32016 45178
rect 1104 45104 32016 45126
rect 7190 45064 7196 45076
rect 7151 45036 7196 45064
rect 7190 45024 7196 45036
rect 7248 45024 7254 45076
rect 10686 45024 10692 45076
rect 10744 45064 10750 45076
rect 10744 45036 12388 45064
rect 10744 45024 10750 45036
rect 7282 44956 7288 45008
rect 7340 44996 7346 45008
rect 7558 44996 7564 45008
rect 7340 44968 7564 44996
rect 7340 44956 7346 44968
rect 7558 44956 7564 44968
rect 7616 44996 7622 45008
rect 7616 44968 7972 44996
rect 7616 44956 7622 44968
rect 7377 44931 7435 44937
rect 7377 44897 7389 44931
rect 7423 44928 7435 44931
rect 7466 44928 7472 44940
rect 7423 44900 7472 44928
rect 7423 44897 7435 44900
rect 7377 44891 7435 44897
rect 7466 44888 7472 44900
rect 7524 44888 7530 44940
rect 7742 44928 7748 44940
rect 7703 44900 7748 44928
rect 7742 44888 7748 44900
rect 7800 44888 7806 44940
rect 7944 44937 7972 44968
rect 11146 44956 11152 45008
rect 11204 44996 11210 45008
rect 12253 44999 12311 45005
rect 12253 44996 12265 44999
rect 11204 44968 12265 44996
rect 11204 44956 11210 44968
rect 12253 44965 12265 44968
rect 12299 44965 12311 44999
rect 12253 44959 12311 44965
rect 7929 44931 7987 44937
rect 7929 44897 7941 44931
rect 7975 44897 7987 44931
rect 10226 44928 10232 44940
rect 10187 44900 10232 44928
rect 7929 44891 7987 44897
rect 10226 44888 10232 44900
rect 10284 44888 10290 44940
rect 10413 44931 10471 44937
rect 10413 44897 10425 44931
rect 10459 44928 10471 44931
rect 10686 44928 10692 44940
rect 10459 44900 10692 44928
rect 10459 44897 10471 44900
rect 10413 44891 10471 44897
rect 10686 44888 10692 44900
rect 10744 44888 10750 44940
rect 10781 44931 10839 44937
rect 10781 44897 10793 44931
rect 10827 44928 10839 44931
rect 10870 44928 10876 44940
rect 10827 44900 10876 44928
rect 10827 44897 10839 44900
rect 10781 44891 10839 44897
rect 10870 44888 10876 44900
rect 10928 44888 10934 44940
rect 11701 44931 11759 44937
rect 11701 44897 11713 44931
rect 11747 44897 11759 44931
rect 11701 44891 11759 44897
rect 12161 44931 12219 44937
rect 12161 44897 12173 44931
rect 12207 44928 12219 44931
rect 12360 44928 12388 45036
rect 13630 45024 13636 45076
rect 13688 45064 13694 45076
rect 14826 45064 14832 45076
rect 13688 45036 14832 45064
rect 13688 45024 13694 45036
rect 14826 45024 14832 45036
rect 14884 45024 14890 45076
rect 15746 45064 15752 45076
rect 14936 45036 15752 45064
rect 12207 44900 12388 44928
rect 13541 44931 13599 44937
rect 12207 44897 12219 44900
rect 12161 44891 12219 44897
rect 13541 44897 13553 44931
rect 13587 44928 13599 44931
rect 13630 44928 13636 44940
rect 13587 44900 13636 44928
rect 13587 44897 13599 44900
rect 13541 44891 13599 44897
rect 7190 44820 7196 44872
rect 7248 44860 7254 44872
rect 7561 44863 7619 44869
rect 7561 44860 7573 44863
rect 7248 44832 7573 44860
rect 7248 44820 7254 44832
rect 7561 44829 7573 44832
rect 7607 44829 7619 44863
rect 7561 44823 7619 44829
rect 7650 44820 7656 44872
rect 7708 44860 7714 44872
rect 9125 44863 9183 44869
rect 9125 44860 9137 44863
rect 7708 44832 9137 44860
rect 7708 44820 7714 44832
rect 9125 44829 9137 44832
rect 9171 44829 9183 44863
rect 9125 44823 9183 44829
rect 9306 44820 9312 44872
rect 9364 44860 9370 44872
rect 9401 44863 9459 44869
rect 9401 44860 9413 44863
rect 9364 44832 9413 44860
rect 9364 44820 9370 44832
rect 9401 44829 9413 44832
rect 9447 44829 9459 44863
rect 9401 44823 9459 44829
rect 9950 44820 9956 44872
rect 10008 44860 10014 44872
rect 10502 44860 10508 44872
rect 10008 44832 10508 44860
rect 10008 44820 10014 44832
rect 10502 44820 10508 44832
rect 10560 44820 10566 44872
rect 10594 44820 10600 44872
rect 10652 44860 10658 44872
rect 11716 44860 11744 44891
rect 13630 44888 13636 44900
rect 13688 44888 13694 44940
rect 14642 44928 14648 44940
rect 14603 44900 14648 44928
rect 14642 44888 14648 44900
rect 14700 44888 14706 44940
rect 14737 44931 14795 44937
rect 14737 44897 14749 44931
rect 14783 44928 14795 44931
rect 14936 44928 14964 45036
rect 15746 45024 15752 45036
rect 15804 45024 15810 45076
rect 17034 45024 17040 45076
rect 17092 45064 17098 45076
rect 17954 45064 17960 45076
rect 17092 45036 17816 45064
rect 17915 45036 17960 45064
rect 17092 45024 17098 45036
rect 15102 44956 15108 45008
rect 15160 44996 15166 45008
rect 15160 44968 15700 44996
rect 15160 44956 15166 44968
rect 14783 44900 14964 44928
rect 15013 44931 15071 44937
rect 14783 44897 14795 44900
rect 14737 44891 14795 44897
rect 15013 44897 15025 44931
rect 15059 44897 15071 44931
rect 15470 44928 15476 44940
rect 15431 44900 15476 44928
rect 15013 44891 15071 44897
rect 12618 44860 12624 44872
rect 10652 44832 10697 44860
rect 11716 44832 12624 44860
rect 10652 44820 10658 44832
rect 12618 44820 12624 44832
rect 12676 44820 12682 44872
rect 13446 44820 13452 44872
rect 13504 44860 13510 44872
rect 13817 44863 13875 44869
rect 13817 44860 13829 44863
rect 13504 44832 13829 44860
rect 13504 44820 13510 44832
rect 13817 44829 13829 44832
rect 13863 44829 13875 44863
rect 15028 44860 15056 44891
rect 15470 44888 15476 44900
rect 15528 44888 15534 44940
rect 15672 44937 15700 44968
rect 15657 44931 15715 44937
rect 15657 44897 15669 44931
rect 15703 44897 15715 44931
rect 15657 44891 15715 44897
rect 15746 44888 15752 44940
rect 15804 44928 15810 44940
rect 15804 44900 15849 44928
rect 15804 44888 15810 44900
rect 15930 44888 15936 44940
rect 15988 44928 15994 44940
rect 16025 44931 16083 44937
rect 16025 44928 16037 44931
rect 15988 44900 16037 44928
rect 15988 44888 15994 44900
rect 16025 44897 16037 44900
rect 16071 44897 16083 44931
rect 16025 44891 16083 44897
rect 17126 44888 17132 44940
rect 17184 44928 17190 44940
rect 17221 44931 17279 44937
rect 17221 44928 17233 44931
rect 17184 44900 17233 44928
rect 17184 44888 17190 44900
rect 17221 44897 17233 44900
rect 17267 44897 17279 44931
rect 17221 44891 17279 44897
rect 17405 44931 17463 44937
rect 17405 44897 17417 44931
rect 17451 44928 17463 44931
rect 17678 44928 17684 44940
rect 17451 44900 17684 44928
rect 17451 44897 17463 44900
rect 17405 44891 17463 44897
rect 17678 44888 17684 44900
rect 17736 44888 17742 44940
rect 17788 44937 17816 45036
rect 17954 45024 17960 45036
rect 18012 45024 18018 45076
rect 18506 45064 18512 45076
rect 18467 45036 18512 45064
rect 18506 45024 18512 45036
rect 18564 45024 18570 45076
rect 21174 45024 21180 45076
rect 21232 45064 21238 45076
rect 22557 45067 22615 45073
rect 22557 45064 22569 45067
rect 21232 45036 22569 45064
rect 21232 45024 21238 45036
rect 22557 45033 22569 45036
rect 22603 45033 22615 45067
rect 23382 45064 23388 45076
rect 23295 45036 23388 45064
rect 22557 45027 22615 45033
rect 21266 44956 21272 45008
rect 21324 44996 21330 45008
rect 21324 44968 21404 44996
rect 21324 44956 21330 44968
rect 17773 44931 17831 44937
rect 17773 44897 17785 44931
rect 17819 44897 17831 44931
rect 17773 44891 17831 44897
rect 15838 44860 15844 44872
rect 15028 44832 15844 44860
rect 13817 44823 13875 44829
rect 15838 44820 15844 44832
rect 15896 44820 15902 44872
rect 17494 44860 17500 44872
rect 17455 44832 17500 44860
rect 17494 44820 17500 44832
rect 17552 44820 17558 44872
rect 17586 44820 17592 44872
rect 17644 44860 17650 44872
rect 17788 44860 17816 44891
rect 17862 44888 17868 44940
rect 17920 44928 17926 44940
rect 18601 44931 18659 44937
rect 18601 44928 18613 44931
rect 17920 44900 18613 44928
rect 17920 44888 17926 44900
rect 18601 44897 18613 44900
rect 18647 44897 18659 44931
rect 18601 44891 18659 44897
rect 19061 44931 19119 44937
rect 19061 44897 19073 44931
rect 19107 44897 19119 44931
rect 19794 44928 19800 44940
rect 19707 44900 19800 44928
rect 19061 44891 19119 44897
rect 18690 44860 18696 44872
rect 17644 44832 17689 44860
rect 17788 44832 18696 44860
rect 17644 44820 17650 44832
rect 18690 44820 18696 44832
rect 18748 44860 18754 44872
rect 19076 44860 19104 44891
rect 19794 44888 19800 44900
rect 19852 44888 19858 44940
rect 20993 44931 21051 44937
rect 20993 44897 21005 44931
rect 21039 44928 21051 44931
rect 21376 44928 21404 44968
rect 22094 44956 22100 45008
rect 22152 44996 22158 45008
rect 23325 44996 23353 45036
rect 23382 45024 23388 45036
rect 23440 45064 23446 45076
rect 23440 45036 24072 45064
rect 23440 45024 23446 45036
rect 22152 44968 23353 44996
rect 22152 44956 22158 44968
rect 23474 44956 23480 45008
rect 23532 44996 23538 45008
rect 24044 44996 24072 45036
rect 24118 45024 24124 45076
rect 24176 45064 24182 45076
rect 24176 45036 24221 45064
rect 24176 45024 24182 45036
rect 23532 44968 23704 44996
rect 24044 44968 24900 44996
rect 23532 44956 23538 44968
rect 21039 44900 21404 44928
rect 21039 44897 21051 44900
rect 20993 44891 21051 44897
rect 18748 44832 19104 44860
rect 18748 44820 18754 44832
rect 7668 44792 7696 44820
rect 7392 44764 7696 44792
rect 10965 44795 11023 44801
rect 7392 44736 7420 44764
rect 10965 44761 10977 44795
rect 11011 44792 11023 44795
rect 12342 44792 12348 44804
rect 11011 44764 12348 44792
rect 11011 44761 11023 44764
rect 10965 44755 11023 44761
rect 12342 44752 12348 44764
rect 12400 44752 12406 44804
rect 14461 44795 14519 44801
rect 14461 44761 14473 44795
rect 14507 44792 14519 44795
rect 16114 44792 16120 44804
rect 14507 44764 16120 44792
rect 14507 44761 14519 44764
rect 14461 44755 14519 44761
rect 16114 44752 16120 44764
rect 16172 44752 16178 44804
rect 16666 44752 16672 44804
rect 16724 44792 16730 44804
rect 19153 44795 19211 44801
rect 19153 44792 19165 44795
rect 16724 44764 19165 44792
rect 16724 44752 16730 44764
rect 19153 44761 19165 44764
rect 19199 44761 19211 44795
rect 19812 44792 19840 44888
rect 21082 44820 21088 44872
rect 21140 44860 21146 44872
rect 21269 44863 21327 44869
rect 21269 44860 21281 44863
rect 21140 44832 21281 44860
rect 21140 44820 21146 44832
rect 21269 44829 21281 44832
rect 21315 44829 21327 44863
rect 21376 44860 21404 44900
rect 21450 44888 21456 44940
rect 21508 44928 21514 44940
rect 21821 44931 21879 44937
rect 21821 44928 21833 44931
rect 21508 44900 21833 44928
rect 21508 44888 21514 44900
rect 21821 44897 21833 44900
rect 21867 44897 21879 44931
rect 22002 44928 22008 44940
rect 21963 44900 22008 44928
rect 21821 44891 21879 44897
rect 22002 44888 22008 44900
rect 22060 44888 22066 44940
rect 22186 44928 22192 44940
rect 22147 44900 22192 44928
rect 22186 44888 22192 44900
rect 22244 44888 22250 44940
rect 22373 44931 22431 44937
rect 22373 44897 22385 44931
rect 22419 44897 22431 44931
rect 22373 44891 22431 44897
rect 22097 44863 22155 44869
rect 22097 44860 22109 44863
rect 21376 44832 22109 44860
rect 21269 44823 21327 44829
rect 22097 44829 22109 44832
rect 22143 44829 22155 44863
rect 22097 44823 22155 44829
rect 22388 44792 22416 44891
rect 23106 44888 23112 44940
rect 23164 44928 23170 44940
rect 23676 44937 23704 44968
rect 23385 44931 23443 44937
rect 23385 44928 23397 44931
rect 23164 44900 23397 44928
rect 23164 44888 23170 44900
rect 23385 44897 23397 44900
rect 23431 44897 23443 44931
rect 23557 44929 23615 44935
rect 23557 44926 23569 44929
rect 23385 44891 23443 44897
rect 23492 44898 23569 44926
rect 19812 44764 22416 44792
rect 23492 44792 23520 44898
rect 23557 44895 23569 44898
rect 23603 44895 23615 44929
rect 23557 44889 23615 44895
rect 23655 44931 23713 44937
rect 23655 44897 23667 44931
rect 23701 44897 23713 44931
rect 23655 44891 23713 44897
rect 23937 44931 23995 44937
rect 23937 44897 23949 44931
rect 23983 44928 23995 44931
rect 24394 44928 24400 44940
rect 23983 44900 24400 44928
rect 23983 44897 23995 44900
rect 23937 44891 23995 44897
rect 24394 44888 24400 44900
rect 24452 44888 24458 44940
rect 24486 44888 24492 44940
rect 24544 44928 24550 44940
rect 24872 44937 24900 44968
rect 24581 44931 24639 44937
rect 24581 44928 24593 44931
rect 24544 44900 24593 44928
rect 24544 44888 24550 44900
rect 24581 44897 24593 44900
rect 24627 44897 24639 44931
rect 24581 44891 24639 44897
rect 24857 44931 24915 44937
rect 24857 44897 24869 44931
rect 24903 44897 24915 44931
rect 24857 44891 24915 44897
rect 24949 44931 25007 44937
rect 24949 44897 24961 44931
rect 24995 44928 25007 44931
rect 25682 44928 25688 44940
rect 24995 44900 25688 44928
rect 24995 44897 25007 44900
rect 24949 44891 25007 44897
rect 25682 44888 25688 44900
rect 25740 44888 25746 44940
rect 26418 44888 26424 44940
rect 26476 44928 26482 44940
rect 28086 44931 28144 44937
rect 28086 44928 28098 44931
rect 26476 44900 28098 44928
rect 26476 44888 26482 44900
rect 28086 44897 28098 44900
rect 28132 44897 28144 44931
rect 28086 44891 28144 44897
rect 23750 44860 23756 44872
rect 23711 44832 23756 44860
rect 23750 44820 23756 44832
rect 23808 44820 23814 44872
rect 24210 44820 24216 44872
rect 24268 44860 24274 44872
rect 26145 44863 26203 44869
rect 26145 44860 26157 44863
rect 24268 44832 26157 44860
rect 24268 44820 24274 44832
rect 26145 44829 26157 44832
rect 26191 44829 26203 44863
rect 26145 44823 26203 44829
rect 28353 44863 28411 44869
rect 28353 44829 28365 44863
rect 28399 44829 28411 44863
rect 28353 44823 28411 44829
rect 24302 44792 24308 44804
rect 23492 44764 24308 44792
rect 19153 44755 19211 44761
rect 24302 44752 24308 44764
rect 24360 44752 24366 44804
rect 24762 44752 24768 44804
rect 24820 44792 24826 44804
rect 25593 44795 25651 44801
rect 25593 44792 25605 44795
rect 24820 44764 25605 44792
rect 24820 44752 24826 44764
rect 25593 44761 25605 44764
rect 25639 44761 25651 44795
rect 25593 44755 25651 44761
rect 7374 44684 7380 44736
rect 7432 44684 7438 44736
rect 10134 44684 10140 44736
rect 10192 44724 10198 44736
rect 11609 44727 11667 44733
rect 11609 44724 11621 44727
rect 10192 44696 11621 44724
rect 10192 44684 10198 44696
rect 11609 44693 11621 44696
rect 11655 44693 11667 44727
rect 11609 44687 11667 44693
rect 14921 44727 14979 44733
rect 14921 44693 14933 44727
rect 14967 44724 14979 44727
rect 15930 44724 15936 44736
rect 14967 44696 15936 44724
rect 14967 44693 14979 44696
rect 14921 44687 14979 44693
rect 15930 44684 15936 44696
rect 15988 44724 15994 44736
rect 16206 44724 16212 44736
rect 15988 44696 16212 44724
rect 15988 44684 15994 44696
rect 16206 44684 16212 44696
rect 16264 44684 16270 44736
rect 16761 44727 16819 44733
rect 16761 44693 16773 44727
rect 16807 44724 16819 44727
rect 16942 44724 16948 44736
rect 16807 44696 16948 44724
rect 16807 44693 16819 44696
rect 16761 44687 16819 44693
rect 16942 44684 16948 44696
rect 17000 44684 17006 44736
rect 19889 44727 19947 44733
rect 19889 44693 19901 44727
rect 19935 44724 19947 44727
rect 22370 44724 22376 44736
rect 19935 44696 22376 44724
rect 19935 44693 19947 44696
rect 19889 44687 19947 44693
rect 22370 44684 22376 44696
rect 22428 44684 22434 44736
rect 24026 44684 24032 44736
rect 24084 44724 24090 44736
rect 24673 44727 24731 44733
rect 24673 44724 24685 44727
rect 24084 44696 24685 44724
rect 24084 44684 24090 44696
rect 24673 44693 24685 44696
rect 24719 44693 24731 44727
rect 24673 44687 24731 44693
rect 24854 44684 24860 44736
rect 24912 44724 24918 44736
rect 25133 44727 25191 44733
rect 25133 44724 25145 44727
rect 24912 44696 25145 44724
rect 24912 44684 24918 44696
rect 25133 44693 25145 44696
rect 25179 44693 25191 44727
rect 25133 44687 25191 44693
rect 26326 44684 26332 44736
rect 26384 44724 26390 44736
rect 26973 44727 27031 44733
rect 26973 44724 26985 44727
rect 26384 44696 26985 44724
rect 26384 44684 26390 44696
rect 26973 44693 26985 44696
rect 27019 44693 27031 44727
rect 26973 44687 27031 44693
rect 27614 44684 27620 44736
rect 27672 44724 27678 44736
rect 28368 44724 28396 44823
rect 30926 44724 30932 44736
rect 27672 44696 28396 44724
rect 30887 44696 30932 44724
rect 27672 44684 27678 44696
rect 30926 44684 30932 44696
rect 30984 44684 30990 44736
rect 1104 44634 32016 44656
rect 1104 44582 6102 44634
rect 6154 44582 6166 44634
rect 6218 44582 6230 44634
rect 6282 44582 6294 44634
rect 6346 44582 6358 44634
rect 6410 44582 16405 44634
rect 16457 44582 16469 44634
rect 16521 44582 16533 44634
rect 16585 44582 16597 44634
rect 16649 44582 16661 44634
rect 16713 44582 26709 44634
rect 26761 44582 26773 44634
rect 26825 44582 26837 44634
rect 26889 44582 26901 44634
rect 26953 44582 26965 44634
rect 27017 44582 32016 44634
rect 1104 44560 32016 44582
rect 2682 44480 2688 44532
rect 2740 44520 2746 44532
rect 9769 44523 9827 44529
rect 9769 44520 9781 44523
rect 2740 44492 9781 44520
rect 2740 44480 2746 44492
rect 9769 44489 9781 44492
rect 9815 44489 9827 44523
rect 18046 44520 18052 44532
rect 9769 44483 9827 44489
rect 12084 44492 14136 44520
rect 12084 44464 12112 44492
rect 7006 44412 7012 44464
rect 7064 44452 7070 44464
rect 7193 44455 7251 44461
rect 7193 44452 7205 44455
rect 7064 44424 7205 44452
rect 7064 44412 7070 44424
rect 7193 44421 7205 44424
rect 7239 44452 7251 44455
rect 7742 44452 7748 44464
rect 7239 44424 7748 44452
rect 7239 44421 7251 44424
rect 7193 44415 7251 44421
rect 7742 44412 7748 44424
rect 7800 44412 7806 44464
rect 9490 44412 9496 44464
rect 9548 44452 9554 44464
rect 12066 44452 12072 44464
rect 9548 44424 12072 44452
rect 9548 44412 9554 44424
rect 12066 44412 12072 44424
rect 12124 44412 12130 44464
rect 8297 44387 8355 44393
rect 8297 44353 8309 44387
rect 8343 44384 8355 44387
rect 10594 44384 10600 44396
rect 8343 44356 10600 44384
rect 8343 44353 8355 44356
rect 8297 44347 8355 44353
rect 10594 44344 10600 44356
rect 10652 44344 10658 44396
rect 14108 44393 14136 44492
rect 15672 44492 18052 44520
rect 14093 44387 14151 44393
rect 14093 44353 14105 44387
rect 14139 44353 14151 44387
rect 14093 44347 14151 44353
rect 14274 44344 14280 44396
rect 14332 44384 14338 44396
rect 14369 44387 14427 44393
rect 14369 44384 14381 44387
rect 14332 44356 14381 44384
rect 14332 44344 14338 44356
rect 14369 44353 14381 44356
rect 14415 44384 14427 44387
rect 14458 44384 14464 44396
rect 14415 44356 14464 44384
rect 14415 44353 14427 44356
rect 14369 44347 14427 44353
rect 14458 44344 14464 44356
rect 14516 44344 14522 44396
rect 5810 44316 5816 44328
rect 5771 44288 5816 44316
rect 5810 44276 5816 44288
rect 5868 44276 5874 44328
rect 8018 44316 8024 44328
rect 7979 44288 8024 44316
rect 8018 44276 8024 44288
rect 8076 44276 8082 44328
rect 8113 44319 8171 44325
rect 8113 44285 8125 44319
rect 8159 44285 8171 44319
rect 8386 44316 8392 44328
rect 8347 44288 8392 44316
rect 8113 44279 8171 44285
rect 1854 44248 1860 44260
rect 1815 44220 1860 44248
rect 1854 44208 1860 44220
rect 1912 44208 1918 44260
rect 6080 44251 6138 44257
rect 6080 44217 6092 44251
rect 6126 44248 6138 44251
rect 6822 44248 6828 44260
rect 6126 44220 6828 44248
rect 6126 44217 6138 44220
rect 6080 44211 6138 44217
rect 6822 44208 6828 44220
rect 6880 44208 6886 44260
rect 7926 44248 7932 44260
rect 6932 44220 7932 44248
rect 2133 44183 2191 44189
rect 2133 44149 2145 44183
rect 2179 44180 2191 44183
rect 6932 44180 6960 44220
rect 7926 44208 7932 44220
rect 7984 44208 7990 44260
rect 8128 44248 8156 44279
rect 8386 44276 8392 44288
rect 8444 44276 8450 44328
rect 10502 44316 10508 44328
rect 9140 44288 10508 44316
rect 9140 44248 9168 44288
rect 10502 44276 10508 44288
rect 10560 44276 10566 44328
rect 12069 44319 12127 44325
rect 12069 44285 12081 44319
rect 12115 44316 12127 44319
rect 12158 44316 12164 44328
rect 12115 44288 12164 44316
rect 12115 44285 12127 44288
rect 12069 44279 12127 44285
rect 9858 44248 9864 44260
rect 8128 44220 9168 44248
rect 9819 44220 9864 44248
rect 9858 44208 9864 44220
rect 9916 44208 9922 44260
rect 11606 44248 11612 44260
rect 11567 44220 11612 44248
rect 11606 44208 11612 44220
rect 11664 44248 11670 44260
rect 12084 44248 12112 44279
rect 12158 44276 12164 44288
rect 12216 44276 12222 44328
rect 12342 44325 12348 44328
rect 12336 44316 12348 44325
rect 12303 44288 12348 44316
rect 12336 44279 12348 44288
rect 12342 44276 12348 44279
rect 12400 44276 12406 44328
rect 15470 44316 15476 44328
rect 15431 44288 15476 44316
rect 15470 44276 15476 44288
rect 15528 44276 15534 44328
rect 15672 44325 15700 44492
rect 18046 44480 18052 44492
rect 18104 44480 18110 44532
rect 22554 44480 22560 44532
rect 22612 44520 22618 44532
rect 23750 44520 23756 44532
rect 22612 44492 23756 44520
rect 22612 44480 22618 44492
rect 23750 44480 23756 44492
rect 23808 44480 23814 44532
rect 24118 44480 24124 44532
rect 24176 44520 24182 44532
rect 27985 44523 28043 44529
rect 27985 44520 27997 44523
rect 24176 44492 27997 44520
rect 24176 44480 24182 44492
rect 27985 44489 27997 44492
rect 28031 44489 28043 44523
rect 27985 44483 28043 44489
rect 17126 44452 17132 44464
rect 16868 44424 17132 44452
rect 15841 44387 15899 44393
rect 15841 44353 15853 44387
rect 15887 44384 15899 44387
rect 16206 44384 16212 44396
rect 15887 44356 16212 44384
rect 15887 44353 15899 44356
rect 15841 44347 15899 44353
rect 16206 44344 16212 44356
rect 16264 44344 16270 44396
rect 15657 44319 15715 44325
rect 15657 44285 15669 44319
rect 15703 44285 15715 44319
rect 15657 44279 15715 44285
rect 15746 44276 15752 44328
rect 15804 44316 15810 44328
rect 16022 44316 16028 44328
rect 15804 44288 15849 44316
rect 15983 44288 16028 44316
rect 15804 44276 15810 44288
rect 16022 44276 16028 44288
rect 16080 44276 16086 44328
rect 16868 44325 16896 44424
rect 17126 44412 17132 44424
rect 17184 44412 17190 44464
rect 21450 44452 21456 44464
rect 20732 44424 21456 44452
rect 17586 44384 17592 44396
rect 17328 44356 17592 44384
rect 16853 44319 16911 44325
rect 16853 44285 16865 44319
rect 16899 44285 16911 44319
rect 17034 44316 17040 44328
rect 16995 44288 17040 44316
rect 16853 44279 16911 44285
rect 17034 44276 17040 44288
rect 17092 44276 17098 44328
rect 17129 44319 17187 44325
rect 17129 44285 17141 44319
rect 17175 44285 17187 44319
rect 17129 44279 17187 44285
rect 17221 44319 17279 44325
rect 17221 44285 17233 44319
rect 17267 44316 17279 44319
rect 17328 44316 17356 44356
rect 17586 44344 17592 44356
rect 17644 44384 17650 44396
rect 18414 44384 18420 44396
rect 17644 44356 18420 44384
rect 17644 44344 17650 44356
rect 18414 44344 18420 44356
rect 18472 44344 18478 44396
rect 20732 44393 20760 44424
rect 21450 44412 21456 44424
rect 21508 44412 21514 44464
rect 22830 44412 22836 44464
rect 22888 44452 22894 44464
rect 24210 44452 24216 44464
rect 22888 44424 24216 44452
rect 22888 44412 22894 44424
rect 24210 44412 24216 44424
rect 24268 44412 24274 44464
rect 24486 44452 24492 44464
rect 24447 44424 24492 44452
rect 24486 44412 24492 44424
rect 24544 44412 24550 44464
rect 27062 44412 27068 44464
rect 27120 44452 27126 44464
rect 27522 44452 27528 44464
rect 27120 44424 27528 44452
rect 27120 44412 27126 44424
rect 27522 44412 27528 44424
rect 27580 44452 27586 44464
rect 28537 44455 28595 44461
rect 28537 44452 28549 44455
rect 27580 44424 28549 44452
rect 27580 44412 27586 44424
rect 28537 44421 28549 44424
rect 28583 44452 28595 44455
rect 29362 44452 29368 44464
rect 28583 44424 29368 44452
rect 28583 44421 28595 44424
rect 28537 44415 28595 44421
rect 29362 44412 29368 44424
rect 29420 44412 29426 44464
rect 20717 44387 20775 44393
rect 20717 44353 20729 44387
rect 20763 44353 20775 44387
rect 20717 44347 20775 44353
rect 20993 44387 21051 44393
rect 20993 44353 21005 44387
rect 21039 44384 21051 44387
rect 22094 44384 22100 44396
rect 21039 44356 22100 44384
rect 21039 44353 21051 44356
rect 20993 44347 21051 44353
rect 22094 44344 22100 44356
rect 22152 44344 22158 44396
rect 22186 44344 22192 44396
rect 22244 44384 22250 44396
rect 22649 44387 22707 44393
rect 22649 44384 22661 44387
rect 22244 44356 22661 44384
rect 22244 44344 22250 44356
rect 22649 44353 22661 44356
rect 22695 44353 22707 44387
rect 22649 44347 22707 44353
rect 22848 44356 24348 44384
rect 17267 44288 17356 44316
rect 17405 44319 17463 44325
rect 17267 44285 17279 44288
rect 17221 44279 17279 44285
rect 17405 44285 17417 44319
rect 17451 44316 17463 44319
rect 17954 44316 17960 44328
rect 17451 44288 17960 44316
rect 17451 44285 17463 44288
rect 17405 44279 17463 44285
rect 13906 44248 13912 44260
rect 11664 44220 12112 44248
rect 12176 44220 13912 44248
rect 11664 44208 11670 44220
rect 2179 44152 6960 44180
rect 7837 44183 7895 44189
rect 2179 44149 2191 44152
rect 2133 44143 2191 44149
rect 7837 44149 7849 44183
rect 7883 44180 7895 44183
rect 9122 44180 9128 44192
rect 7883 44152 9128 44180
rect 7883 44149 7895 44152
rect 7837 44143 7895 44149
rect 9122 44140 9128 44152
rect 9180 44140 9186 44192
rect 9214 44140 9220 44192
rect 9272 44180 9278 44192
rect 9769 44183 9827 44189
rect 9272 44152 9317 44180
rect 9272 44140 9278 44152
rect 9769 44149 9781 44183
rect 9815 44180 9827 44183
rect 12176 44180 12204 44220
rect 13906 44208 13912 44220
rect 13964 44248 13970 44260
rect 16942 44248 16948 44260
rect 13964 44220 16948 44248
rect 13964 44208 13970 44220
rect 16942 44208 16948 44220
rect 17000 44208 17006 44260
rect 17144 44248 17172 44279
rect 17954 44276 17960 44288
rect 18012 44316 18018 44328
rect 18233 44319 18291 44325
rect 18233 44316 18245 44319
rect 18012 44288 18245 44316
rect 18012 44276 18018 44288
rect 18233 44285 18245 44288
rect 18279 44285 18291 44319
rect 18233 44279 18291 44285
rect 19245 44319 19303 44325
rect 19245 44285 19257 44319
rect 19291 44285 19303 44319
rect 19245 44279 19303 44285
rect 17144 44220 17264 44248
rect 17236 44192 17264 44220
rect 17310 44208 17316 44260
rect 17368 44248 17374 44260
rect 18141 44251 18199 44257
rect 18141 44248 18153 44251
rect 17368 44220 18153 44248
rect 17368 44208 17374 44220
rect 18141 44217 18153 44220
rect 18187 44217 18199 44251
rect 18141 44211 18199 44217
rect 9815 44152 12204 44180
rect 9815 44149 9827 44152
rect 9769 44143 9827 44149
rect 12250 44140 12256 44192
rect 12308 44180 12314 44192
rect 13449 44183 13507 44189
rect 13449 44180 13461 44183
rect 12308 44152 13461 44180
rect 12308 44140 12314 44152
rect 13449 44149 13461 44152
rect 13495 44149 13507 44183
rect 13449 44143 13507 44149
rect 16209 44183 16267 44189
rect 16209 44149 16221 44183
rect 16255 44180 16267 44183
rect 16390 44180 16396 44192
rect 16255 44152 16396 44180
rect 16255 44149 16267 44152
rect 16209 44143 16267 44149
rect 16390 44140 16396 44152
rect 16448 44140 16454 44192
rect 17218 44140 17224 44192
rect 17276 44140 17282 44192
rect 17586 44180 17592 44192
rect 17547 44152 17592 44180
rect 17586 44140 17592 44152
rect 17644 44140 17650 44192
rect 17678 44140 17684 44192
rect 17736 44180 17742 44192
rect 19260 44180 19288 44279
rect 21266 44276 21272 44328
rect 21324 44316 21330 44328
rect 21453 44319 21511 44325
rect 21453 44316 21465 44319
rect 21324 44288 21465 44316
rect 21324 44276 21330 44288
rect 21453 44285 21465 44288
rect 21499 44316 21511 44319
rect 22002 44316 22008 44328
rect 21499 44288 22008 44316
rect 21499 44285 21511 44288
rect 21453 44279 21511 44285
rect 22002 44276 22008 44288
rect 22060 44276 22066 44328
rect 22465 44319 22523 44325
rect 22465 44285 22477 44319
rect 22511 44285 22523 44319
rect 22738 44316 22744 44328
rect 22699 44288 22744 44316
rect 22465 44279 22523 44285
rect 22480 44248 22508 44279
rect 22738 44276 22744 44288
rect 22796 44276 22802 44328
rect 22848 44325 22876 44356
rect 22833 44319 22891 44325
rect 22833 44285 22845 44319
rect 22879 44285 22891 44319
rect 23014 44316 23020 44328
rect 22975 44288 23020 44316
rect 22833 44279 22891 44285
rect 23014 44276 23020 44288
rect 23072 44276 23078 44328
rect 23658 44316 23664 44328
rect 23619 44288 23664 44316
rect 23658 44276 23664 44288
rect 23716 44276 23722 44328
rect 24210 44248 24216 44260
rect 22480 44220 24216 44248
rect 24210 44208 24216 44220
rect 24268 44208 24274 44260
rect 17736 44152 19288 44180
rect 19337 44183 19395 44189
rect 17736 44140 17742 44152
rect 19337 44149 19349 44183
rect 19383 44180 19395 44183
rect 19426 44180 19432 44192
rect 19383 44152 19432 44180
rect 19383 44149 19395 44152
rect 19337 44143 19395 44149
rect 19426 44140 19432 44152
rect 19484 44140 19490 44192
rect 20622 44140 20628 44192
rect 20680 44180 20686 44192
rect 20806 44180 20812 44192
rect 20680 44152 20812 44180
rect 20680 44140 20686 44152
rect 20806 44140 20812 44152
rect 20864 44140 20870 44192
rect 21450 44140 21456 44192
rect 21508 44180 21514 44192
rect 21545 44183 21603 44189
rect 21545 44180 21557 44183
rect 21508 44152 21557 44180
rect 21508 44140 21514 44152
rect 21545 44149 21557 44152
rect 21591 44149 21603 44183
rect 22278 44180 22284 44192
rect 22239 44152 22284 44180
rect 21545 44143 21603 44149
rect 22278 44140 22284 44152
rect 22336 44140 22342 44192
rect 22370 44140 22376 44192
rect 22428 44180 22434 44192
rect 23569 44183 23627 44189
rect 23569 44180 23581 44183
rect 22428 44152 23581 44180
rect 22428 44140 22434 44152
rect 23569 44149 23581 44152
rect 23615 44149 23627 44183
rect 24320 44180 24348 44356
rect 24397 44319 24455 44325
rect 24397 44285 24409 44319
rect 24443 44316 24455 44319
rect 24578 44316 24584 44328
rect 24443 44288 24584 44316
rect 24443 44285 24455 44288
rect 24397 44279 24455 44285
rect 24578 44276 24584 44288
rect 24636 44276 24642 44328
rect 26973 44319 27031 44325
rect 24964 44288 26924 44316
rect 24964 44180 24992 44288
rect 26602 44208 26608 44260
rect 26660 44248 26666 44260
rect 26706 44251 26764 44257
rect 26706 44248 26718 44251
rect 26660 44220 26718 44248
rect 26660 44208 26666 44220
rect 26706 44217 26718 44220
rect 26752 44217 26764 44251
rect 26896 44248 26924 44288
rect 26973 44285 26985 44319
rect 27019 44316 27031 44319
rect 27614 44316 27620 44328
rect 27019 44288 27620 44316
rect 27019 44285 27031 44288
rect 26973 44279 27031 44285
rect 27614 44276 27620 44288
rect 27672 44276 27678 44328
rect 31110 44316 31116 44328
rect 31071 44288 31116 44316
rect 31110 44276 31116 44288
rect 31168 44276 31174 44328
rect 27338 44248 27344 44260
rect 26896 44220 27344 44248
rect 26706 44211 26764 44217
rect 27338 44208 27344 44220
rect 27396 44208 27402 44260
rect 24320 44152 24992 44180
rect 25133 44183 25191 44189
rect 23569 44143 23627 44149
rect 25133 44149 25145 44183
rect 25179 44180 25191 44183
rect 25314 44180 25320 44192
rect 25179 44152 25320 44180
rect 25179 44149 25191 44152
rect 25133 44143 25191 44149
rect 25314 44140 25320 44152
rect 25372 44140 25378 44192
rect 25593 44183 25651 44189
rect 25593 44149 25605 44183
rect 25639 44180 25651 44183
rect 25866 44180 25872 44192
rect 25639 44152 25872 44180
rect 25639 44149 25651 44152
rect 25593 44143 25651 44149
rect 25866 44140 25872 44152
rect 25924 44140 25930 44192
rect 26234 44140 26240 44192
rect 26292 44180 26298 44192
rect 27433 44183 27491 44189
rect 27433 44180 27445 44183
rect 26292 44152 27445 44180
rect 26292 44140 26298 44152
rect 27433 44149 27445 44152
rect 27479 44149 27491 44183
rect 30650 44180 30656 44192
rect 30611 44152 30656 44180
rect 27433 44143 27491 44149
rect 30650 44140 30656 44152
rect 30708 44140 30714 44192
rect 31297 44183 31355 44189
rect 31297 44149 31309 44183
rect 31343 44180 31355 44183
rect 31343 44152 32076 44180
rect 31343 44149 31355 44152
rect 31297 44143 31355 44149
rect 1104 44090 32016 44112
rect 1104 44038 11253 44090
rect 11305 44038 11317 44090
rect 11369 44038 11381 44090
rect 11433 44038 11445 44090
rect 11497 44038 11509 44090
rect 11561 44038 21557 44090
rect 21609 44038 21621 44090
rect 21673 44038 21685 44090
rect 21737 44038 21749 44090
rect 21801 44038 21813 44090
rect 21865 44038 32016 44090
rect 1104 44016 32016 44038
rect 6822 43976 6828 43988
rect 6783 43948 6828 43976
rect 6822 43936 6828 43948
rect 6880 43936 6886 43988
rect 11793 43979 11851 43985
rect 11793 43945 11805 43979
rect 11839 43976 11851 43979
rect 14642 43976 14648 43988
rect 11839 43948 14648 43976
rect 11839 43945 11851 43948
rect 11793 43939 11851 43945
rect 14642 43936 14648 43948
rect 14700 43936 14706 43988
rect 17218 43936 17224 43988
rect 17276 43976 17282 43988
rect 17276 43948 17724 43976
rect 17276 43936 17282 43948
rect 0 43908 800 43922
rect 1581 43911 1639 43917
rect 1581 43908 1593 43911
rect 0 43880 1593 43908
rect 0 43866 800 43880
rect 1581 43877 1593 43880
rect 1627 43908 1639 43911
rect 1854 43908 1860 43920
rect 1627 43880 1860 43908
rect 1627 43877 1639 43880
rect 1581 43871 1639 43877
rect 1854 43868 1860 43880
rect 1912 43868 1918 43920
rect 12250 43908 12256 43920
rect 10888 43880 12256 43908
rect 10888 43852 10916 43880
rect 12250 43868 12256 43880
rect 12308 43868 12314 43920
rect 14550 43908 14556 43920
rect 12406 43880 14556 43908
rect 7006 43840 7012 43852
rect 6967 43812 7012 43840
rect 7006 43800 7012 43812
rect 7064 43800 7070 43852
rect 7377 43843 7435 43849
rect 7377 43809 7389 43843
rect 7423 43840 7435 43843
rect 7466 43840 7472 43852
rect 7423 43812 7472 43840
rect 7423 43809 7435 43812
rect 7377 43803 7435 43809
rect 7466 43800 7472 43812
rect 7524 43800 7530 43852
rect 7558 43800 7564 43852
rect 7616 43840 7622 43852
rect 8849 43843 8907 43849
rect 7616 43812 7661 43840
rect 7616 43800 7622 43812
rect 8849 43809 8861 43843
rect 8895 43840 8907 43843
rect 9490 43840 9496 43852
rect 8895 43812 9496 43840
rect 8895 43809 8907 43812
rect 8849 43803 8907 43809
rect 9490 43800 9496 43812
rect 9548 43800 9554 43852
rect 10870 43840 10876 43852
rect 10783 43812 10876 43840
rect 10870 43800 10876 43812
rect 10928 43800 10934 43852
rect 11885 43843 11943 43849
rect 11885 43809 11897 43843
rect 11931 43840 11943 43843
rect 12406 43840 12434 43880
rect 14384 43849 14412 43880
rect 14550 43868 14556 43880
rect 14608 43868 14614 43920
rect 15746 43868 15752 43920
rect 15804 43868 15810 43920
rect 16298 43908 16304 43920
rect 15948 43880 16304 43908
rect 11931 43812 12434 43840
rect 12612 43843 12670 43849
rect 11931 43809 11943 43812
rect 11885 43803 11943 43809
rect 12612 43809 12624 43843
rect 12658 43840 12670 43843
rect 14185 43843 14243 43849
rect 14185 43840 14197 43843
rect 12658 43812 14197 43840
rect 12658 43809 12670 43812
rect 12612 43803 12670 43809
rect 14185 43809 14197 43812
rect 14231 43809 14243 43843
rect 14185 43803 14243 43809
rect 14369 43843 14427 43849
rect 14369 43809 14381 43843
rect 14415 43809 14427 43843
rect 14369 43803 14427 43809
rect 14737 43843 14795 43849
rect 14737 43809 14749 43843
rect 14783 43809 14795 43843
rect 14918 43840 14924 43852
rect 14879 43812 14924 43840
rect 14737 43803 14795 43809
rect 7190 43772 7196 43784
rect 7103 43744 7196 43772
rect 7190 43732 7196 43744
rect 7248 43732 7254 43784
rect 7282 43732 7288 43784
rect 7340 43772 7346 43784
rect 8570 43772 8576 43784
rect 7340 43744 7385 43772
rect 8531 43744 8576 43772
rect 7340 43732 7346 43744
rect 8570 43732 8576 43744
rect 8628 43732 8634 43784
rect 9306 43772 9312 43784
rect 9267 43744 9312 43772
rect 9306 43732 9312 43744
rect 9364 43732 9370 43784
rect 9585 43775 9643 43781
rect 9585 43741 9597 43775
rect 9631 43772 9643 43775
rect 9950 43772 9956 43784
rect 9631 43744 9956 43772
rect 9631 43741 9643 43744
rect 9585 43735 9643 43741
rect 9950 43732 9956 43744
rect 10008 43732 10014 43784
rect 11606 43732 11612 43784
rect 11664 43772 11670 43784
rect 12345 43775 12403 43781
rect 12345 43772 12357 43775
rect 11664 43744 12357 43772
rect 11664 43732 11670 43744
rect 12345 43741 12357 43744
rect 12391 43741 12403 43775
rect 12345 43735 12403 43741
rect 7208 43704 7236 43732
rect 8588 43704 8616 43732
rect 7208 43676 8616 43704
rect 13725 43707 13783 43713
rect 13725 43673 13737 43707
rect 13771 43704 13783 43707
rect 14384 43704 14412 43803
rect 14458 43732 14464 43784
rect 14516 43772 14522 43784
rect 14553 43775 14611 43781
rect 14553 43772 14565 43775
rect 14516 43744 14565 43772
rect 14516 43732 14522 43744
rect 14553 43741 14565 43744
rect 14599 43741 14611 43775
rect 14553 43735 14611 43741
rect 14645 43775 14703 43781
rect 14645 43741 14657 43775
rect 14691 43741 14703 43775
rect 14752 43772 14780 43803
rect 14918 43800 14924 43812
rect 14976 43800 14982 43852
rect 15562 43840 15568 43852
rect 15523 43812 15568 43840
rect 15562 43800 15568 43812
rect 15620 43800 15626 43852
rect 15764 43840 15792 43868
rect 15948 43849 15976 43880
rect 16298 43868 16304 43880
rect 16356 43868 16362 43920
rect 17488 43911 17546 43917
rect 17488 43877 17500 43911
rect 17534 43908 17546 43911
rect 17586 43908 17592 43920
rect 17534 43880 17592 43908
rect 17534 43877 17546 43880
rect 17488 43871 17546 43877
rect 17586 43868 17592 43880
rect 17644 43868 17650 43920
rect 17696 43908 17724 43948
rect 17954 43936 17960 43988
rect 18012 43976 18018 43988
rect 18601 43979 18659 43985
rect 18601 43976 18613 43979
rect 18012 43948 18613 43976
rect 18012 43936 18018 43948
rect 18601 43945 18613 43948
rect 18647 43945 18659 43979
rect 18601 43939 18659 43945
rect 20346 43936 20352 43988
rect 20404 43936 20410 43988
rect 24210 43936 24216 43988
rect 24268 43976 24274 43988
rect 24581 43979 24639 43985
rect 24581 43976 24593 43979
rect 24268 43948 24593 43976
rect 24268 43936 24274 43948
rect 24581 43945 24593 43948
rect 24627 43945 24639 43979
rect 26418 43976 26424 43988
rect 26379 43948 26424 43976
rect 24581 43939 24639 43945
rect 26418 43936 26424 43948
rect 26476 43936 26482 43988
rect 29362 43976 29368 43988
rect 29323 43948 29368 43976
rect 29362 43936 29368 43948
rect 29420 43936 29426 43988
rect 20364 43908 20392 43936
rect 24854 43908 24860 43920
rect 17696 43880 19380 43908
rect 20364 43880 20760 43908
rect 15841 43843 15899 43849
rect 15841 43840 15853 43843
rect 15764 43812 15853 43840
rect 15841 43809 15853 43812
rect 15887 43809 15899 43843
rect 15841 43803 15899 43809
rect 15933 43843 15991 43849
rect 15933 43809 15945 43843
rect 15979 43809 15991 43843
rect 16114 43840 16120 43852
rect 16075 43812 16120 43840
rect 15933 43803 15991 43809
rect 16114 43800 16120 43812
rect 16172 43800 16178 43852
rect 16761 43843 16819 43849
rect 16761 43809 16773 43843
rect 16807 43840 16819 43843
rect 18966 43840 18972 43852
rect 16807 43812 18972 43840
rect 16807 43809 16819 43812
rect 16761 43803 16819 43809
rect 18966 43800 18972 43812
rect 19024 43800 19030 43852
rect 19352 43849 19380 43880
rect 19337 43843 19395 43849
rect 19337 43809 19349 43843
rect 19383 43809 19395 43843
rect 19337 43803 19395 43809
rect 20254 43800 20260 43852
rect 20312 43840 20318 43852
rect 20349 43843 20407 43849
rect 20349 43840 20361 43843
rect 20312 43812 20361 43840
rect 20312 43800 20318 43812
rect 20349 43809 20361 43812
rect 20395 43809 20407 43843
rect 20530 43840 20536 43852
rect 20491 43812 20536 43840
rect 20349 43803 20407 43809
rect 20530 43800 20536 43812
rect 20588 43800 20594 43852
rect 20732 43849 20760 43880
rect 22572 43880 24860 43908
rect 20717 43843 20775 43849
rect 20717 43809 20729 43843
rect 20763 43809 20775 43843
rect 20717 43803 20775 43809
rect 20901 43843 20959 43849
rect 20901 43809 20913 43843
rect 20947 43840 20959 43843
rect 21266 43840 21272 43852
rect 20947 43812 21272 43840
rect 20947 43809 20959 43812
rect 20901 43803 20959 43809
rect 21266 43800 21272 43812
rect 21324 43800 21330 43852
rect 21358 43800 21364 43852
rect 21416 43840 21422 43852
rect 22005 43843 22063 43849
rect 22005 43840 22017 43843
rect 21416 43812 22017 43840
rect 21416 43800 21422 43812
rect 22005 43809 22017 43812
rect 22051 43809 22063 43843
rect 22370 43840 22376 43852
rect 22331 43812 22376 43840
rect 22005 43803 22063 43809
rect 22370 43800 22376 43812
rect 22428 43800 22434 43852
rect 22572 43849 22600 43880
rect 24854 43868 24860 43880
rect 24912 43868 24918 43920
rect 32048 43908 32076 44152
rect 32320 43908 33120 43922
rect 32048 43880 33120 43908
rect 32320 43866 33120 43880
rect 22557 43843 22615 43849
rect 22557 43809 22569 43843
rect 22603 43809 22615 43843
rect 22557 43803 22615 43809
rect 23106 43800 23112 43852
rect 23164 43840 23170 43852
rect 23477 43843 23535 43849
rect 23477 43840 23489 43843
rect 23164 43812 23489 43840
rect 23164 43800 23170 43812
rect 23477 43809 23489 43812
rect 23523 43809 23535 43843
rect 23477 43803 23535 43809
rect 24394 43800 24400 43852
rect 24452 43840 24458 43852
rect 24673 43843 24731 43849
rect 24673 43840 24685 43843
rect 24452 43812 24685 43840
rect 24452 43800 24458 43812
rect 24673 43809 24685 43812
rect 24719 43809 24731 43843
rect 25682 43840 25688 43852
rect 25643 43812 25688 43840
rect 24673 43803 24731 43809
rect 25682 43800 25688 43812
rect 25740 43800 25746 43852
rect 25866 43840 25872 43852
rect 25827 43812 25872 43840
rect 25866 43800 25872 43812
rect 25924 43800 25930 43852
rect 26234 43840 26240 43852
rect 26195 43812 26240 43840
rect 26234 43800 26240 43812
rect 26292 43800 26298 43852
rect 27154 43800 27160 43852
rect 27212 43840 27218 43852
rect 27689 43843 27747 43849
rect 27689 43840 27701 43843
rect 27212 43812 27701 43840
rect 27212 43800 27218 43812
rect 27689 43809 27701 43812
rect 27735 43809 27747 43843
rect 27689 43803 27747 43809
rect 15194 43772 15200 43784
rect 14752 43744 15200 43772
rect 14645 43735 14703 43741
rect 14660 43704 14688 43735
rect 15194 43732 15200 43744
rect 15252 43732 15258 43784
rect 15749 43775 15807 43781
rect 15749 43741 15761 43775
rect 15795 43772 15807 43775
rect 16206 43772 16212 43784
rect 15795 43744 16212 43772
rect 15795 43741 15807 43744
rect 15749 43735 15807 43741
rect 16206 43732 16212 43744
rect 16264 43732 16270 43784
rect 17221 43775 17279 43781
rect 17221 43741 17233 43775
rect 17267 43741 17279 43775
rect 17221 43735 17279 43741
rect 19061 43775 19119 43781
rect 19061 43741 19073 43775
rect 19107 43741 19119 43775
rect 19061 43735 19119 43741
rect 13771 43676 14412 43704
rect 14476 43676 14688 43704
rect 13771 43673 13783 43676
rect 13725 43667 13783 43673
rect 14476 43648 14504 43676
rect 15930 43664 15936 43716
rect 15988 43704 15994 43716
rect 16390 43704 16396 43716
rect 15988 43676 16396 43704
rect 15988 43664 15994 43676
rect 16390 43664 16396 43676
rect 16448 43664 16454 43716
rect 2130 43636 2136 43648
rect 2091 43608 2136 43636
rect 2130 43596 2136 43608
rect 2188 43596 2194 43648
rect 5813 43639 5871 43645
rect 5813 43605 5825 43639
rect 5859 43636 5871 43639
rect 6730 43636 6736 43648
rect 5859 43608 6736 43636
rect 5859 43605 5871 43608
rect 5813 43599 5871 43605
rect 6730 43596 6736 43608
rect 6788 43596 6794 43648
rect 10686 43596 10692 43648
rect 10744 43636 10750 43648
rect 10781 43639 10839 43645
rect 10781 43636 10793 43639
rect 10744 43608 10793 43636
rect 10744 43596 10750 43608
rect 10781 43605 10793 43608
rect 10827 43605 10839 43639
rect 10781 43599 10839 43605
rect 14458 43596 14464 43648
rect 14516 43596 14522 43648
rect 15286 43596 15292 43648
rect 15344 43636 15350 43648
rect 15381 43639 15439 43645
rect 15381 43636 15393 43639
rect 15344 43608 15393 43636
rect 15344 43596 15350 43608
rect 15381 43605 15393 43608
rect 15427 43605 15439 43639
rect 17236 43636 17264 43735
rect 19076 43704 19104 43735
rect 20438 43732 20444 43784
rect 20496 43772 20502 43784
rect 20625 43775 20683 43781
rect 20625 43772 20637 43775
rect 20496 43744 20637 43772
rect 20496 43732 20502 43744
rect 20625 43741 20637 43744
rect 20671 43741 20683 43775
rect 20625 43735 20683 43741
rect 21082 43732 21088 43784
rect 21140 43732 21146 43784
rect 22186 43772 22192 43784
rect 22147 43744 22192 43772
rect 22186 43732 22192 43744
rect 22244 43732 22250 43784
rect 22281 43775 22339 43781
rect 22281 43741 22293 43775
rect 22327 43772 22339 43775
rect 22738 43772 22744 43784
rect 22327 43744 22744 43772
rect 22327 43741 22339 43744
rect 22281 43735 22339 43741
rect 22738 43732 22744 43744
rect 22796 43772 22802 43784
rect 22922 43772 22928 43784
rect 22796 43744 22928 43772
rect 22796 43732 22802 43744
rect 22922 43732 22928 43744
rect 22980 43732 22986 43784
rect 23201 43775 23259 43781
rect 23201 43741 23213 43775
rect 23247 43741 23259 43775
rect 23201 43735 23259 43741
rect 21100 43704 21128 43732
rect 19076 43676 21128 43704
rect 22094 43664 22100 43716
rect 22152 43704 22158 43716
rect 23216 43704 23244 43735
rect 23290 43732 23296 43784
rect 23348 43772 23354 43784
rect 24412 43772 24440 43800
rect 23348 43744 24440 43772
rect 25961 43775 26019 43781
rect 23348 43732 23354 43744
rect 25961 43741 25973 43775
rect 26007 43741 26019 43775
rect 25961 43735 26019 43741
rect 26053 43775 26111 43781
rect 26053 43741 26065 43775
rect 26099 43772 26111 43775
rect 26326 43772 26332 43784
rect 26099 43744 26332 43772
rect 26099 43741 26111 43744
rect 26053 43735 26111 43741
rect 22152 43676 23244 43704
rect 25976 43704 26004 43735
rect 26326 43732 26332 43744
rect 26384 43732 26390 43784
rect 27433 43775 27491 43781
rect 27433 43741 27445 43775
rect 27479 43741 27491 43775
rect 27433 43735 27491 43741
rect 26142 43704 26148 43716
rect 25976 43676 26148 43704
rect 22152 43664 22158 43676
rect 26142 43664 26148 43676
rect 26200 43664 26206 43716
rect 18506 43636 18512 43648
rect 17236 43608 18512 43636
rect 15381 43599 15439 43605
rect 18506 43596 18512 43608
rect 18564 43596 18570 43648
rect 20162 43596 20168 43648
rect 20220 43636 20226 43648
rect 21085 43639 21143 43645
rect 21085 43636 21097 43639
rect 20220 43608 21097 43636
rect 20220 43596 20226 43608
rect 21085 43605 21097 43608
rect 21131 43605 21143 43639
rect 21085 43599 21143 43605
rect 21821 43639 21879 43645
rect 21821 43605 21833 43639
rect 21867 43636 21879 43639
rect 23198 43636 23204 43648
rect 21867 43608 23204 43636
rect 21867 43605 21879 43608
rect 21821 43599 21879 43605
rect 23198 43596 23204 43608
rect 23256 43596 23262 43648
rect 25222 43636 25228 43648
rect 25183 43608 25228 43636
rect 25222 43596 25228 43608
rect 25280 43596 25286 43648
rect 27448 43636 27476 43735
rect 27614 43636 27620 43648
rect 27448 43608 27620 43636
rect 27614 43596 27620 43608
rect 27672 43596 27678 43648
rect 28718 43596 28724 43648
rect 28776 43636 28782 43648
rect 28813 43639 28871 43645
rect 28813 43636 28825 43639
rect 28776 43608 28825 43636
rect 28776 43596 28782 43608
rect 28813 43605 28825 43608
rect 28859 43605 28871 43639
rect 28813 43599 28871 43605
rect 30469 43639 30527 43645
rect 30469 43605 30481 43639
rect 30515 43636 30527 43639
rect 31018 43636 31024 43648
rect 30515 43608 31024 43636
rect 30515 43605 30527 43608
rect 30469 43599 30527 43605
rect 31018 43596 31024 43608
rect 31076 43596 31082 43648
rect 1104 43546 32016 43568
rect 1104 43494 6102 43546
rect 6154 43494 6166 43546
rect 6218 43494 6230 43546
rect 6282 43494 6294 43546
rect 6346 43494 6358 43546
rect 6410 43494 16405 43546
rect 16457 43494 16469 43546
rect 16521 43494 16533 43546
rect 16585 43494 16597 43546
rect 16649 43494 16661 43546
rect 16713 43494 26709 43546
rect 26761 43494 26773 43546
rect 26825 43494 26837 43546
rect 26889 43494 26901 43546
rect 26953 43494 26965 43546
rect 27017 43494 32016 43546
rect 1104 43472 32016 43494
rect 5626 43392 5632 43444
rect 5684 43432 5690 43444
rect 5684 43404 9260 43432
rect 5684 43392 5690 43404
rect 9232 43364 9260 43404
rect 9306 43392 9312 43444
rect 9364 43432 9370 43444
rect 9364 43404 12480 43432
rect 9364 43392 9370 43404
rect 10318 43364 10324 43376
rect 9232 43336 10324 43364
rect 10318 43324 10324 43336
rect 10376 43324 10382 43376
rect 5810 43256 5816 43308
rect 5868 43296 5874 43308
rect 5997 43299 6055 43305
rect 5997 43296 6009 43299
rect 5868 43268 6009 43296
rect 5868 43256 5874 43268
rect 5997 43265 6009 43268
rect 6043 43265 6055 43299
rect 9858 43296 9864 43308
rect 5997 43259 6055 43265
rect 8128 43268 9864 43296
rect 8128 43228 8156 43268
rect 9858 43256 9864 43268
rect 9916 43256 9922 43308
rect 9950 43256 9956 43308
rect 10008 43296 10014 43308
rect 12452 43305 12480 43404
rect 15654 43392 15660 43444
rect 15712 43432 15718 43444
rect 17770 43432 17776 43444
rect 15712 43404 17776 43432
rect 15712 43392 15718 43404
rect 17770 43392 17776 43404
rect 17828 43392 17834 43444
rect 23845 43435 23903 43441
rect 23845 43401 23857 43435
rect 23891 43432 23903 43435
rect 24670 43432 24676 43444
rect 23891 43404 24676 43432
rect 23891 43401 23903 43404
rect 23845 43395 23903 43401
rect 24670 43392 24676 43404
rect 24728 43392 24734 43444
rect 27154 43432 27160 43444
rect 27115 43404 27160 43432
rect 27154 43392 27160 43404
rect 27212 43392 27218 43444
rect 30653 43435 30711 43441
rect 30653 43401 30665 43435
rect 30699 43432 30711 43435
rect 30926 43432 30932 43444
rect 30699 43404 30932 43432
rect 30699 43401 30711 43404
rect 30653 43395 30711 43401
rect 30926 43392 30932 43404
rect 30984 43392 30990 43444
rect 31110 43392 31116 43444
rect 31168 43432 31174 43444
rect 31297 43435 31355 43441
rect 31297 43432 31309 43435
rect 31168 43404 31309 43432
rect 31168 43392 31174 43404
rect 31297 43401 31309 43404
rect 31343 43401 31355 43435
rect 31297 43395 31355 43401
rect 21082 43324 21088 43376
rect 21140 43364 21146 43376
rect 21140 43336 22094 43364
rect 21140 43324 21146 43336
rect 10965 43299 11023 43305
rect 10965 43296 10977 43299
rect 10008 43268 10977 43296
rect 10008 43256 10014 43268
rect 10965 43265 10977 43268
rect 11011 43265 11023 43299
rect 10965 43259 11023 43265
rect 12437 43299 12495 43305
rect 12437 43265 12449 43299
rect 12483 43296 12495 43299
rect 12526 43296 12532 43308
rect 12483 43268 12532 43296
rect 12483 43265 12495 43268
rect 12437 43259 12495 43265
rect 12526 43256 12532 43268
rect 12584 43256 12590 43308
rect 12713 43299 12771 43305
rect 12713 43265 12725 43299
rect 12759 43296 12771 43299
rect 14458 43296 14464 43308
rect 12759 43268 14464 43296
rect 12759 43265 12771 43268
rect 12713 43259 12771 43265
rect 14458 43256 14464 43268
rect 14516 43256 14522 43308
rect 16577 43299 16635 43305
rect 16577 43265 16589 43299
rect 16623 43296 16635 43299
rect 16942 43296 16948 43308
rect 16623 43268 16948 43296
rect 16623 43265 16635 43268
rect 16577 43259 16635 43265
rect 16942 43256 16948 43268
rect 17000 43296 17006 43308
rect 17126 43296 17132 43308
rect 17000 43268 17132 43296
rect 17000 43256 17006 43268
rect 17126 43256 17132 43268
rect 17184 43256 17190 43308
rect 18414 43296 18420 43308
rect 18375 43268 18420 43296
rect 18414 43256 18420 43268
rect 18472 43256 18478 43308
rect 20901 43299 20959 43305
rect 20901 43296 20913 43299
rect 19536 43268 20913 43296
rect 4908 43200 8156 43228
rect 8205 43231 8263 43237
rect 1489 43095 1547 43101
rect 1489 43061 1501 43095
rect 1535 43092 1547 43095
rect 1578 43092 1584 43104
rect 1535 43064 1584 43092
rect 1535 43061 1547 43064
rect 1489 43055 1547 43061
rect 1578 43052 1584 43064
rect 1636 43052 1642 43104
rect 1762 43052 1768 43104
rect 1820 43092 1826 43104
rect 1949 43095 2007 43101
rect 1949 43092 1961 43095
rect 1820 43064 1961 43092
rect 1820 43052 1826 43064
rect 1949 43061 1961 43064
rect 1995 43061 2007 43095
rect 1949 43055 2007 43061
rect 2593 43095 2651 43101
rect 2593 43061 2605 43095
rect 2639 43092 2651 43095
rect 2866 43092 2872 43104
rect 2639 43064 2872 43092
rect 2639 43061 2651 43064
rect 2593 43055 2651 43061
rect 2866 43052 2872 43064
rect 2924 43052 2930 43104
rect 2958 43052 2964 43104
rect 3016 43092 3022 43104
rect 3053 43095 3111 43101
rect 3053 43092 3065 43095
rect 3016 43064 3065 43092
rect 3016 43052 3022 43064
rect 3053 43061 3065 43064
rect 3099 43061 3111 43095
rect 3053 43055 3111 43061
rect 4154 43052 4160 43104
rect 4212 43092 4218 43104
rect 4908 43101 4936 43200
rect 8205 43197 8217 43231
rect 8251 43197 8263 43231
rect 8205 43191 8263 43197
rect 6264 43163 6322 43169
rect 6264 43129 6276 43163
rect 6310 43160 6322 43163
rect 7282 43160 7288 43172
rect 6310 43132 7288 43160
rect 6310 43129 6322 43132
rect 6264 43123 6322 43129
rect 7282 43120 7288 43132
rect 7340 43120 7346 43172
rect 8220 43160 8248 43191
rect 9214 43188 9220 43240
rect 9272 43228 9278 43240
rect 9401 43231 9459 43237
rect 9401 43228 9413 43231
rect 9272 43200 9413 43228
rect 9272 43188 9278 43200
rect 9401 43197 9413 43200
rect 9447 43197 9459 43231
rect 9401 43191 9459 43197
rect 9677 43231 9735 43237
rect 9677 43197 9689 43231
rect 9723 43228 9735 43231
rect 10226 43228 10232 43240
rect 9723 43200 10232 43228
rect 9723 43197 9735 43200
rect 9677 43191 9735 43197
rect 10226 43188 10232 43200
rect 10284 43228 10290 43240
rect 10689 43231 10747 43237
rect 10689 43228 10701 43231
rect 10284 43200 10701 43228
rect 10284 43188 10290 43200
rect 10689 43197 10701 43200
rect 10735 43197 10747 43231
rect 10870 43228 10876 43240
rect 10831 43200 10876 43228
rect 10689 43191 10747 43197
rect 10870 43188 10876 43200
rect 10928 43188 10934 43240
rect 11054 43188 11060 43240
rect 11112 43228 11118 43240
rect 11241 43231 11299 43237
rect 11112 43200 11157 43228
rect 11112 43188 11118 43200
rect 11241 43197 11253 43231
rect 11287 43228 11299 43231
rect 11287 43200 12434 43228
rect 11287 43197 11299 43200
rect 11241 43191 11299 43197
rect 7484 43132 8248 43160
rect 7484 43104 7512 43132
rect 11698 43120 11704 43172
rect 11756 43160 11762 43172
rect 11885 43163 11943 43169
rect 11885 43160 11897 43163
rect 11756 43132 11897 43160
rect 11756 43120 11762 43132
rect 11885 43129 11897 43132
rect 11931 43129 11943 43163
rect 12406 43160 12434 43200
rect 14366 43188 14372 43240
rect 14424 43228 14430 43240
rect 15470 43228 15476 43240
rect 14424 43200 15476 43228
rect 14424 43188 14430 43200
rect 15470 43188 15476 43200
rect 15528 43188 15534 43240
rect 15562 43188 15568 43240
rect 15620 43228 15626 43240
rect 16301 43231 16359 43237
rect 16301 43228 16313 43231
rect 15620 43200 16313 43228
rect 15620 43188 15626 43200
rect 16301 43197 16313 43200
rect 16347 43197 16359 43231
rect 16301 43191 16359 43197
rect 18693 43231 18751 43237
rect 18693 43197 18705 43231
rect 18739 43228 18751 43231
rect 19334 43228 19340 43240
rect 18739 43200 19340 43228
rect 18739 43197 18751 43200
rect 18693 43191 18751 43197
rect 19334 43188 19340 43200
rect 19392 43228 19398 43240
rect 19536 43237 19564 43268
rect 20901 43265 20913 43268
rect 20947 43296 20959 43299
rect 22066 43296 22094 43336
rect 26142 43324 26148 43376
rect 26200 43364 26206 43376
rect 26200 43336 26924 43364
rect 26200 43324 26206 43336
rect 22465 43299 22523 43305
rect 22465 43296 22477 43299
rect 20947 43268 21496 43296
rect 22066 43268 22477 43296
rect 20947 43265 20959 43268
rect 20901 43259 20959 43265
rect 19521 43231 19579 43237
rect 19521 43228 19533 43231
rect 19392 43200 19533 43228
rect 19392 43188 19398 43200
rect 19521 43197 19533 43200
rect 19567 43197 19579 43231
rect 19521 43191 19579 43197
rect 20346 43188 20352 43240
rect 20404 43228 20410 43240
rect 21468 43237 21496 43268
rect 22465 43265 22477 43268
rect 22511 43265 22523 43299
rect 22465 43259 22523 43265
rect 22741 43299 22799 43305
rect 22741 43265 22753 43299
rect 22787 43296 22799 43299
rect 23474 43296 23480 43308
rect 22787 43268 23480 43296
rect 22787 43265 22799 43268
rect 22741 43259 22799 43265
rect 23474 43256 23480 43268
rect 23532 43256 23538 43308
rect 23750 43256 23756 43308
rect 23808 43296 23814 43308
rect 23808 43268 24532 43296
rect 23808 43256 23814 43268
rect 20625 43231 20683 43237
rect 20625 43228 20637 43231
rect 20404 43200 20637 43228
rect 20404 43188 20410 43200
rect 20625 43197 20637 43200
rect 20671 43197 20683 43231
rect 20625 43191 20683 43197
rect 21453 43231 21511 43237
rect 21453 43197 21465 43231
rect 21499 43197 21511 43231
rect 24394 43228 24400 43240
rect 24355 43200 24400 43228
rect 21453 43191 21511 43197
rect 24394 43188 24400 43200
rect 24452 43188 24458 43240
rect 24504 43228 24532 43268
rect 26326 43256 26332 43308
rect 26384 43296 26390 43308
rect 26789 43299 26847 43305
rect 26789 43296 26801 43299
rect 26384 43268 26801 43296
rect 26384 43256 26390 43268
rect 26789 43265 26801 43268
rect 26835 43265 26847 43299
rect 26789 43259 26847 43265
rect 26896 43240 26924 43336
rect 26418 43228 26424 43240
rect 24504 43200 24808 43228
rect 26379 43200 26424 43228
rect 12618 43160 12624 43172
rect 12406 43132 12624 43160
rect 11885 43123 11943 43129
rect 12618 43120 12624 43132
rect 12676 43160 12682 43172
rect 13262 43160 13268 43172
rect 12676 43132 13268 43160
rect 12676 43120 12682 43132
rect 13262 43120 13268 43132
rect 13320 43120 13326 43172
rect 15228 43163 15286 43169
rect 15228 43129 15240 43163
rect 15274 43160 15286 43163
rect 15378 43160 15384 43172
rect 15274 43132 15384 43160
rect 15274 43129 15286 43132
rect 15228 43123 15286 43129
rect 15378 43120 15384 43132
rect 15436 43120 15442 43172
rect 22462 43120 22468 43172
rect 22520 43160 22526 43172
rect 24642 43163 24700 43169
rect 24642 43160 24654 43163
rect 22520 43132 24654 43160
rect 22520 43120 22526 43132
rect 24642 43129 24654 43132
rect 24688 43129 24700 43163
rect 24642 43123 24700 43129
rect 4893 43095 4951 43101
rect 4893 43092 4905 43095
rect 4212 43064 4905 43092
rect 4212 43052 4218 43064
rect 4893 43061 4905 43064
rect 4939 43061 4951 43095
rect 4893 43055 4951 43061
rect 5537 43095 5595 43101
rect 5537 43061 5549 43095
rect 5583 43092 5595 43095
rect 5626 43092 5632 43104
rect 5583 43064 5632 43092
rect 5583 43061 5595 43064
rect 5537 43055 5595 43061
rect 5626 43052 5632 43064
rect 5684 43052 5690 43104
rect 7377 43095 7435 43101
rect 7377 43061 7389 43095
rect 7423 43092 7435 43095
rect 7466 43092 7472 43104
rect 7423 43064 7472 43092
rect 7423 43061 7435 43064
rect 7377 43055 7435 43061
rect 7466 43052 7472 43064
rect 7524 43052 7530 43104
rect 8297 43095 8355 43101
rect 8297 43061 8309 43095
rect 8343 43092 8355 43095
rect 9490 43092 9496 43104
rect 8343 43064 9496 43092
rect 8343 43061 8355 43064
rect 8297 43055 8355 43061
rect 9490 43052 9496 43064
rect 9548 43052 9554 43104
rect 11425 43095 11483 43101
rect 11425 43061 11437 43095
rect 11471 43092 11483 43095
rect 11790 43092 11796 43104
rect 11471 43064 11796 43092
rect 11471 43061 11483 43064
rect 11425 43055 11483 43061
rect 11790 43052 11796 43064
rect 11848 43052 11854 43104
rect 14093 43095 14151 43101
rect 14093 43061 14105 43095
rect 14139 43092 14151 43095
rect 15102 43092 15108 43104
rect 14139 43064 15108 43092
rect 14139 43061 14151 43064
rect 14093 43055 14151 43061
rect 15102 43052 15108 43064
rect 15160 43052 15166 43104
rect 17402 43052 17408 43104
rect 17460 43092 17466 43104
rect 19429 43095 19487 43101
rect 19429 43092 19441 43095
rect 17460 43064 19441 43092
rect 17460 43052 17466 43064
rect 19429 43061 19441 43064
rect 19475 43061 19487 43095
rect 19429 43055 19487 43061
rect 21545 43095 21603 43101
rect 21545 43061 21557 43095
rect 21591 43092 21603 43095
rect 22554 43092 22560 43104
rect 21591 43064 22560 43092
rect 21591 43061 21603 43064
rect 21545 43055 21603 43061
rect 22554 43052 22560 43064
rect 22612 43052 22618 43104
rect 22646 43052 22652 43104
rect 22704 43092 22710 43104
rect 23934 43092 23940 43104
rect 22704 43064 23940 43092
rect 22704 43052 22710 43064
rect 23934 43052 23940 43064
rect 23992 43052 23998 43104
rect 24780 43092 24808 43200
rect 26418 43188 26424 43200
rect 26476 43188 26482 43240
rect 26605 43231 26663 43237
rect 26605 43197 26617 43231
rect 26651 43197 26663 43231
rect 26605 43191 26663 43197
rect 26697 43231 26755 43237
rect 26697 43197 26709 43231
rect 26743 43228 26755 43231
rect 26878 43228 26884 43240
rect 26743 43200 26884 43228
rect 26743 43197 26755 43200
rect 26697 43191 26755 43197
rect 26234 43120 26240 43172
rect 26292 43160 26298 43172
rect 26620 43160 26648 43191
rect 26878 43188 26884 43200
rect 26936 43188 26942 43240
rect 26973 43231 27031 43237
rect 26973 43197 26985 43231
rect 27019 43197 27031 43231
rect 27614 43228 27620 43240
rect 27527 43200 27620 43228
rect 26973 43191 27031 43197
rect 26988 43160 27016 43191
rect 27614 43188 27620 43200
rect 27672 43228 27678 43240
rect 28626 43228 28632 43240
rect 27672 43200 28632 43228
rect 27672 43188 27678 43200
rect 28626 43188 28632 43200
rect 28684 43188 28690 43240
rect 31110 43228 31116 43240
rect 31071 43200 31116 43228
rect 31110 43188 31116 43200
rect 31168 43188 31174 43240
rect 27706 43160 27712 43172
rect 26292 43132 26740 43160
rect 26988 43132 27712 43160
rect 26292 43120 26298 43132
rect 25777 43095 25835 43101
rect 25777 43092 25789 43095
rect 24780 43064 25789 43092
rect 25777 43061 25789 43064
rect 25823 43092 25835 43095
rect 26142 43092 26148 43104
rect 25823 43064 26148 43092
rect 25823 43061 25835 43064
rect 25777 43055 25835 43061
rect 26142 43052 26148 43064
rect 26200 43052 26206 43104
rect 26712 43092 26740 43132
rect 27706 43120 27712 43132
rect 27764 43120 27770 43172
rect 27884 43163 27942 43169
rect 27884 43129 27896 43163
rect 27930 43160 27942 43163
rect 28258 43160 28264 43172
rect 27930 43132 28264 43160
rect 27930 43129 27942 43132
rect 27884 43123 27942 43129
rect 28258 43120 28264 43132
rect 28316 43120 28322 43172
rect 27154 43092 27160 43104
rect 26712 43064 27160 43092
rect 27154 43052 27160 43064
rect 27212 43052 27218 43104
rect 28997 43095 29055 43101
rect 28997 43061 29009 43095
rect 29043 43092 29055 43095
rect 29178 43092 29184 43104
rect 29043 43064 29184 43092
rect 29043 43061 29055 43064
rect 28997 43055 29055 43061
rect 29178 43052 29184 43064
rect 29236 43052 29242 43104
rect 29546 43092 29552 43104
rect 29507 43064 29552 43092
rect 29546 43052 29552 43064
rect 29604 43052 29610 43104
rect 1104 43002 32016 43024
rect 1104 42950 11253 43002
rect 11305 42950 11317 43002
rect 11369 42950 11381 43002
rect 11433 42950 11445 43002
rect 11497 42950 11509 43002
rect 11561 42950 21557 43002
rect 21609 42950 21621 43002
rect 21673 42950 21685 43002
rect 21737 42950 21749 43002
rect 21801 42950 21813 43002
rect 21865 42950 32016 43002
rect 1104 42928 32016 42950
rect 9214 42848 9220 42900
rect 9272 42848 9278 42900
rect 9398 42848 9404 42900
rect 9456 42848 9462 42900
rect 9950 42848 9956 42900
rect 10008 42888 10014 42900
rect 15378 42888 15384 42900
rect 10008 42860 15056 42888
rect 15339 42860 15384 42888
rect 10008 42848 10014 42860
rect 9232 42820 9260 42848
rect 8312 42792 9260 42820
rect 9416 42820 9444 42848
rect 11790 42829 11796 42832
rect 11784 42820 11796 42829
rect 9416 42792 9536 42820
rect 5718 42752 5724 42764
rect 5679 42724 5724 42752
rect 5718 42712 5724 42724
rect 5776 42712 5782 42764
rect 7006 42712 7012 42764
rect 7064 42752 7070 42764
rect 7285 42755 7343 42761
rect 7285 42752 7297 42755
rect 7064 42724 7297 42752
rect 7064 42712 7070 42724
rect 7285 42721 7297 42724
rect 7331 42721 7343 42755
rect 7285 42715 7343 42721
rect 7558 42712 7564 42764
rect 7616 42752 7622 42764
rect 8018 42752 8024 42764
rect 7616 42724 8024 42752
rect 7616 42712 7622 42724
rect 8018 42712 8024 42724
rect 8076 42752 8082 42764
rect 8205 42755 8263 42761
rect 8205 42752 8217 42755
rect 8076 42724 8217 42752
rect 8076 42712 8082 42724
rect 8205 42721 8217 42724
rect 8251 42721 8263 42755
rect 8205 42715 8263 42721
rect 4525 42687 4583 42693
rect 4525 42653 4537 42687
rect 4571 42684 4583 42687
rect 5166 42684 5172 42696
rect 4571 42656 5172 42684
rect 4571 42653 4583 42656
rect 4525 42647 4583 42653
rect 5166 42644 5172 42656
rect 5224 42644 5230 42696
rect 5736 42616 5764 42712
rect 6825 42687 6883 42693
rect 6825 42653 6837 42687
rect 6871 42684 6883 42687
rect 7834 42684 7840 42696
rect 6871 42656 7840 42684
rect 6871 42653 6883 42656
rect 6825 42647 6883 42653
rect 7834 42644 7840 42656
rect 7892 42684 7898 42696
rect 7929 42687 7987 42693
rect 7929 42684 7941 42687
rect 7892 42656 7941 42684
rect 7892 42644 7898 42656
rect 7929 42653 7941 42656
rect 7975 42684 7987 42687
rect 8312 42684 8340 42792
rect 9122 42712 9128 42764
rect 9180 42752 9186 42764
rect 9508 42761 9536 42792
rect 10520 42792 10732 42820
rect 11751 42792 11796 42820
rect 10520 42764 10548 42792
rect 9217 42755 9275 42761
rect 9217 42752 9229 42755
rect 9180 42724 9229 42752
rect 9180 42712 9186 42724
rect 9217 42721 9229 42724
rect 9263 42721 9275 42755
rect 9217 42715 9275 42721
rect 9401 42755 9459 42761
rect 9401 42721 9413 42755
rect 9447 42721 9459 42755
rect 9401 42715 9459 42721
rect 9493 42755 9551 42761
rect 9493 42721 9505 42755
rect 9539 42721 9551 42755
rect 9766 42752 9772 42764
rect 9727 42724 9772 42752
rect 9493 42715 9551 42721
rect 7975 42656 8340 42684
rect 7975 42653 7987 42656
rect 7929 42647 7987 42653
rect 7190 42616 7196 42628
rect 5736 42588 7196 42616
rect 7190 42576 7196 42588
rect 7248 42576 7254 42628
rect 9416 42616 9444 42715
rect 9766 42712 9772 42724
rect 9824 42712 9830 42764
rect 10502 42712 10508 42764
rect 10560 42712 10566 42764
rect 10704 42761 10732 42792
rect 11784 42783 11796 42792
rect 11790 42780 11796 42783
rect 11848 42780 11854 42832
rect 14918 42820 14924 42832
rect 14660 42792 14924 42820
rect 10597 42755 10655 42761
rect 10597 42721 10609 42755
rect 10643 42721 10655 42755
rect 10597 42715 10655 42721
rect 10689 42755 10747 42761
rect 10689 42721 10701 42755
rect 10735 42721 10747 42755
rect 10962 42752 10968 42764
rect 10923 42724 10968 42752
rect 10689 42715 10747 42721
rect 9582 42684 9588 42696
rect 9543 42656 9588 42684
rect 9582 42644 9588 42656
rect 9640 42644 9646 42696
rect 10612 42684 10640 42715
rect 10962 42712 10968 42724
rect 11020 42712 11026 42764
rect 11517 42755 11575 42761
rect 11517 42721 11529 42755
rect 11563 42752 11575 42755
rect 11606 42752 11612 42764
rect 11563 42724 11612 42752
rect 11563 42721 11575 42724
rect 11517 42715 11575 42721
rect 11606 42712 11612 42724
rect 11664 42712 11670 42764
rect 12986 42712 12992 42764
rect 13044 42752 13050 42764
rect 14660 42761 14688 42792
rect 14918 42780 14924 42792
rect 14976 42780 14982 42832
rect 15028 42820 15056 42860
rect 15378 42848 15384 42860
rect 15436 42848 15442 42900
rect 22554 42848 22560 42900
rect 22612 42848 22618 42900
rect 23474 42848 23480 42900
rect 23532 42888 23538 42900
rect 28258 42888 28264 42900
rect 23532 42860 23888 42888
rect 28219 42860 28264 42888
rect 23532 42848 23538 42860
rect 20898 42820 20904 42832
rect 15028 42792 20904 42820
rect 20898 42780 20904 42792
rect 20956 42820 20962 42832
rect 21358 42820 21364 42832
rect 20956 42792 21364 42820
rect 20956 42780 20962 42792
rect 21358 42780 21364 42792
rect 21416 42780 21422 42832
rect 22572 42820 22600 42848
rect 23492 42820 23520 42848
rect 22572 42792 22784 42820
rect 13633 42755 13691 42761
rect 13633 42752 13645 42755
rect 13044 42724 13645 42752
rect 13044 42712 13050 42724
rect 13633 42721 13645 42724
rect 13679 42752 13691 42755
rect 14645 42755 14703 42761
rect 14645 42752 14657 42755
rect 13679 42724 14657 42752
rect 13679 42721 13691 42724
rect 13633 42715 13691 42721
rect 14645 42721 14657 42724
rect 14691 42721 14703 42755
rect 14826 42752 14832 42764
rect 14787 42724 14832 42752
rect 14645 42715 14703 42721
rect 14826 42712 14832 42724
rect 14884 42712 14890 42764
rect 15194 42752 15200 42764
rect 15107 42724 15200 42752
rect 15194 42712 15200 42724
rect 15252 42752 15258 42764
rect 15841 42755 15899 42761
rect 15841 42752 15853 42755
rect 15252 42724 15853 42752
rect 15252 42712 15258 42724
rect 15841 42721 15853 42724
rect 15887 42721 15899 42755
rect 16942 42752 16948 42764
rect 16903 42724 16948 42752
rect 15841 42715 15899 42721
rect 16942 42712 16948 42724
rect 17000 42712 17006 42764
rect 17129 42755 17187 42761
rect 17129 42721 17141 42755
rect 17175 42752 17187 42755
rect 17175 42724 17448 42752
rect 17175 42721 17187 42724
rect 17129 42715 17187 42721
rect 11146 42684 11152 42696
rect 10612 42656 11152 42684
rect 11146 42644 11152 42656
rect 11204 42644 11210 42696
rect 13357 42687 13415 42693
rect 13357 42653 13369 42687
rect 13403 42684 13415 42687
rect 13446 42684 13452 42696
rect 13403 42656 13452 42684
rect 13403 42653 13415 42656
rect 13357 42647 13415 42653
rect 13446 42644 13452 42656
rect 13504 42644 13510 42696
rect 14458 42644 14464 42696
rect 14516 42684 14522 42696
rect 14921 42687 14979 42693
rect 14921 42684 14933 42687
rect 14516 42656 14933 42684
rect 14516 42644 14522 42656
rect 14921 42653 14933 42656
rect 14967 42653 14979 42687
rect 14921 42647 14979 42653
rect 15010 42644 15016 42696
rect 15068 42684 15074 42696
rect 17218 42684 17224 42696
rect 15068 42656 15113 42684
rect 17179 42656 17224 42684
rect 15068 42644 15074 42656
rect 17218 42644 17224 42656
rect 17276 42644 17282 42696
rect 17313 42687 17371 42693
rect 17313 42653 17325 42687
rect 17359 42653 17371 42687
rect 17420 42684 17448 42724
rect 17494 42712 17500 42764
rect 17552 42752 17558 42764
rect 17678 42752 17684 42764
rect 17552 42724 17684 42752
rect 17552 42712 17558 42724
rect 17678 42712 17684 42724
rect 17736 42712 17742 42764
rect 18506 42712 18512 42764
rect 18564 42752 18570 42764
rect 18601 42755 18659 42761
rect 18601 42752 18613 42755
rect 18564 42724 18613 42752
rect 18564 42712 18570 42724
rect 18601 42721 18613 42724
rect 18647 42721 18659 42755
rect 18601 42715 18659 42721
rect 18868 42755 18926 42761
rect 18868 42721 18880 42755
rect 18914 42752 18926 42755
rect 19242 42752 19248 42764
rect 18914 42724 19248 42752
rect 18914 42721 18926 42724
rect 18868 42715 18926 42721
rect 19242 42712 19248 42724
rect 19300 42712 19306 42764
rect 19334 42712 19340 42764
rect 19392 42752 19398 42764
rect 20441 42755 20499 42761
rect 20441 42752 20453 42755
rect 19392 42724 20453 42752
rect 19392 42712 19398 42724
rect 20441 42721 20453 42724
rect 20487 42721 20499 42755
rect 20441 42715 20499 42721
rect 22373 42755 22431 42761
rect 22373 42721 22385 42755
rect 22419 42752 22431 42755
rect 22462 42752 22468 42764
rect 22419 42724 22468 42752
rect 22419 42721 22431 42724
rect 22373 42715 22431 42721
rect 22462 42712 22468 42724
rect 22520 42712 22526 42764
rect 22756 42761 22784 42792
rect 22848 42792 23520 42820
rect 22848 42761 22876 42792
rect 23557 42765 23615 42771
rect 22557 42755 22615 42761
rect 22557 42721 22569 42755
rect 22603 42721 22615 42755
rect 22557 42715 22615 42721
rect 22741 42755 22799 42761
rect 22741 42721 22753 42755
rect 22787 42721 22799 42755
rect 22741 42715 22799 42721
rect 22833 42755 22891 42761
rect 22833 42721 22845 42755
rect 22879 42721 22891 42755
rect 22833 42715 22891 42721
rect 22925 42755 22983 42761
rect 22925 42721 22937 42755
rect 22971 42721 22983 42755
rect 23106 42752 23112 42764
rect 23067 42724 23112 42752
rect 22925 42715 22983 42721
rect 17954 42684 17960 42696
rect 17420 42656 17960 42684
rect 17313 42647 17371 42653
rect 10778 42616 10784 42628
rect 9416 42588 10784 42616
rect 10778 42576 10784 42588
rect 10836 42576 10842 42628
rect 13464 42616 13492 42644
rect 15562 42616 15568 42628
rect 13464 42588 15568 42616
rect 15562 42576 15568 42588
rect 15620 42576 15626 42628
rect 15838 42576 15844 42628
rect 15896 42616 15902 42628
rect 15933 42619 15991 42625
rect 15933 42616 15945 42619
rect 15896 42588 15945 42616
rect 15896 42576 15902 42588
rect 15933 42585 15945 42588
rect 15979 42585 15991 42619
rect 17328 42616 17356 42647
rect 17954 42644 17960 42656
rect 18012 42644 18018 42696
rect 20717 42687 20775 42693
rect 20717 42653 20729 42687
rect 20763 42684 20775 42687
rect 20990 42684 20996 42696
rect 20763 42656 20996 42684
rect 20763 42653 20775 42656
rect 20717 42647 20775 42653
rect 20990 42644 20996 42656
rect 21048 42644 21054 42696
rect 17402 42616 17408 42628
rect 17328 42588 17408 42616
rect 15933 42579 15991 42585
rect 17402 42576 17408 42588
rect 17460 42576 17466 42628
rect 20530 42616 20536 42628
rect 19996 42588 20536 42616
rect 1486 42548 1492 42560
rect 1447 42520 1492 42548
rect 1486 42508 1492 42520
rect 1544 42508 1550 42560
rect 2038 42548 2044 42560
rect 1999 42520 2044 42548
rect 2038 42508 2044 42520
rect 2096 42508 2102 42560
rect 2314 42508 2320 42560
rect 2372 42548 2378 42560
rect 2501 42551 2559 42557
rect 2501 42548 2513 42551
rect 2372 42520 2513 42548
rect 2372 42508 2378 42520
rect 2501 42517 2513 42520
rect 2547 42517 2559 42551
rect 3050 42548 3056 42560
rect 3011 42520 3056 42548
rect 2501 42511 2559 42517
rect 3050 42508 3056 42520
rect 3108 42508 3114 42560
rect 3973 42551 4031 42557
rect 3973 42517 3985 42551
rect 4019 42548 4031 42551
rect 4154 42548 4160 42560
rect 4019 42520 4160 42548
rect 4019 42517 4031 42520
rect 3973 42511 4031 42517
rect 4154 42508 4160 42520
rect 4212 42508 4218 42560
rect 4246 42508 4252 42560
rect 4304 42548 4310 42560
rect 5169 42551 5227 42557
rect 5169 42548 5181 42551
rect 4304 42520 5181 42548
rect 4304 42508 4310 42520
rect 5169 42517 5181 42520
rect 5215 42517 5227 42551
rect 5169 42511 5227 42517
rect 7377 42551 7435 42557
rect 7377 42517 7389 42551
rect 7423 42548 7435 42551
rect 9122 42548 9128 42560
rect 7423 42520 9128 42548
rect 7423 42517 7435 42520
rect 7377 42511 7435 42517
rect 9122 42508 9128 42520
rect 9180 42508 9186 42560
rect 9953 42551 10011 42557
rect 9953 42517 9965 42551
rect 9999 42548 10011 42551
rect 10042 42548 10048 42560
rect 9999 42520 10048 42548
rect 9999 42517 10011 42520
rect 9953 42511 10011 42517
rect 10042 42508 10048 42520
rect 10100 42508 10106 42560
rect 10134 42508 10140 42560
rect 10192 42548 10198 42560
rect 10413 42551 10471 42557
rect 10413 42548 10425 42551
rect 10192 42520 10425 42548
rect 10192 42508 10198 42520
rect 10413 42517 10425 42520
rect 10459 42517 10471 42551
rect 10413 42511 10471 42517
rect 10594 42508 10600 42560
rect 10652 42548 10658 42560
rect 10873 42551 10931 42557
rect 10873 42548 10885 42551
rect 10652 42520 10885 42548
rect 10652 42508 10658 42520
rect 10873 42517 10885 42520
rect 10919 42517 10931 42551
rect 10873 42511 10931 42517
rect 12897 42551 12955 42557
rect 12897 42517 12909 42551
rect 12943 42548 12955 42551
rect 13262 42548 13268 42560
rect 12943 42520 13268 42548
rect 12943 42517 12955 42520
rect 12897 42511 12955 42517
rect 13262 42508 13268 42520
rect 13320 42508 13326 42560
rect 16114 42508 16120 42560
rect 16172 42548 16178 42560
rect 17310 42548 17316 42560
rect 16172 42520 17316 42548
rect 16172 42508 16178 42520
rect 17310 42508 17316 42520
rect 17368 42508 17374 42560
rect 17678 42548 17684 42560
rect 17639 42520 17684 42548
rect 17678 42508 17684 42520
rect 17736 42508 17742 42560
rect 19518 42508 19524 42560
rect 19576 42548 19582 42560
rect 19996 42557 20024 42588
rect 20530 42576 20536 42588
rect 20588 42576 20594 42628
rect 22572 42616 22600 42715
rect 22646 42644 22652 42696
rect 22704 42684 22710 42696
rect 22940 42684 22968 42715
rect 23106 42712 23112 42724
rect 23164 42752 23170 42764
rect 23557 42762 23569 42765
rect 23492 42752 23569 42762
rect 23164 42734 23569 42752
rect 23164 42724 23520 42734
rect 23557 42731 23569 42734
rect 23603 42731 23615 42765
rect 23750 42752 23756 42764
rect 23557 42725 23615 42731
rect 23663 42724 23756 42752
rect 23164 42712 23170 42724
rect 23750 42712 23756 42724
rect 23808 42712 23814 42764
rect 23860 42761 23888 42860
rect 28258 42848 28264 42860
rect 28316 42848 28322 42900
rect 27614 42820 27620 42832
rect 26160 42792 27620 42820
rect 23845 42755 23903 42761
rect 23845 42721 23857 42755
rect 23891 42721 23903 42755
rect 23845 42715 23903 42721
rect 24121 42755 24179 42761
rect 24121 42721 24133 42755
rect 24167 42752 24179 42755
rect 24210 42752 24216 42764
rect 24167 42724 24216 42752
rect 24167 42721 24179 42724
rect 24121 42715 24179 42721
rect 24210 42712 24216 42724
rect 24268 42712 24274 42764
rect 25038 42712 25044 42764
rect 25096 42752 25102 42764
rect 26160 42752 26188 42792
rect 27614 42780 27620 42792
rect 27672 42780 27678 42832
rect 28000 42792 28764 42820
rect 25096 42724 26188 42752
rect 25096 42712 25102 42724
rect 26234 42712 26240 42764
rect 26292 42752 26298 42764
rect 27525 42755 27583 42761
rect 27525 42752 27537 42755
rect 26292 42724 26337 42752
rect 26436 42724 27537 42752
rect 26292 42712 26298 42724
rect 23768 42684 23796 42712
rect 26436 42696 26464 42724
rect 27525 42721 27537 42724
rect 27571 42721 27583 42755
rect 27525 42715 27583 42721
rect 27706 42712 27712 42764
rect 27764 42752 27770 42764
rect 28000 42752 28028 42792
rect 28736 42764 28764 42792
rect 27764 42724 28028 42752
rect 28077 42755 28135 42761
rect 27764 42712 27770 42724
rect 28077 42721 28089 42755
rect 28123 42721 28135 42755
rect 28718 42752 28724 42764
rect 28679 42724 28724 42752
rect 28077 42715 28135 42721
rect 22704 42656 22968 42684
rect 23492 42656 23796 42684
rect 23937 42687 23995 42693
rect 22704 42644 22710 42656
rect 23492 42616 23520 42656
rect 23937 42653 23949 42687
rect 23983 42653 23995 42687
rect 23937 42647 23995 42653
rect 22572 42588 23520 42616
rect 23566 42576 23572 42628
rect 23624 42616 23630 42628
rect 23952 42616 23980 42647
rect 24946 42644 24952 42696
rect 25004 42684 25010 42696
rect 25225 42687 25283 42693
rect 25004 42656 25049 42684
rect 25004 42644 25010 42656
rect 25225 42653 25237 42687
rect 25271 42684 25283 42687
rect 25682 42684 25688 42696
rect 25271 42656 25688 42684
rect 25271 42653 25283 42656
rect 25225 42647 25283 42653
rect 25682 42644 25688 42656
rect 25740 42684 25746 42696
rect 26418 42684 26424 42696
rect 25740 42656 26424 42684
rect 25740 42644 25746 42656
rect 26418 42644 26424 42656
rect 26476 42644 26482 42696
rect 26970 42644 26976 42696
rect 27028 42684 27034 42696
rect 27798 42684 27804 42696
rect 27028 42656 27804 42684
rect 27028 42644 27034 42656
rect 27798 42644 27804 42656
rect 27856 42644 27862 42696
rect 27890 42644 27896 42696
rect 27948 42684 27954 42696
rect 28092 42684 28120 42715
rect 28718 42712 28724 42724
rect 28776 42712 28782 42764
rect 29362 42752 29368 42764
rect 29323 42724 29368 42752
rect 29362 42712 29368 42724
rect 29420 42712 29426 42764
rect 30650 42712 30656 42764
rect 30708 42752 30714 42764
rect 30929 42755 30987 42761
rect 30929 42752 30941 42755
rect 30708 42724 30941 42752
rect 30708 42712 30714 42724
rect 30929 42721 30941 42724
rect 30975 42752 30987 42755
rect 31202 42752 31208 42764
rect 30975 42724 31208 42752
rect 30975 42721 30987 42724
rect 30929 42715 30987 42721
rect 31202 42712 31208 42724
rect 31260 42712 31266 42764
rect 29178 42684 29184 42696
rect 27948 42656 27993 42684
rect 28092 42656 29184 42684
rect 27948 42644 27954 42656
rect 29178 42644 29184 42656
rect 29236 42644 29242 42696
rect 29457 42619 29515 42625
rect 29457 42616 29469 42619
rect 23624 42588 23980 42616
rect 24044 42588 24440 42616
rect 23624 42576 23630 42588
rect 19981 42551 20039 42557
rect 19981 42548 19993 42551
rect 19576 42520 19993 42548
rect 19576 42508 19582 42520
rect 19981 42517 19993 42520
rect 20027 42517 20039 42551
rect 19981 42511 20039 42517
rect 20070 42508 20076 42560
rect 20128 42548 20134 42560
rect 21821 42551 21879 42557
rect 21821 42548 21833 42551
rect 20128 42520 21833 42548
rect 20128 42508 20134 42520
rect 21821 42517 21833 42520
rect 21867 42548 21879 42551
rect 22738 42548 22744 42560
rect 21867 42520 22744 42548
rect 21867 42517 21879 42520
rect 21821 42511 21879 42517
rect 22738 42508 22744 42520
rect 22796 42508 22802 42560
rect 23106 42508 23112 42560
rect 23164 42548 23170 42560
rect 24044 42548 24072 42588
rect 24302 42548 24308 42560
rect 23164 42520 24072 42548
rect 24263 42520 24308 42548
rect 23164 42508 23170 42520
rect 24302 42508 24308 42520
rect 24360 42508 24366 42560
rect 24412 42548 24440 42588
rect 25424 42588 29469 42616
rect 25424 42548 25452 42588
rect 29457 42585 29469 42588
rect 29503 42585 29515 42619
rect 29457 42579 29515 42585
rect 26326 42548 26332 42560
rect 24412 42520 25452 42548
rect 26287 42520 26332 42548
rect 26326 42508 26332 42520
rect 26384 42508 26390 42560
rect 26510 42508 26516 42560
rect 26568 42548 26574 42560
rect 26973 42551 27031 42557
rect 26973 42548 26985 42551
rect 26568 42520 26985 42548
rect 26568 42508 26574 42520
rect 26973 42517 26985 42520
rect 27019 42517 27031 42551
rect 26973 42511 27031 42517
rect 27430 42508 27436 42560
rect 27488 42548 27494 42560
rect 28813 42551 28871 42557
rect 28813 42548 28825 42551
rect 27488 42520 28825 42548
rect 27488 42508 27494 42520
rect 28813 42517 28825 42520
rect 28859 42517 28871 42551
rect 28813 42511 28871 42517
rect 30101 42551 30159 42557
rect 30101 42517 30113 42551
rect 30147 42548 30159 42551
rect 30374 42548 30380 42560
rect 30147 42520 30380 42548
rect 30147 42517 30159 42520
rect 30101 42511 30159 42517
rect 30374 42508 30380 42520
rect 30432 42508 30438 42560
rect 1104 42458 32016 42480
rect 1104 42406 6102 42458
rect 6154 42406 6166 42458
rect 6218 42406 6230 42458
rect 6282 42406 6294 42458
rect 6346 42406 6358 42458
rect 6410 42406 16405 42458
rect 16457 42406 16469 42458
rect 16521 42406 16533 42458
rect 16585 42406 16597 42458
rect 16649 42406 16661 42458
rect 16713 42406 26709 42458
rect 26761 42406 26773 42458
rect 26825 42406 26837 42458
rect 26889 42406 26901 42458
rect 26953 42406 26965 42458
rect 27017 42406 32016 42458
rect 1104 42384 32016 42406
rect 4982 42344 4988 42356
rect 4943 42316 4988 42344
rect 4982 42304 4988 42316
rect 5040 42304 5046 42356
rect 7282 42344 7288 42356
rect 7243 42316 7288 42344
rect 7282 42304 7288 42316
rect 7340 42304 7346 42356
rect 9950 42344 9956 42356
rect 7576 42316 9956 42344
rect 3237 42279 3295 42285
rect 3237 42245 3249 42279
rect 3283 42276 3295 42279
rect 7576 42276 7604 42316
rect 9950 42304 9956 42316
rect 10008 42304 10014 42356
rect 10152 42316 10364 42344
rect 3283 42248 7604 42276
rect 3283 42245 3295 42248
rect 3237 42239 3295 42245
rect 7650 42236 7656 42288
rect 7708 42276 7714 42288
rect 8570 42276 8576 42288
rect 7708 42248 8576 42276
rect 7708 42236 7714 42248
rect 8570 42236 8576 42248
rect 8628 42236 8634 42288
rect 9398 42236 9404 42288
rect 9456 42276 9462 42288
rect 10152 42276 10180 42316
rect 9456 42248 10180 42276
rect 9456 42236 9462 42248
rect 3881 42211 3939 42217
rect 3881 42177 3893 42211
rect 3927 42208 3939 42211
rect 5626 42208 5632 42220
rect 3927 42180 5632 42208
rect 3927 42177 3939 42180
rect 3881 42171 3939 42177
rect 5626 42168 5632 42180
rect 5684 42168 5690 42220
rect 7374 42168 7380 42220
rect 7432 42208 7438 42220
rect 7736 42211 7794 42217
rect 7736 42208 7748 42211
rect 7432 42180 7748 42208
rect 7432 42168 7438 42180
rect 7736 42177 7748 42180
rect 7782 42177 7794 42211
rect 7736 42171 7794 42177
rect 9309 42211 9367 42217
rect 9309 42177 9321 42211
rect 9355 42208 9367 42211
rect 10336 42208 10364 42316
rect 11054 42304 11060 42356
rect 11112 42344 11118 42356
rect 11609 42347 11667 42353
rect 11609 42344 11621 42347
rect 11112 42316 11621 42344
rect 11112 42304 11118 42316
rect 11609 42313 11621 42316
rect 11655 42344 11667 42347
rect 11882 42344 11888 42356
rect 11655 42316 11888 42344
rect 11655 42313 11667 42316
rect 11609 42307 11667 42313
rect 11882 42304 11888 42316
rect 11940 42304 11946 42356
rect 19426 42344 19432 42356
rect 17420 42316 19432 42344
rect 13449 42279 13507 42285
rect 13449 42276 13461 42279
rect 12176 42248 13461 42276
rect 12176 42217 12204 42248
rect 13449 42245 13461 42248
rect 13495 42276 13507 42279
rect 16390 42276 16396 42288
rect 13495 42248 15976 42276
rect 13495 42245 13507 42248
rect 13449 42239 13507 42245
rect 10407 42211 10465 42217
rect 10407 42208 10419 42211
rect 9355 42180 9628 42208
rect 10336 42180 10419 42208
rect 9355 42177 9367 42180
rect 9309 42171 9367 42177
rect 1857 42143 1915 42149
rect 1857 42140 1869 42143
rect 768 42112 1869 42140
rect 768 42004 796 42112
rect 1857 42109 1869 42112
rect 1903 42140 1915 42143
rect 2130 42140 2136 42152
rect 1903 42112 2136 42140
rect 1903 42109 1915 42112
rect 1857 42103 1915 42109
rect 2130 42100 2136 42112
rect 2188 42100 2194 42152
rect 2225 42143 2283 42149
rect 2225 42109 2237 42143
rect 2271 42140 2283 42143
rect 5534 42140 5540 42152
rect 2271 42112 5540 42140
rect 2271 42109 2283 42112
rect 2225 42103 2283 42109
rect 5534 42100 5540 42112
rect 5592 42100 5598 42152
rect 6638 42140 6644 42152
rect 6599 42112 6644 42140
rect 6638 42100 6644 42112
rect 6696 42100 6702 42152
rect 7466 42140 7472 42152
rect 7427 42112 7472 42140
rect 7466 42100 7472 42112
rect 7524 42100 7530 42152
rect 7650 42140 7656 42152
rect 7611 42112 7656 42140
rect 7650 42100 7656 42112
rect 7708 42100 7714 42152
rect 7837 42141 7895 42147
rect 7837 42107 7849 42141
rect 7883 42107 7895 42141
rect 8018 42140 8024 42152
rect 7979 42112 8024 42140
rect 7837 42101 7895 42107
rect 5629 42075 5687 42081
rect 5629 42041 5641 42075
rect 5675 42072 5687 42075
rect 6546 42072 6552 42084
rect 5675 42044 6552 42072
rect 5675 42041 5687 42044
rect 5629 42035 5687 42041
rect 6546 42032 6552 42044
rect 6604 42032 6610 42084
rect 7852 42072 7880 42101
rect 8018 42100 8024 42112
rect 8076 42100 8082 42152
rect 8938 42140 8944 42152
rect 8899 42112 8944 42140
rect 8938 42100 8944 42112
rect 8996 42100 9002 42152
rect 9122 42140 9128 42152
rect 9083 42112 9128 42140
rect 9122 42100 9128 42112
rect 9180 42100 9186 42152
rect 9217 42143 9275 42149
rect 9217 42109 9229 42143
rect 9263 42109 9275 42143
rect 9490 42140 9496 42152
rect 9451 42112 9496 42140
rect 9217 42103 9275 42109
rect 8110 42072 8116 42084
rect 7852 42044 8116 42072
rect 8110 42032 8116 42044
rect 8168 42032 8174 42084
rect 9232 42072 9260 42103
rect 9490 42100 9496 42112
rect 9548 42100 9554 42152
rect 9600 42084 9628 42180
rect 10407 42177 10419 42180
rect 10453 42177 10465 42211
rect 10407 42171 10465 42177
rect 12161 42211 12219 42217
rect 12161 42177 12173 42211
rect 12207 42177 12219 42211
rect 12161 42171 12219 42177
rect 13078 42168 13084 42220
rect 13136 42208 13142 42220
rect 14461 42211 14519 42217
rect 14461 42208 14473 42211
rect 13136 42180 14473 42208
rect 13136 42168 13142 42180
rect 14461 42177 14473 42180
rect 14507 42208 14519 42211
rect 15010 42208 15016 42220
rect 14507 42180 15016 42208
rect 14507 42177 14519 42180
rect 14461 42171 14519 42177
rect 15010 42168 15016 42180
rect 15068 42168 15074 42220
rect 10134 42140 10140 42152
rect 10095 42112 10140 42140
rect 10134 42100 10140 42112
rect 10192 42100 10198 42152
rect 10226 42100 10232 42152
rect 10284 42150 10290 42152
rect 10321 42150 10379 42151
rect 10284 42145 10379 42150
rect 10284 42122 10333 42145
rect 10284 42100 10290 42122
rect 10321 42111 10333 42122
rect 10367 42111 10379 42145
rect 10505 42143 10563 42149
rect 10505 42118 10517 42143
rect 10321 42105 10379 42111
rect 10428 42109 10517 42118
rect 10551 42109 10563 42143
rect 10428 42103 10563 42109
rect 10689 42143 10747 42149
rect 10689 42109 10701 42143
rect 10735 42140 10747 42143
rect 10778 42140 10784 42152
rect 10735 42112 10784 42140
rect 10735 42109 10747 42112
rect 10689 42103 10747 42109
rect 10428 42090 10548 42103
rect 10778 42100 10784 42112
rect 10836 42100 10842 42152
rect 11517 42143 11575 42149
rect 11517 42109 11529 42143
rect 11563 42140 11575 42143
rect 12066 42140 12072 42152
rect 11563 42112 12072 42140
rect 11563 42109 11575 42112
rect 11517 42103 11575 42109
rect 12066 42100 12072 42112
rect 12124 42140 12130 42152
rect 12437 42143 12495 42149
rect 12437 42140 12449 42143
rect 12124 42112 12449 42140
rect 12124 42100 12130 42112
rect 12437 42109 12449 42112
rect 12483 42140 12495 42143
rect 13354 42140 13360 42152
rect 12483 42112 13360 42140
rect 12483 42109 12495 42112
rect 12437 42103 12495 42109
rect 13354 42100 13360 42112
rect 13412 42100 13418 42152
rect 14277 42143 14335 42149
rect 14277 42109 14289 42143
rect 14323 42109 14335 42143
rect 14550 42140 14556 42152
rect 14511 42112 14556 42140
rect 14277 42103 14335 42109
rect 9398 42072 9404 42084
rect 9232 42044 9404 42072
rect 9398 42032 9404 42044
rect 9456 42032 9462 42084
rect 9582 42032 9588 42084
rect 9640 42072 9646 42084
rect 10428 42072 10456 42090
rect 9640 42044 10456 42072
rect 9640 42032 9646 42044
rect 12986 42032 12992 42084
rect 13044 42072 13050 42084
rect 14292 42072 14320 42103
rect 14550 42100 14556 42112
rect 14608 42100 14614 42152
rect 14642 42100 14648 42152
rect 14700 42140 14706 42152
rect 14829 42143 14887 42149
rect 14700 42112 14745 42140
rect 14700 42100 14706 42112
rect 14829 42109 14841 42143
rect 14875 42109 14887 42143
rect 14829 42103 14887 42109
rect 14734 42072 14740 42084
rect 13044 42044 14228 42072
rect 14292 42044 14740 42072
rect 13044 42032 13050 42044
rect 4433 42007 4491 42013
rect 768 41976 888 42004
rect 0 41868 800 41882
rect 860 41868 888 41976
rect 4433 41973 4445 42007
rect 4479 42004 4491 42007
rect 4798 42004 4804 42016
rect 4479 41976 4804 42004
rect 4479 41973 4491 41976
rect 4433 41967 4491 41973
rect 4798 41964 4804 41976
rect 4856 41964 4862 42016
rect 5994 41964 6000 42016
rect 6052 42004 6058 42016
rect 6089 42007 6147 42013
rect 6089 42004 6101 42007
rect 6052 41976 6101 42004
rect 6052 41964 6058 41976
rect 6089 41973 6101 41976
rect 6135 41973 6147 42007
rect 6089 41967 6147 41973
rect 6733 42007 6791 42013
rect 6733 41973 6745 42007
rect 6779 42004 6791 42007
rect 9490 42004 9496 42016
rect 6779 41976 9496 42004
rect 6779 41973 6791 41976
rect 6733 41967 6791 41973
rect 9490 41964 9496 41976
rect 9548 41964 9554 42016
rect 9674 42004 9680 42016
rect 9635 41976 9680 42004
rect 9674 41964 9680 41976
rect 9732 41964 9738 42016
rect 10873 42007 10931 42013
rect 10873 41973 10885 42007
rect 10919 42004 10931 42007
rect 10962 42004 10968 42016
rect 10919 41976 10968 42004
rect 10919 41973 10931 41976
rect 10873 41967 10931 41973
rect 10962 41964 10968 41976
rect 11020 41964 11026 42016
rect 13722 41964 13728 42016
rect 13780 42004 13786 42016
rect 14093 42007 14151 42013
rect 14093 42004 14105 42007
rect 13780 41976 14105 42004
rect 13780 41964 13786 41976
rect 14093 41973 14105 41976
rect 14139 41973 14151 42007
rect 14200 42004 14228 42044
rect 14734 42032 14740 42044
rect 14792 42032 14798 42084
rect 14844 42004 14872 42103
rect 15948 42072 15976 42248
rect 16224 42248 16396 42276
rect 16114 42208 16120 42220
rect 16040 42180 16120 42208
rect 16040 42149 16068 42180
rect 16114 42168 16120 42180
rect 16172 42168 16178 42220
rect 16224 42208 16252 42248
rect 16390 42236 16396 42248
rect 16448 42236 16454 42288
rect 16292 42211 16350 42217
rect 16292 42208 16304 42211
rect 16224 42180 16304 42208
rect 16292 42177 16304 42180
rect 16338 42177 16350 42211
rect 17420 42208 17448 42316
rect 19426 42304 19432 42316
rect 19484 42304 19490 42356
rect 21266 42344 21272 42356
rect 21227 42316 21272 42344
rect 21266 42304 21272 42316
rect 21324 42304 21330 42356
rect 22925 42347 22983 42353
rect 22925 42313 22937 42347
rect 22971 42344 22983 42347
rect 23014 42344 23020 42356
rect 22971 42316 23020 42344
rect 22971 42313 22983 42316
rect 22925 42307 22983 42313
rect 23014 42304 23020 42316
rect 23072 42304 23078 42356
rect 26326 42344 26332 42356
rect 24228 42316 26332 42344
rect 23382 42276 23388 42288
rect 22020 42248 22968 42276
rect 23295 42248 23388 42276
rect 16292 42171 16350 42177
rect 16408 42180 17448 42208
rect 18417 42211 18475 42217
rect 16025 42143 16083 42149
rect 16025 42109 16037 42143
rect 16071 42109 16083 42143
rect 16206 42140 16212 42152
rect 16167 42112 16212 42140
rect 16025 42103 16083 42109
rect 16206 42100 16212 42112
rect 16264 42100 16270 42152
rect 16408 42151 16436 42180
rect 18417 42177 18429 42211
rect 18463 42208 18475 42211
rect 18506 42208 18512 42220
rect 18463 42180 18512 42208
rect 18463 42177 18475 42180
rect 18417 42171 18475 42177
rect 18506 42168 18512 42180
rect 18564 42168 18570 42220
rect 21450 42168 21456 42220
rect 21508 42208 21514 42220
rect 22020 42217 22048 42248
rect 22940 42220 22968 42248
rect 23382 42236 23388 42248
rect 23440 42276 23446 42288
rect 24026 42276 24032 42288
rect 23440 42248 24032 42276
rect 23440 42236 23446 42248
rect 24026 42236 24032 42248
rect 24084 42236 24090 42288
rect 22005 42211 22063 42217
rect 21508 42180 21956 42208
rect 21508 42168 21514 42180
rect 16393 42145 16451 42151
rect 16393 42111 16405 42145
rect 16439 42111 16451 42145
rect 16393 42105 16451 42111
rect 16577 42143 16635 42149
rect 16577 42109 16589 42143
rect 16623 42140 16635 42143
rect 16850 42140 16856 42152
rect 16623 42112 16856 42140
rect 16623 42109 16635 42112
rect 16577 42103 16635 42109
rect 16850 42100 16856 42112
rect 16908 42100 16914 42152
rect 17678 42100 17684 42152
rect 17736 42140 17742 42152
rect 18150 42143 18208 42149
rect 18150 42140 18162 42143
rect 17736 42112 18162 42140
rect 17736 42100 17742 42112
rect 18150 42109 18162 42112
rect 18196 42109 18208 42143
rect 18150 42103 18208 42109
rect 19245 42143 19303 42149
rect 19245 42109 19257 42143
rect 19291 42109 19303 42143
rect 19245 42103 19303 42109
rect 19889 42143 19947 42149
rect 19889 42109 19901 42143
rect 19935 42140 19947 42143
rect 20714 42140 20720 42152
rect 19935 42112 20720 42140
rect 19935 42109 19947 42112
rect 19889 42103 19947 42109
rect 15948 42044 17908 42072
rect 15378 42004 15384 42016
rect 14200 41976 14872 42004
rect 15339 41976 15384 42004
rect 14093 41967 14151 41973
rect 15378 41964 15384 41976
rect 15436 41964 15442 42016
rect 15838 42004 15844 42016
rect 15799 41976 15844 42004
rect 15838 41964 15844 41976
rect 15896 41964 15902 42016
rect 16206 41964 16212 42016
rect 16264 42004 16270 42016
rect 16942 42004 16948 42016
rect 16264 41976 16948 42004
rect 16264 41964 16270 41976
rect 16942 41964 16948 41976
rect 17000 41964 17006 42016
rect 17037 42007 17095 42013
rect 17037 41973 17049 42007
rect 17083 42004 17095 42007
rect 17126 42004 17132 42016
rect 17083 41976 17132 42004
rect 17083 41973 17095 41976
rect 17037 41967 17095 41973
rect 17126 41964 17132 41976
rect 17184 42004 17190 42016
rect 17494 42004 17500 42016
rect 17184 41976 17500 42004
rect 17184 41964 17190 41976
rect 17494 41964 17500 41976
rect 17552 41964 17558 42016
rect 17880 42004 17908 42044
rect 17954 42032 17960 42084
rect 18012 42072 18018 42084
rect 19260 42072 19288 42103
rect 20714 42100 20720 42112
rect 20772 42100 20778 42152
rect 21729 42143 21787 42149
rect 21729 42109 21741 42143
rect 21775 42140 21787 42143
rect 21818 42140 21824 42152
rect 21775 42112 21824 42140
rect 21775 42109 21787 42112
rect 21729 42103 21787 42109
rect 21818 42100 21824 42112
rect 21876 42100 21882 42152
rect 21928 42149 21956 42180
rect 22005 42177 22017 42211
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 22097 42211 22155 42217
rect 22097 42177 22109 42211
rect 22143 42208 22155 42211
rect 22186 42208 22192 42220
rect 22143 42180 22192 42208
rect 22143 42177 22155 42180
rect 22097 42171 22155 42177
rect 22186 42168 22192 42180
rect 22244 42208 22250 42220
rect 22830 42208 22836 42220
rect 22244 42180 22836 42208
rect 22244 42168 22250 42180
rect 22830 42168 22836 42180
rect 22888 42168 22894 42220
rect 22922 42168 22928 42220
rect 22980 42168 22986 42220
rect 21913 42143 21971 42149
rect 21913 42109 21925 42143
rect 21959 42109 21971 42143
rect 21913 42103 21971 42109
rect 22292 42143 22350 42149
rect 22292 42109 22304 42143
rect 22338 42140 22350 42143
rect 23106 42140 23112 42152
rect 22338 42112 22968 42140
rect 23067 42112 23112 42140
rect 22338 42109 22350 42112
rect 22292 42103 22350 42109
rect 20162 42081 20168 42084
rect 20156 42072 20168 42081
rect 18012 42044 19288 42072
rect 20123 42044 20168 42072
rect 18012 42032 18018 42044
rect 20156 42035 20168 42044
rect 20162 42032 20168 42035
rect 20220 42032 20226 42084
rect 22940 42072 22968 42112
rect 23106 42100 23112 42112
rect 23164 42100 23170 42152
rect 23201 42143 23259 42149
rect 23201 42109 23213 42143
rect 23247 42140 23259 42143
rect 23290 42140 23296 42152
rect 23247 42112 23296 42140
rect 23247 42109 23259 42112
rect 23201 42103 23259 42109
rect 23290 42100 23296 42112
rect 23348 42100 23354 42152
rect 23477 42143 23535 42149
rect 23477 42109 23489 42143
rect 23523 42140 23535 42143
rect 24228 42140 24256 42316
rect 26326 42304 26332 42316
rect 26384 42304 26390 42356
rect 26602 42304 26608 42356
rect 26660 42344 26666 42356
rect 26973 42347 27031 42353
rect 26973 42344 26985 42347
rect 26660 42316 26985 42344
rect 26660 42304 26666 42316
rect 26973 42313 26985 42316
rect 27019 42313 27031 42347
rect 29362 42344 29368 42356
rect 26973 42307 27031 42313
rect 27080 42316 29368 42344
rect 24394 42140 24400 42152
rect 23523 42112 24256 42140
rect 24307 42112 24400 42140
rect 23523 42109 23535 42112
rect 23477 42103 23535 42109
rect 24394 42100 24400 42112
rect 24452 42140 24458 42152
rect 25038 42140 25044 42152
rect 24452 42112 25044 42140
rect 24452 42100 24458 42112
rect 25038 42100 25044 42112
rect 25096 42100 25102 42152
rect 26234 42100 26240 42152
rect 26292 42130 26298 42152
rect 26425 42145 26483 42151
rect 26694 42149 26700 42152
rect 26425 42130 26437 42145
rect 26471 42130 26483 42145
rect 26292 42102 26327 42130
rect 26292 42100 26298 42102
rect 26237 42099 26249 42100
rect 26283 42099 26295 42100
rect 26237 42093 26295 42099
rect 23934 42072 23940 42084
rect 22940 42044 23940 42072
rect 23934 42032 23940 42044
rect 23992 42032 23998 42084
rect 24302 42032 24308 42084
rect 24360 42072 24366 42084
rect 24642 42075 24700 42081
rect 26418 42078 26424 42130
rect 26476 42105 26483 42130
rect 26513 42143 26571 42149
rect 26513 42109 26525 42143
rect 26559 42109 26571 42143
rect 26476 42078 26482 42105
rect 26513 42103 26571 42109
rect 26651 42143 26700 42149
rect 26651 42109 26663 42143
rect 26697 42109 26700 42143
rect 26651 42103 26700 42109
rect 24642 42072 24654 42075
rect 24360 42044 24654 42072
rect 24360 42032 24366 42044
rect 24642 42041 24654 42044
rect 24688 42041 24700 42075
rect 26528 42072 26556 42103
rect 26694 42100 26700 42103
rect 26752 42100 26758 42152
rect 26786 42100 26792 42152
rect 26844 42140 26850 42152
rect 26844 42112 26889 42140
rect 26844 42100 26850 42112
rect 26878 42072 26884 42084
rect 26528 42044 26884 42072
rect 24642 42035 24700 42041
rect 26878 42032 26884 42044
rect 26936 42032 26942 42084
rect 18598 42004 18604 42016
rect 17880 41976 18604 42004
rect 18598 41964 18604 41976
rect 18656 41964 18662 42016
rect 19337 42007 19395 42013
rect 19337 41973 19349 42007
rect 19383 42004 19395 42007
rect 19518 42004 19524 42016
rect 19383 41976 19524 42004
rect 19383 41973 19395 41976
rect 19337 41967 19395 41973
rect 19518 41964 19524 41976
rect 19576 41964 19582 42016
rect 22186 41964 22192 42016
rect 22244 42004 22250 42016
rect 22465 42007 22523 42013
rect 22465 42004 22477 42007
rect 22244 41976 22477 42004
rect 22244 41964 22250 41976
rect 22465 41973 22477 41976
rect 22511 41973 22523 42007
rect 22465 41967 22523 41973
rect 22554 41964 22560 42016
rect 22612 42004 22618 42016
rect 23382 42004 23388 42016
rect 22612 41976 23388 42004
rect 22612 41964 22618 41976
rect 23382 41964 23388 41976
rect 23440 41964 23446 42016
rect 23658 41964 23664 42016
rect 23716 42004 23722 42016
rect 24210 42004 24216 42016
rect 23716 41976 24216 42004
rect 23716 41964 23722 41976
rect 24210 41964 24216 41976
rect 24268 42004 24274 42016
rect 25777 42007 25835 42013
rect 25777 42004 25789 42007
rect 24268 41976 25789 42004
rect 24268 41964 24274 41976
rect 25777 41973 25789 41976
rect 25823 42004 25835 42007
rect 27080 42004 27108 42316
rect 29362 42304 29368 42316
rect 29420 42304 29426 42356
rect 27890 42236 27896 42288
rect 27948 42276 27954 42288
rect 27948 42248 29960 42276
rect 27948 42236 27954 42248
rect 29932 42220 29960 42248
rect 28902 42168 28908 42220
rect 28960 42208 28966 42220
rect 29825 42211 29883 42217
rect 29825 42208 29837 42211
rect 28960 42180 29837 42208
rect 28960 42168 28966 42180
rect 29825 42177 29837 42180
rect 29871 42177 29883 42211
rect 29825 42171 29883 42177
rect 29914 42168 29920 42220
rect 29972 42208 29978 42220
rect 29972 42180 30065 42208
rect 29972 42168 29978 42180
rect 27154 42100 27160 42152
rect 27212 42140 27218 42152
rect 27433 42143 27491 42149
rect 27433 42140 27445 42143
rect 27212 42112 27445 42140
rect 27212 42100 27218 42112
rect 27433 42109 27445 42112
rect 27479 42109 27491 42143
rect 27433 42103 27491 42109
rect 28261 42143 28319 42149
rect 28261 42109 28273 42143
rect 28307 42109 28319 42143
rect 28261 42103 28319 42109
rect 28997 42143 29055 42149
rect 28997 42109 29009 42143
rect 29043 42140 29055 42143
rect 29086 42140 29092 42152
rect 29043 42112 29092 42140
rect 29043 42109 29055 42112
rect 28997 42103 29055 42109
rect 28169 42075 28227 42081
rect 28169 42072 28181 42075
rect 27356 42044 28181 42072
rect 27356 42016 27384 42044
rect 28169 42041 28181 42044
rect 28215 42041 28227 42075
rect 28276 42072 28304 42103
rect 29086 42100 29092 42112
rect 29144 42100 29150 42152
rect 29270 42100 29276 42152
rect 29328 42140 29334 42152
rect 29549 42143 29607 42149
rect 29549 42140 29561 42143
rect 29328 42112 29561 42140
rect 29328 42100 29334 42112
rect 29549 42109 29561 42112
rect 29595 42109 29607 42143
rect 29549 42103 29607 42109
rect 29733 42143 29791 42149
rect 29733 42109 29745 42143
rect 29779 42109 29791 42143
rect 29733 42103 29791 42109
rect 30101 42143 30159 42149
rect 30101 42109 30113 42143
rect 30147 42140 30159 42143
rect 30466 42140 30472 42152
rect 30147 42112 30472 42140
rect 30147 42109 30159 42112
rect 30101 42103 30159 42109
rect 29104 42072 29132 42100
rect 29748 42072 29776 42103
rect 30466 42100 30472 42112
rect 30524 42100 30530 42152
rect 31110 42140 31116 42152
rect 31071 42112 31116 42140
rect 31110 42100 31116 42112
rect 31168 42100 31174 42152
rect 30006 42072 30012 42084
rect 28276 42044 29040 42072
rect 29104 42044 30012 42072
rect 28169 42035 28227 42041
rect 25823 41976 27108 42004
rect 25823 41973 25835 41976
rect 25777 41967 25835 41973
rect 27338 41964 27344 42016
rect 27396 41964 27402 42016
rect 27522 42004 27528 42016
rect 27483 41976 27528 42004
rect 27522 41964 27528 41976
rect 27580 41964 27586 42016
rect 28258 41964 28264 42016
rect 28316 42004 28322 42016
rect 28905 42007 28963 42013
rect 28905 42004 28917 42007
rect 28316 41976 28917 42004
rect 28316 41964 28322 41976
rect 28905 41973 28917 41976
rect 28951 41973 28963 42007
rect 29012 42004 29040 42044
rect 30006 42032 30012 42044
rect 30064 42032 30070 42084
rect 29178 42004 29184 42016
rect 29012 41976 29184 42004
rect 28905 41967 28963 41973
rect 29178 41964 29184 41976
rect 29236 41964 29242 42016
rect 30282 42004 30288 42016
rect 30243 41976 30288 42004
rect 30282 41964 30288 41976
rect 30340 41964 30346 42016
rect 31297 42007 31355 42013
rect 31297 41973 31309 42007
rect 31343 42004 31355 42007
rect 31343 41976 32076 42004
rect 31343 41973 31355 41976
rect 31297 41967 31355 41973
rect 0 41840 888 41868
rect 1104 41914 32016 41936
rect 1104 41862 11253 41914
rect 11305 41862 11317 41914
rect 11369 41862 11381 41914
rect 11433 41862 11445 41914
rect 11497 41862 11509 41914
rect 11561 41862 21557 41914
rect 21609 41862 21621 41914
rect 21673 41862 21685 41914
rect 21737 41862 21749 41914
rect 21801 41862 21813 41914
rect 21865 41862 32016 41914
rect 1104 41840 32016 41862
rect 32048 41868 32076 41976
rect 32320 41868 33120 41882
rect 32048 41840 33120 41868
rect 0 41826 800 41840
rect 32320 41826 33120 41840
rect 2682 41800 2688 41812
rect 2643 41772 2688 41800
rect 2682 41760 2688 41772
rect 2740 41760 2746 41812
rect 8754 41800 8760 41812
rect 3620 41772 8760 41800
rect 2133 41735 2191 41741
rect 2133 41701 2145 41735
rect 2179 41732 2191 41735
rect 3620 41732 3648 41772
rect 8754 41760 8760 41772
rect 8812 41760 8818 41812
rect 8938 41760 8944 41812
rect 8996 41800 9002 41812
rect 9401 41803 9459 41809
rect 9401 41800 9413 41803
rect 8996 41772 9413 41800
rect 8996 41760 9002 41772
rect 9401 41769 9413 41772
rect 9447 41769 9459 41803
rect 9401 41763 9459 41769
rect 12526 41760 12532 41812
rect 12584 41800 12590 41812
rect 17865 41803 17923 41809
rect 17865 41800 17877 41803
rect 12584 41772 17877 41800
rect 12584 41760 12590 41772
rect 17865 41769 17877 41772
rect 17911 41769 17923 41803
rect 17865 41763 17923 41769
rect 20530 41760 20536 41812
rect 20588 41800 20594 41812
rect 20588 41772 23888 41800
rect 20588 41760 20594 41772
rect 5810 41732 5816 41744
rect 2179 41704 3648 41732
rect 3712 41704 5816 41732
rect 2179 41701 2191 41704
rect 2133 41695 2191 41701
rect 3712 41676 3740 41704
rect 5810 41692 5816 41704
rect 5868 41692 5874 41744
rect 7500 41735 7558 41741
rect 7500 41701 7512 41735
rect 7546 41732 7558 41735
rect 8205 41735 8263 41741
rect 8205 41732 8217 41735
rect 7546 41704 8217 41732
rect 7546 41701 7558 41704
rect 7500 41695 7558 41701
rect 8205 41701 8217 41704
rect 8251 41701 8263 41735
rect 9766 41732 9772 41744
rect 9679 41704 9772 41732
rect 8205 41695 8263 41701
rect 3694 41664 3700 41676
rect 3607 41636 3700 41664
rect 3694 41624 3700 41636
rect 3752 41624 3758 41676
rect 3964 41667 4022 41673
rect 3964 41633 3976 41667
rect 4010 41664 4022 41667
rect 4522 41664 4528 41676
rect 4010 41636 4528 41664
rect 4010 41633 4022 41636
rect 3964 41627 4022 41633
rect 4522 41624 4528 41636
rect 4580 41624 4586 41676
rect 6638 41624 6644 41676
rect 6696 41664 6702 41676
rect 8110 41664 8116 41676
rect 6696 41636 8116 41664
rect 6696 41624 6702 41636
rect 8110 41624 8116 41636
rect 8168 41664 8174 41676
rect 8389 41667 8447 41673
rect 8389 41664 8401 41667
rect 8168 41636 8401 41664
rect 8168 41624 8174 41636
rect 8389 41633 8401 41636
rect 8435 41633 8447 41667
rect 8570 41664 8576 41676
rect 8531 41636 8576 41664
rect 8389 41627 8447 41633
rect 8570 41624 8576 41636
rect 8628 41624 8634 41676
rect 8757 41667 8815 41673
rect 8757 41633 8769 41667
rect 8803 41664 8815 41667
rect 8846 41664 8852 41676
rect 8803 41636 8852 41664
rect 8803 41633 8815 41636
rect 8757 41627 8815 41633
rect 8846 41624 8852 41636
rect 8904 41624 8910 41676
rect 8941 41667 8999 41673
rect 8941 41633 8953 41667
rect 8987 41664 8999 41667
rect 9306 41664 9312 41676
rect 8987 41636 9312 41664
rect 8987 41633 8999 41636
rect 8941 41627 8999 41633
rect 9306 41624 9312 41636
rect 9364 41624 9370 41676
rect 9490 41624 9496 41676
rect 9548 41664 9554 41676
rect 9692 41673 9720 41704
rect 9766 41692 9772 41704
rect 9824 41732 9830 41744
rect 10410 41732 10416 41744
rect 9824 41704 10416 41732
rect 9824 41692 9830 41704
rect 10410 41692 10416 41704
rect 10468 41692 10474 41744
rect 14182 41732 14188 41744
rect 14143 41704 14188 41732
rect 14182 41692 14188 41704
rect 14240 41692 14246 41744
rect 15746 41692 15752 41744
rect 15804 41732 15810 41744
rect 16298 41732 16304 41744
rect 15804 41704 16304 41732
rect 15804 41692 15810 41704
rect 16298 41692 16304 41704
rect 16356 41732 16362 41744
rect 16356 41704 16988 41732
rect 16356 41692 16362 41704
rect 9585 41667 9643 41673
rect 9585 41664 9597 41667
rect 9548 41636 9597 41664
rect 9548 41624 9554 41636
rect 9585 41633 9597 41636
rect 9631 41633 9643 41667
rect 9585 41627 9643 41633
rect 9677 41667 9735 41673
rect 9677 41633 9689 41667
rect 9723 41633 9735 41667
rect 9677 41627 9735 41633
rect 9953 41667 10011 41673
rect 9953 41633 9965 41667
rect 9999 41633 10011 41667
rect 9953 41627 10011 41633
rect 5350 41556 5356 41608
rect 5408 41596 5414 41608
rect 5721 41599 5779 41605
rect 5721 41596 5733 41599
rect 5408 41568 5733 41596
rect 5408 41556 5414 41568
rect 5721 41565 5733 41568
rect 5767 41565 5779 41599
rect 5721 41559 5779 41565
rect 7745 41599 7803 41605
rect 7745 41565 7757 41599
rect 7791 41596 7803 41599
rect 8294 41596 8300 41608
rect 7791 41568 8300 41596
rect 7791 41565 7803 41568
rect 7745 41559 7803 41565
rect 8294 41556 8300 41568
rect 8352 41556 8358 41608
rect 8662 41556 8668 41608
rect 8720 41596 8726 41608
rect 8720 41568 8765 41596
rect 8720 41556 8726 41568
rect 9214 41556 9220 41608
rect 9272 41596 9278 41608
rect 9968 41596 9996 41627
rect 10042 41624 10048 41676
rect 10100 41664 10106 41676
rect 10781 41667 10839 41673
rect 10781 41664 10793 41667
rect 10100 41636 10793 41664
rect 10100 41624 10106 41636
rect 10781 41633 10793 41636
rect 10827 41633 10839 41667
rect 10781 41627 10839 41633
rect 12069 41667 12127 41673
rect 12069 41633 12081 41667
rect 12115 41664 12127 41667
rect 12802 41664 12808 41676
rect 12115 41636 12808 41664
rect 12115 41633 12127 41636
rect 12069 41627 12127 41633
rect 12802 41624 12808 41636
rect 12860 41624 12866 41676
rect 13078 41664 13084 41676
rect 13039 41636 13084 41664
rect 13078 41624 13084 41636
rect 13136 41624 13142 41676
rect 13354 41664 13360 41676
rect 13315 41636 13360 41664
rect 13354 41624 13360 41636
rect 13412 41624 13418 41676
rect 16206 41624 16212 41676
rect 16264 41664 16270 41676
rect 16960 41673 16988 41704
rect 17310 41692 17316 41744
rect 17368 41732 17374 41744
rect 22189 41735 22247 41741
rect 17368 41704 21036 41732
rect 17368 41692 17374 41704
rect 16669 41667 16727 41673
rect 16669 41664 16681 41667
rect 16264 41636 16681 41664
rect 16264 41624 16270 41636
rect 16669 41633 16681 41636
rect 16715 41633 16727 41667
rect 16669 41627 16727 41633
rect 16853 41667 16911 41673
rect 16853 41633 16865 41667
rect 16899 41633 16911 41667
rect 16853 41627 16911 41633
rect 16945 41667 17003 41673
rect 16945 41633 16957 41667
rect 16991 41633 17003 41667
rect 16945 41627 17003 41633
rect 17221 41667 17279 41673
rect 17221 41633 17233 41667
rect 17267 41633 17279 41667
rect 17221 41627 17279 41633
rect 18969 41667 19027 41673
rect 18969 41633 18981 41667
rect 19015 41664 19027 41667
rect 19334 41664 19340 41676
rect 19015 41636 19340 41664
rect 19015 41633 19027 41636
rect 18969 41627 19027 41633
rect 9272 41568 9996 41596
rect 9272 41556 9278 41568
rect 10318 41556 10324 41608
rect 10376 41596 10382 41608
rect 10689 41599 10747 41605
rect 10689 41596 10701 41599
rect 10376 41568 10701 41596
rect 10376 41556 10382 41568
rect 10689 41565 10701 41568
rect 10735 41565 10747 41599
rect 10689 41559 10747 41565
rect 12618 41556 12624 41608
rect 12676 41596 12682 41608
rect 13096 41596 13124 41624
rect 12676 41568 13124 41596
rect 12676 41556 12682 41568
rect 15194 41556 15200 41608
rect 15252 41596 15258 41608
rect 16868 41596 16896 41627
rect 17034 41596 17040 41608
rect 15252 41568 16896 41596
rect 16995 41568 17040 41596
rect 15252 41556 15258 41568
rect 17034 41556 17040 41568
rect 17092 41556 17098 41608
rect 6365 41531 6423 41537
rect 4632 41500 6040 41528
rect 1581 41463 1639 41469
rect 1581 41429 1593 41463
rect 1627 41460 1639 41463
rect 1854 41460 1860 41472
rect 1627 41432 1860 41460
rect 1627 41429 1639 41432
rect 1581 41423 1639 41429
rect 1854 41420 1860 41432
rect 1912 41420 1918 41472
rect 3234 41460 3240 41472
rect 3147 41432 3240 41460
rect 3234 41420 3240 41432
rect 3292 41460 3298 41472
rect 4632 41460 4660 41500
rect 3292 41432 4660 41460
rect 5077 41463 5135 41469
rect 3292 41420 3298 41432
rect 5077 41429 5089 41463
rect 5123 41460 5135 41463
rect 5626 41460 5632 41472
rect 5123 41432 5632 41460
rect 5123 41429 5135 41432
rect 5077 41423 5135 41429
rect 5626 41420 5632 41432
rect 5684 41420 5690 41472
rect 6012 41460 6040 41500
rect 6365 41497 6377 41531
rect 6411 41528 6423 41531
rect 6638 41528 6644 41540
rect 6411 41500 6644 41528
rect 6411 41497 6423 41500
rect 6365 41491 6423 41497
rect 6638 41488 6644 41500
rect 6696 41488 6702 41540
rect 10134 41528 10140 41540
rect 7760 41500 10140 41528
rect 7760 41460 7788 41500
rect 10134 41488 10140 41500
rect 10192 41488 10198 41540
rect 10594 41528 10600 41540
rect 10244 41500 10600 41528
rect 9858 41460 9864 41472
rect 6012 41432 7788 41460
rect 9771 41432 9864 41460
rect 9858 41420 9864 41432
rect 9916 41460 9922 41472
rect 10244 41460 10272 41500
rect 10594 41488 10600 41500
rect 10652 41488 10658 41540
rect 11977 41531 12035 41537
rect 11977 41497 11989 41531
rect 12023 41528 12035 41531
rect 17236 41528 17264 41627
rect 19334 41624 19340 41636
rect 19392 41624 19398 41676
rect 20254 41664 20260 41676
rect 20215 41636 20260 41664
rect 20254 41624 20260 41636
rect 20312 41624 20318 41676
rect 21008 41673 21036 41704
rect 22189 41701 22201 41735
rect 22235 41732 22247 41735
rect 23290 41732 23296 41744
rect 22235 41704 23296 41732
rect 22235 41701 22247 41704
rect 22189 41695 22247 41701
rect 23290 41692 23296 41704
rect 23348 41692 23354 41744
rect 20993 41667 21051 41673
rect 20993 41633 21005 41667
rect 21039 41633 21051 41667
rect 20993 41627 21051 41633
rect 21266 41624 21272 41676
rect 21324 41664 21330 41676
rect 21821 41667 21879 41673
rect 21821 41664 21833 41667
rect 21324 41636 21833 41664
rect 21324 41624 21330 41636
rect 21821 41633 21833 41636
rect 21867 41633 21879 41667
rect 21821 41627 21879 41633
rect 22005 41667 22063 41673
rect 22005 41633 22017 41667
rect 22051 41633 22063 41667
rect 22005 41627 22063 41633
rect 18598 41556 18604 41608
rect 18656 41596 18662 41608
rect 19245 41599 19303 41605
rect 19245 41596 19257 41599
rect 18656 41568 19257 41596
rect 18656 41556 18662 41568
rect 19245 41565 19257 41568
rect 19291 41565 19303 41599
rect 19245 41559 19303 41565
rect 20533 41599 20591 41605
rect 20533 41565 20545 41599
rect 20579 41565 20591 41599
rect 22020 41596 22048 41627
rect 22094 41624 22100 41676
rect 22152 41664 22158 41676
rect 23201 41667 23259 41673
rect 23201 41664 23213 41667
rect 22152 41636 23213 41664
rect 22152 41624 22158 41636
rect 23201 41633 23213 41636
rect 23247 41633 23259 41667
rect 23201 41627 23259 41633
rect 23385 41667 23443 41673
rect 23385 41633 23397 41667
rect 23431 41664 23443 41667
rect 23474 41664 23480 41676
rect 23431 41636 23480 41664
rect 23431 41633 23443 41636
rect 23385 41627 23443 41633
rect 23474 41624 23480 41636
rect 23532 41624 23538 41676
rect 23860 41673 23888 41772
rect 23934 41760 23940 41812
rect 23992 41800 23998 41812
rect 23992 41772 24037 41800
rect 23992 41760 23998 41772
rect 25866 41760 25872 41812
rect 25924 41800 25930 41812
rect 26786 41800 26792 41812
rect 25924 41772 26792 41800
rect 25924 41760 25930 41772
rect 26786 41760 26792 41772
rect 26844 41760 26850 41812
rect 30006 41800 30012 41812
rect 28828 41772 29868 41800
rect 29967 41772 30012 41800
rect 25406 41692 25412 41744
rect 25464 41732 25470 41744
rect 28828 41732 28856 41772
rect 25464 41704 28856 41732
rect 28896 41735 28954 41741
rect 25464 41692 25470 41704
rect 28896 41701 28908 41735
rect 28942 41732 28954 41735
rect 28994 41732 29000 41744
rect 28942 41704 29000 41732
rect 28942 41701 28954 41704
rect 28896 41695 28954 41701
rect 28994 41692 29000 41704
rect 29052 41692 29058 41744
rect 29840 41732 29868 41772
rect 30006 41760 30012 41772
rect 30064 41760 30070 41812
rect 30926 41760 30932 41812
rect 30984 41800 30990 41812
rect 31021 41803 31079 41809
rect 31021 41800 31033 41803
rect 30984 41772 31033 41800
rect 30984 41760 30990 41772
rect 31021 41769 31033 41772
rect 31067 41769 31079 41803
rect 31021 41763 31079 41769
rect 31110 41732 31116 41744
rect 29840 41704 31116 41732
rect 31110 41692 31116 41704
rect 31168 41692 31174 41744
rect 23845 41667 23903 41673
rect 23845 41633 23857 41667
rect 23891 41633 23903 41667
rect 23845 41627 23903 41633
rect 24854 41624 24860 41676
rect 24912 41664 24918 41676
rect 25038 41664 25044 41676
rect 24912 41636 25044 41664
rect 24912 41624 24918 41636
rect 25038 41624 25044 41636
rect 25096 41624 25102 41676
rect 25308 41667 25366 41673
rect 25308 41633 25320 41667
rect 25354 41664 25366 41667
rect 25774 41664 25780 41676
rect 25354 41636 25780 41664
rect 25354 41633 25366 41636
rect 25308 41627 25366 41633
rect 25774 41624 25780 41636
rect 25832 41624 25838 41676
rect 26786 41624 26792 41676
rect 26844 41664 26850 41676
rect 27065 41667 27123 41673
rect 27065 41664 27077 41667
rect 26844 41636 27077 41664
rect 26844 41624 26850 41636
rect 27065 41633 27077 41636
rect 27111 41633 27123 41667
rect 27065 41627 27123 41633
rect 28169 41667 28227 41673
rect 28169 41633 28181 41667
rect 28215 41664 28227 41667
rect 30466 41664 30472 41676
rect 28215 41636 30472 41664
rect 28215 41633 28227 41636
rect 28169 41627 28227 41633
rect 30466 41624 30472 41636
rect 30524 41624 30530 41676
rect 22278 41596 22284 41608
rect 22020 41568 22284 41596
rect 20533 41559 20591 41565
rect 12023 41500 17264 41528
rect 20548 41528 20576 41559
rect 22278 41556 22284 41568
rect 22336 41556 22342 41608
rect 26142 41556 26148 41608
rect 26200 41596 26206 41608
rect 26694 41596 26700 41608
rect 26200 41568 26700 41596
rect 26200 41556 26206 41568
rect 26694 41556 26700 41568
rect 26752 41556 26758 41608
rect 28626 41596 28632 41608
rect 28587 41568 28632 41596
rect 28626 41556 28632 41568
rect 28684 41556 28690 41608
rect 22002 41528 22008 41540
rect 20548 41500 22008 41528
rect 12023 41497 12035 41500
rect 11977 41491 12035 41497
rect 22002 41488 22008 41500
rect 22060 41528 22066 41540
rect 23382 41528 23388 41540
rect 22060 41500 23388 41528
rect 22060 41488 22066 41500
rect 23382 41488 23388 41500
rect 23440 41488 23446 41540
rect 26234 41488 26240 41540
rect 26292 41528 26298 41540
rect 26878 41528 26884 41540
rect 26292 41500 26884 41528
rect 26292 41488 26298 41500
rect 26878 41488 26884 41500
rect 26936 41528 26942 41540
rect 27798 41528 27804 41540
rect 26936 41500 27804 41528
rect 26936 41488 26942 41500
rect 27798 41488 27804 41500
rect 27856 41488 27862 41540
rect 10410 41460 10416 41472
rect 9916 41432 10272 41460
rect 10371 41432 10416 41460
rect 9916 41420 9922 41432
rect 10410 41420 10416 41432
rect 10468 41420 10474 41472
rect 10778 41460 10784 41472
rect 10739 41432 10784 41460
rect 10778 41420 10784 41432
rect 10836 41420 10842 41472
rect 15470 41460 15476 41472
rect 15431 41432 15476 41460
rect 15470 41420 15476 41432
rect 15528 41420 15534 41472
rect 15746 41420 15752 41472
rect 15804 41460 15810 41472
rect 17405 41463 17463 41469
rect 17405 41460 17417 41463
rect 15804 41432 17417 41460
rect 15804 41420 15810 41432
rect 17405 41429 17417 41432
rect 17451 41429 17463 41463
rect 17405 41423 17463 41429
rect 19334 41420 19340 41472
rect 19392 41460 19398 41472
rect 21085 41463 21143 41469
rect 21085 41460 21097 41463
rect 19392 41432 21097 41460
rect 19392 41420 19398 41432
rect 21085 41429 21097 41432
rect 21131 41429 21143 41463
rect 21085 41423 21143 41429
rect 22738 41420 22744 41472
rect 22796 41460 22802 41472
rect 23017 41463 23075 41469
rect 23017 41460 23029 41463
rect 22796 41432 23029 41460
rect 22796 41420 22802 41432
rect 23017 41429 23029 41432
rect 23063 41429 23075 41463
rect 23017 41423 23075 41429
rect 24581 41463 24639 41469
rect 24581 41429 24593 41463
rect 24627 41460 24639 41463
rect 24946 41460 24952 41472
rect 24627 41432 24952 41460
rect 24627 41429 24639 41432
rect 24581 41423 24639 41429
rect 24946 41420 24952 41432
rect 25004 41420 25010 41472
rect 25038 41420 25044 41472
rect 25096 41460 25102 41472
rect 25314 41460 25320 41472
rect 25096 41432 25320 41460
rect 25096 41420 25102 41432
rect 25314 41420 25320 41432
rect 25372 41420 25378 41472
rect 26418 41460 26424 41472
rect 26331 41432 26424 41460
rect 26418 41420 26424 41432
rect 26476 41460 26482 41472
rect 26602 41460 26608 41472
rect 26476 41432 26608 41460
rect 26476 41420 26482 41432
rect 26602 41420 26608 41432
rect 26660 41420 26666 41472
rect 27154 41460 27160 41472
rect 27115 41432 27160 41460
rect 27154 41420 27160 41432
rect 27212 41420 27218 41472
rect 27890 41420 27896 41472
rect 27948 41460 27954 41472
rect 28077 41463 28135 41469
rect 28077 41460 28089 41463
rect 27948 41432 28089 41460
rect 27948 41420 27954 41432
rect 28077 41429 28089 41432
rect 28123 41429 28135 41463
rect 30466 41460 30472 41472
rect 30427 41432 30472 41460
rect 28077 41423 28135 41429
rect 30466 41420 30472 41432
rect 30524 41420 30530 41472
rect 1104 41370 32016 41392
rect 1104 41318 6102 41370
rect 6154 41318 6166 41370
rect 6218 41318 6230 41370
rect 6282 41318 6294 41370
rect 6346 41318 6358 41370
rect 6410 41318 16405 41370
rect 16457 41318 16469 41370
rect 16521 41318 16533 41370
rect 16585 41318 16597 41370
rect 16649 41318 16661 41370
rect 16713 41318 26709 41370
rect 26761 41318 26773 41370
rect 26825 41318 26837 41370
rect 26889 41318 26901 41370
rect 26953 41318 26965 41370
rect 27017 41318 32016 41370
rect 1104 41296 32016 41318
rect 2041 41259 2099 41265
rect 2041 41225 2053 41259
rect 2087 41256 2099 41259
rect 3234 41256 3240 41268
rect 2087 41228 3240 41256
rect 2087 41225 2099 41228
rect 2041 41219 2099 41225
rect 3234 41216 3240 41228
rect 3292 41216 3298 41268
rect 4065 41259 4123 41265
rect 4065 41225 4077 41259
rect 4111 41256 4123 41259
rect 4338 41256 4344 41268
rect 4111 41228 4344 41256
rect 4111 41225 4123 41228
rect 4065 41219 4123 41225
rect 4338 41216 4344 41228
rect 4396 41216 4402 41268
rect 4430 41216 4436 41268
rect 4488 41256 4494 41268
rect 8297 41259 8355 41265
rect 4488 41228 5764 41256
rect 4488 41216 4494 41228
rect 3970 41120 3976 41132
rect 3883 41092 3976 41120
rect 3896 41061 3924 41092
rect 3970 41080 3976 41092
rect 4028 41120 4034 41132
rect 4028 41092 4752 41120
rect 4028 41080 4034 41092
rect 3881 41055 3939 41061
rect 3881 41021 3893 41055
rect 3927 41021 3939 41055
rect 3881 41015 3939 41021
rect 4065 41055 4123 41061
rect 4065 41021 4077 41055
rect 4111 41021 4123 41055
rect 4065 41015 4123 41021
rect 1489 40987 1547 40993
rect 1489 40953 1501 40987
rect 1535 40984 1547 40987
rect 3510 40984 3516 40996
rect 1535 40956 3516 40984
rect 1535 40953 1547 40956
rect 1489 40947 1547 40953
rect 3510 40944 3516 40956
rect 3568 40944 3574 40996
rect 3786 40944 3792 40996
rect 3844 40984 3850 40996
rect 4080 40984 4108 41015
rect 4430 41012 4436 41064
rect 4488 41052 4494 41064
rect 4724 41061 4752 41092
rect 4525 41055 4583 41061
rect 4525 41052 4537 41055
rect 4488 41024 4537 41052
rect 4488 41012 4494 41024
rect 4525 41021 4537 41024
rect 4571 41021 4583 41055
rect 4525 41015 4583 41021
rect 4709 41055 4767 41061
rect 4709 41021 4721 41055
rect 4755 41021 4767 41055
rect 4709 41015 4767 41021
rect 4801 41055 4859 41061
rect 4801 41021 4813 41055
rect 4847 41021 4859 41055
rect 4801 41015 4859 41021
rect 4893 41055 4951 41061
rect 4893 41021 4905 41055
rect 4939 41052 4951 41055
rect 5074 41052 5080 41064
rect 4939 41024 5080 41052
rect 4939 41021 4951 41024
rect 4893 41015 4951 41021
rect 4816 40984 4844 41015
rect 5074 41012 5080 41024
rect 5132 41012 5138 41064
rect 5442 41012 5448 41064
rect 5500 41052 5506 41064
rect 5629 41055 5687 41061
rect 5629 41052 5641 41055
rect 5500 41024 5641 41052
rect 5500 41012 5506 41024
rect 5629 41021 5641 41024
rect 5675 41021 5687 41055
rect 5736 41052 5764 41228
rect 8297 41225 8309 41259
rect 8343 41256 8355 41259
rect 9214 41256 9220 41268
rect 8343 41228 9220 41256
rect 8343 41225 8355 41228
rect 8297 41219 8355 41225
rect 9214 41216 9220 41228
rect 9272 41216 9278 41268
rect 13081 41259 13139 41265
rect 13081 41225 13093 41259
rect 13127 41256 13139 41259
rect 13814 41256 13820 41268
rect 13127 41228 13820 41256
rect 13127 41225 13139 41228
rect 13081 41219 13139 41225
rect 13814 41216 13820 41228
rect 13872 41256 13878 41268
rect 14826 41256 14832 41268
rect 13872 41228 14832 41256
rect 13872 41216 13878 41228
rect 14826 41216 14832 41228
rect 14884 41216 14890 41268
rect 16301 41259 16359 41265
rect 16301 41225 16313 41259
rect 16347 41256 16359 41259
rect 16850 41256 16856 41268
rect 16347 41228 16856 41256
rect 16347 41225 16359 41228
rect 16301 41219 16359 41225
rect 16850 41216 16856 41228
rect 16908 41216 16914 41268
rect 16945 41259 17003 41265
rect 16945 41225 16957 41259
rect 16991 41256 17003 41259
rect 17034 41256 17040 41268
rect 16991 41228 17040 41256
rect 16991 41225 17003 41228
rect 16945 41219 17003 41225
rect 17034 41216 17040 41228
rect 17092 41216 17098 41268
rect 17218 41216 17224 41268
rect 17276 41256 17282 41268
rect 18598 41256 18604 41268
rect 17276 41228 17908 41256
rect 18559 41228 18604 41256
rect 17276 41216 17282 41228
rect 9674 41148 9680 41200
rect 9732 41188 9738 41200
rect 10505 41191 10563 41197
rect 10505 41188 10517 41191
rect 9732 41160 10517 41188
rect 9732 41148 9738 41160
rect 10505 41157 10517 41160
rect 10551 41157 10563 41191
rect 10505 41151 10563 41157
rect 12802 41148 12808 41200
rect 12860 41188 12866 41200
rect 14093 41191 14151 41197
rect 14093 41188 14105 41191
rect 12860 41160 14105 41188
rect 12860 41148 12866 41160
rect 14093 41157 14105 41160
rect 14139 41188 14151 41191
rect 14274 41188 14280 41200
rect 14139 41160 14280 41188
rect 14139 41157 14151 41160
rect 14093 41151 14151 41157
rect 14274 41148 14280 41160
rect 14332 41148 14338 41200
rect 17770 41188 17776 41200
rect 17731 41160 17776 41188
rect 17770 41148 17776 41160
rect 17828 41148 17834 41200
rect 17880 41188 17908 41228
rect 18598 41216 18604 41228
rect 18656 41216 18662 41268
rect 19242 41256 19248 41268
rect 19203 41228 19248 41256
rect 19242 41216 19248 41228
rect 19300 41216 19306 41268
rect 20990 41256 20996 41268
rect 19628 41228 20996 41256
rect 19518 41188 19524 41200
rect 17880 41160 19524 41188
rect 19518 41148 19524 41160
rect 19576 41148 19582 41200
rect 8294 41080 8300 41132
rect 8352 41120 8358 41132
rect 11054 41120 11060 41132
rect 8352 41092 11060 41120
rect 8352 41080 8358 41092
rect 11054 41080 11060 41092
rect 11112 41120 11118 41132
rect 11606 41120 11612 41132
rect 11112 41092 11612 41120
rect 11112 41080 11118 41092
rect 11606 41080 11612 41092
rect 11664 41120 11670 41132
rect 11701 41123 11759 41129
rect 11701 41120 11713 41123
rect 11664 41092 11713 41120
rect 11664 41080 11670 41092
rect 11701 41089 11713 41092
rect 11747 41089 11759 41123
rect 11701 41083 11759 41089
rect 16114 41080 16120 41132
rect 16172 41120 16178 41132
rect 16850 41120 16856 41132
rect 16172 41092 16856 41120
rect 16172 41080 16178 41092
rect 16850 41080 16856 41092
rect 16908 41120 16914 41132
rect 16908 41092 18184 41120
rect 16908 41080 16914 41092
rect 5813 41055 5871 41061
rect 5813 41052 5825 41055
rect 5736 41024 5825 41052
rect 5629 41015 5687 41021
rect 5813 41021 5825 41024
rect 5859 41021 5871 41055
rect 5813 41015 5871 41021
rect 8205 41055 8263 41061
rect 8205 41021 8217 41055
rect 8251 41052 8263 41055
rect 8478 41052 8484 41064
rect 8251 41024 8484 41052
rect 8251 41021 8263 41024
rect 8205 41015 8263 41021
rect 8478 41012 8484 41024
rect 8536 41052 8542 41064
rect 8846 41052 8852 41064
rect 8536 41024 8852 41052
rect 8536 41012 8542 41024
rect 8846 41012 8852 41024
rect 8904 41012 8910 41064
rect 8941 41055 8999 41061
rect 8941 41021 8953 41055
rect 8987 41021 8999 41055
rect 8941 41015 8999 41021
rect 9217 41055 9275 41061
rect 9217 41021 9229 41055
rect 9263 41052 9275 41055
rect 9306 41052 9312 41064
rect 9263 41024 9312 41052
rect 9263 41021 9275 41024
rect 9217 41015 9275 41021
rect 3844 40956 4108 40984
rect 4172 40956 4844 40984
rect 5169 40987 5227 40993
rect 3844 40944 3850 40956
rect 2498 40916 2504 40928
rect 2459 40888 2504 40916
rect 2498 40876 2504 40888
rect 2556 40876 2562 40928
rect 3237 40919 3295 40925
rect 3237 40885 3249 40919
rect 3283 40916 3295 40919
rect 3602 40916 3608 40928
rect 3283 40888 3608 40916
rect 3283 40885 3295 40888
rect 3237 40879 3295 40885
rect 3602 40876 3608 40888
rect 3660 40916 3666 40928
rect 4172 40916 4200 40956
rect 5169 40953 5181 40987
rect 5215 40984 5227 40987
rect 5902 40984 5908 40996
rect 5215 40956 5908 40984
rect 5215 40953 5227 40956
rect 5169 40947 5227 40953
rect 5902 40944 5908 40956
rect 5960 40944 5966 40996
rect 7745 40987 7803 40993
rect 7745 40953 7757 40987
rect 7791 40984 7803 40987
rect 7834 40984 7840 40996
rect 7791 40956 7840 40984
rect 7791 40953 7803 40956
rect 7745 40947 7803 40953
rect 7834 40944 7840 40956
rect 7892 40984 7898 40996
rect 8570 40984 8576 40996
rect 7892 40956 8576 40984
rect 7892 40944 7898 40956
rect 8570 40944 8576 40956
rect 8628 40984 8634 40996
rect 8956 40984 8984 41015
rect 9306 41012 9312 41024
rect 9364 41012 9370 41064
rect 10226 41052 10232 41064
rect 10187 41024 10232 41052
rect 10226 41012 10232 41024
rect 10284 41012 10290 41064
rect 10410 41052 10416 41064
rect 10371 41024 10416 41052
rect 10410 41012 10416 41024
rect 10468 41012 10474 41064
rect 10594 41052 10600 41064
rect 10555 41024 10600 41052
rect 10594 41012 10600 41024
rect 10652 41012 10658 41064
rect 10686 41012 10692 41064
rect 10744 41052 10750 41064
rect 10744 41024 10789 41052
rect 10744 41012 10750 41024
rect 13078 41012 13084 41064
rect 13136 41052 13142 41064
rect 15470 41052 15476 41064
rect 13136 41024 15476 41052
rect 13136 41012 13142 41024
rect 15470 41012 15476 41024
rect 15528 41012 15534 41064
rect 15933 41055 15991 41061
rect 15933 41021 15945 41055
rect 15979 41021 15991 41055
rect 15933 41015 15991 41021
rect 16301 41055 16359 41061
rect 16301 41021 16313 41055
rect 16347 41052 16359 41055
rect 16942 41052 16948 41064
rect 16347 41024 16948 41052
rect 16347 41021 16359 41024
rect 16301 41015 16359 41021
rect 8628 40956 8984 40984
rect 8628 40944 8634 40956
rect 10134 40944 10140 40996
rect 10192 40984 10198 40996
rect 10612 40984 10640 41012
rect 10192 40956 10640 40984
rect 11968 40987 12026 40993
rect 10192 40944 10198 40956
rect 11968 40953 11980 40987
rect 12014 40984 12026 40987
rect 12250 40984 12256 40996
rect 12014 40956 12256 40984
rect 12014 40953 12026 40956
rect 11968 40947 12026 40953
rect 12250 40944 12256 40956
rect 12308 40944 12314 40996
rect 14366 40944 14372 40996
rect 14424 40984 14430 40996
rect 15206 40987 15264 40993
rect 15206 40984 15218 40987
rect 14424 40956 15218 40984
rect 14424 40944 14430 40956
rect 15206 40953 15218 40956
rect 15252 40953 15264 40987
rect 15206 40947 15264 40953
rect 5718 40916 5724 40928
rect 3660 40888 4200 40916
rect 5679 40888 5724 40916
rect 3660 40876 3666 40888
rect 5718 40876 5724 40888
rect 5776 40876 5782 40928
rect 6641 40919 6699 40925
rect 6641 40885 6653 40919
rect 6687 40916 6699 40919
rect 6822 40916 6828 40928
rect 6687 40888 6828 40916
rect 6687 40885 6699 40888
rect 6641 40879 6699 40885
rect 6822 40876 6828 40888
rect 6880 40876 6886 40928
rect 7098 40916 7104 40928
rect 7059 40888 7104 40916
rect 7098 40876 7104 40888
rect 7156 40876 7162 40928
rect 10870 40916 10876 40928
rect 10831 40888 10876 40916
rect 10870 40876 10876 40888
rect 10928 40876 10934 40928
rect 14734 40876 14740 40928
rect 14792 40916 14798 40928
rect 15948 40916 15976 41015
rect 16942 41012 16948 41024
rect 17000 41012 17006 41064
rect 17129 41055 17187 41061
rect 17129 41021 17141 41055
rect 17175 41052 17187 41055
rect 17218 41052 17224 41064
rect 17175 41024 17224 41052
rect 17175 41021 17187 41024
rect 17129 41015 17187 41021
rect 17218 41012 17224 41024
rect 17276 41012 17282 41064
rect 17310 40984 17316 40996
rect 17223 40956 17316 40984
rect 17310 40944 17316 40956
rect 17368 40984 17374 40996
rect 17678 40984 17684 40996
rect 17368 40956 17684 40984
rect 17368 40944 17374 40956
rect 17678 40944 17684 40956
rect 17736 40944 17742 40996
rect 17954 40984 17960 40996
rect 17867 40956 17960 40984
rect 17954 40944 17960 40956
rect 18012 40944 18018 40996
rect 18156 40993 18184 41092
rect 19242 41080 19248 41132
rect 19300 41120 19306 41132
rect 19300 41092 19564 41120
rect 19300 41080 19306 41092
rect 19426 41052 19432 41064
rect 19387 41024 19432 41052
rect 19426 41012 19432 41024
rect 19484 41012 19490 41064
rect 18141 40987 18199 40993
rect 18141 40953 18153 40987
rect 18187 40984 18199 40987
rect 19334 40984 19340 40996
rect 18187 40956 19340 40984
rect 18187 40953 18199 40956
rect 18141 40947 18199 40953
rect 19334 40944 19340 40956
rect 19392 40944 19398 40996
rect 19536 40984 19564 41092
rect 19628 41061 19656 41228
rect 20990 41216 20996 41228
rect 21048 41216 21054 41268
rect 21266 41216 21272 41268
rect 21324 41256 21330 41268
rect 22557 41259 22615 41265
rect 22557 41256 22569 41259
rect 21324 41228 22569 41256
rect 21324 41216 21330 41228
rect 22557 41225 22569 41228
rect 22603 41225 22615 41259
rect 22557 41219 22615 41225
rect 23293 41259 23351 41265
rect 23293 41225 23305 41259
rect 23339 41256 23351 41259
rect 23474 41256 23480 41268
rect 23339 41228 23480 41256
rect 23339 41225 23351 41228
rect 23293 41219 23351 41225
rect 20438 41188 20444 41200
rect 19720 41160 20444 41188
rect 19720 41129 19748 41160
rect 20438 41148 20444 41160
rect 20496 41148 20502 41200
rect 21082 41188 21088 41200
rect 20824 41160 21088 41188
rect 19696 41123 19754 41129
rect 19696 41089 19708 41123
rect 19742 41089 19754 41123
rect 19696 41083 19754 41089
rect 20070 41080 20076 41132
rect 20128 41120 20134 41132
rect 20824 41129 20852 41160
rect 21082 41148 21088 41160
rect 21140 41148 21146 41200
rect 22572 41188 22600 41219
rect 23474 41216 23480 41228
rect 23532 41256 23538 41268
rect 24302 41256 24308 41268
rect 23532 41228 24308 41256
rect 23532 41216 23538 41228
rect 24302 41216 24308 41228
rect 24360 41216 24366 41268
rect 25774 41256 25780 41268
rect 25735 41228 25780 41256
rect 25774 41216 25780 41228
rect 25832 41216 25838 41268
rect 24578 41188 24584 41200
rect 22572 41160 24584 41188
rect 24578 41148 24584 41160
rect 24636 41148 24642 41200
rect 26326 41148 26332 41200
rect 26384 41188 26390 41200
rect 26384 41160 26556 41188
rect 26384 41148 26390 41160
rect 20809 41123 20867 41129
rect 20809 41120 20821 41123
rect 20128 41092 20821 41120
rect 20128 41080 20134 41092
rect 20809 41089 20821 41092
rect 20855 41089 20867 41123
rect 20809 41083 20867 41089
rect 23014 41080 23020 41132
rect 23072 41120 23078 41132
rect 23201 41123 23259 41129
rect 23201 41120 23213 41123
rect 23072 41092 23213 41120
rect 23072 41080 23078 41092
rect 23201 41089 23213 41092
rect 23247 41089 23259 41123
rect 25130 41120 25136 41132
rect 23201 41083 23259 41089
rect 24412 41092 25136 41120
rect 19613 41055 19671 41061
rect 19613 41021 19625 41055
rect 19659 41021 19671 41055
rect 19613 41015 19671 41021
rect 19797 41055 19855 41061
rect 19797 41021 19809 41055
rect 19843 41021 19855 41055
rect 19797 41015 19855 41021
rect 19981 41055 20039 41061
rect 19981 41021 19993 41055
rect 20027 41052 20039 41055
rect 20346 41052 20352 41064
rect 20027 41024 20352 41052
rect 20027 41021 20039 41024
rect 19981 41015 20039 41021
rect 19812 40984 19840 41015
rect 20346 41012 20352 41024
rect 20404 41012 20410 41064
rect 20438 41012 20444 41064
rect 20496 41052 20502 41064
rect 21085 41055 21143 41061
rect 21085 41052 21097 41055
rect 20496 41024 21097 41052
rect 20496 41012 20502 41024
rect 21085 41021 21097 41024
rect 21131 41021 21143 41055
rect 21085 41015 21143 41021
rect 22278 41012 22284 41064
rect 22336 41052 22342 41064
rect 22373 41055 22431 41061
rect 22373 41052 22385 41055
rect 22336 41024 22385 41052
rect 22336 41012 22342 41024
rect 22373 41021 22385 41024
rect 22419 41052 22431 41055
rect 22462 41052 22468 41064
rect 22419 41024 22468 41052
rect 22419 41021 22431 41024
rect 22373 41015 22431 41021
rect 22462 41012 22468 41024
rect 22520 41012 22526 41064
rect 22649 41055 22707 41061
rect 22649 41021 22661 41055
rect 22695 41021 22707 41055
rect 23106 41052 23112 41064
rect 23067 41024 23112 41052
rect 22649 41015 22707 41021
rect 22664 40984 22692 41015
rect 23106 41012 23112 41024
rect 23164 41012 23170 41064
rect 23474 41012 23480 41064
rect 23532 41052 23538 41064
rect 24412 41061 24440 41092
rect 25130 41080 25136 41092
rect 25188 41080 25194 41132
rect 26142 41120 26148 41132
rect 26103 41092 26148 41120
rect 26142 41080 26148 41092
rect 26200 41080 26206 41132
rect 24397 41055 24455 41061
rect 24397 41052 24409 41055
rect 23532 41024 24409 41052
rect 23532 41012 23538 41024
rect 24397 41021 24409 41024
rect 24443 41021 24455 41055
rect 24397 41015 24455 41021
rect 24673 41055 24731 41061
rect 24673 41021 24685 41055
rect 24719 41021 24731 41055
rect 24673 41015 24731 41021
rect 25961 41055 26019 41061
rect 25961 41021 25973 41055
rect 26007 41021 26019 41055
rect 26234 41052 26240 41064
rect 26195 41024 26240 41052
rect 25961 41015 26019 41021
rect 19536 40956 22692 40984
rect 24210 40944 24216 40996
rect 24268 40984 24274 40996
rect 24688 40984 24716 41015
rect 24268 40956 24716 40984
rect 25976 40984 26004 41015
rect 26234 41012 26240 41024
rect 26292 41012 26298 41064
rect 26326 41012 26332 41064
rect 26384 41052 26390 41064
rect 26528 41061 26556 41160
rect 28626 41120 28632 41132
rect 28587 41092 28632 41120
rect 28626 41080 28632 41092
rect 28684 41120 28690 41132
rect 29641 41123 29699 41129
rect 29641 41120 29653 41123
rect 28684 41092 29653 41120
rect 28684 41080 28690 41092
rect 29641 41089 29653 41092
rect 29687 41089 29699 41123
rect 29641 41083 29699 41089
rect 26513 41055 26571 41061
rect 26384 41024 26429 41052
rect 26384 41012 26390 41024
rect 26513 41021 26525 41055
rect 26559 41021 26571 41055
rect 26513 41015 26571 41021
rect 26973 41055 27031 41061
rect 26973 41021 26985 41055
rect 27019 41052 27031 41055
rect 27062 41052 27068 41064
rect 27019 41024 27068 41052
rect 27019 41021 27031 41024
rect 26973 41015 27031 41021
rect 27062 41012 27068 41024
rect 27120 41012 27126 41064
rect 29908 41055 29966 41061
rect 29908 41021 29920 41055
rect 29954 41052 29966 41055
rect 30282 41052 30288 41064
rect 29954 41024 30288 41052
rect 29954 41021 29966 41024
rect 29908 41015 29966 41021
rect 30282 41012 30288 41024
rect 30340 41012 30346 41064
rect 26602 40984 26608 40996
rect 25976 40956 26608 40984
rect 24268 40944 24274 40956
rect 26602 40944 26608 40956
rect 26660 40944 26666 40996
rect 14792 40888 15976 40916
rect 14792 40876 14798 40888
rect 16206 40876 16212 40928
rect 16264 40916 16270 40928
rect 16485 40919 16543 40925
rect 16485 40916 16497 40919
rect 16264 40888 16497 40916
rect 16264 40876 16270 40888
rect 16485 40885 16497 40888
rect 16531 40885 16543 40919
rect 16485 40879 16543 40885
rect 16942 40876 16948 40928
rect 17000 40916 17006 40928
rect 17972 40916 18000 40944
rect 17000 40888 18000 40916
rect 17000 40876 17006 40888
rect 18598 40876 18604 40928
rect 18656 40916 18662 40928
rect 19702 40916 19708 40928
rect 18656 40888 19708 40916
rect 18656 40876 18662 40888
rect 19702 40876 19708 40888
rect 19760 40876 19766 40928
rect 21910 40876 21916 40928
rect 21968 40916 21974 40928
rect 22097 40919 22155 40925
rect 22097 40916 22109 40919
rect 21968 40888 22109 40916
rect 21968 40876 21974 40888
rect 22097 40885 22109 40888
rect 22143 40885 22155 40919
rect 22097 40879 22155 40885
rect 22278 40876 22284 40928
rect 22336 40916 22342 40928
rect 23477 40919 23535 40925
rect 23477 40916 23489 40919
rect 22336 40888 23489 40916
rect 22336 40876 22342 40888
rect 23477 40885 23489 40888
rect 23523 40885 23535 40919
rect 23477 40879 23535 40885
rect 30558 40876 30564 40928
rect 30616 40916 30622 40928
rect 31018 40916 31024 40928
rect 30616 40888 31024 40916
rect 30616 40876 30622 40888
rect 31018 40876 31024 40888
rect 31076 40876 31082 40928
rect 1104 40826 32016 40848
rect 1104 40774 11253 40826
rect 11305 40774 11317 40826
rect 11369 40774 11381 40826
rect 11433 40774 11445 40826
rect 11497 40774 11509 40826
rect 11561 40774 21557 40826
rect 21609 40774 21621 40826
rect 21673 40774 21685 40826
rect 21737 40774 21749 40826
rect 21801 40774 21813 40826
rect 21865 40774 32016 40826
rect 1104 40752 32016 40774
rect 2866 40712 2872 40724
rect 1872 40684 2872 40712
rect 1394 40536 1400 40588
rect 1452 40576 1458 40588
rect 1872 40585 1900 40684
rect 2866 40672 2872 40684
rect 2924 40672 2930 40724
rect 3970 40672 3976 40724
rect 4028 40712 4034 40724
rect 4065 40715 4123 40721
rect 4065 40712 4077 40715
rect 4028 40684 4077 40712
rect 4028 40672 4034 40684
rect 4065 40681 4077 40684
rect 4111 40681 4123 40715
rect 4065 40675 4123 40681
rect 7837 40715 7895 40721
rect 7837 40681 7849 40715
rect 7883 40712 7895 40715
rect 8478 40712 8484 40724
rect 7883 40684 8484 40712
rect 7883 40681 7895 40684
rect 7837 40675 7895 40681
rect 8478 40672 8484 40684
rect 8536 40672 8542 40724
rect 10226 40672 10232 40724
rect 10284 40712 10290 40724
rect 10781 40715 10839 40721
rect 10781 40712 10793 40715
rect 10284 40684 10793 40712
rect 10284 40672 10290 40684
rect 10781 40681 10793 40684
rect 10827 40681 10839 40715
rect 12250 40712 12256 40724
rect 12211 40684 12256 40712
rect 10781 40675 10839 40681
rect 12250 40672 12256 40684
rect 12308 40672 12314 40724
rect 13814 40712 13820 40724
rect 12452 40684 13820 40712
rect 2774 40644 2780 40656
rect 2700 40616 2780 40644
rect 1857 40579 1915 40585
rect 1857 40576 1869 40579
rect 1452 40548 1869 40576
rect 1452 40536 1458 40548
rect 1857 40545 1869 40548
rect 1903 40545 1915 40579
rect 1857 40539 1915 40545
rect 2700 40517 2728 40616
rect 2774 40604 2780 40616
rect 2832 40644 2838 40656
rect 3694 40644 3700 40656
rect 2832 40616 3700 40644
rect 2832 40604 2838 40616
rect 3694 40604 3700 40616
rect 3752 40604 3758 40656
rect 5442 40644 5448 40656
rect 4724 40616 5448 40644
rect 2952 40579 3010 40585
rect 2952 40545 2964 40579
rect 2998 40576 3010 40579
rect 3234 40576 3240 40588
rect 2998 40548 3240 40576
rect 2998 40545 3010 40548
rect 2952 40539 3010 40545
rect 3234 40536 3240 40548
rect 3292 40536 3298 40588
rect 3326 40536 3332 40588
rect 3384 40576 3390 40588
rect 3786 40576 3792 40588
rect 3384 40548 3792 40576
rect 3384 40536 3390 40548
rect 3786 40536 3792 40548
rect 3844 40576 3850 40588
rect 4724 40585 4752 40616
rect 5442 40604 5448 40616
rect 5500 40604 5506 40656
rect 8294 40644 8300 40656
rect 6472 40616 8300 40644
rect 4525 40579 4583 40585
rect 4525 40576 4537 40579
rect 3844 40548 4537 40576
rect 3844 40536 3850 40548
rect 4525 40545 4537 40548
rect 4571 40545 4583 40579
rect 4525 40539 4583 40545
rect 4709 40579 4767 40585
rect 4709 40545 4721 40579
rect 4755 40545 4767 40579
rect 4709 40539 4767 40545
rect 2685 40511 2743 40517
rect 2685 40477 2697 40511
rect 2731 40477 2743 40511
rect 2685 40471 2743 40477
rect 4062 40468 4068 40520
rect 4120 40508 4126 40520
rect 4724 40508 4752 40539
rect 4798 40536 4804 40588
rect 4856 40576 4862 40588
rect 4939 40579 4997 40585
rect 4856 40548 4901 40576
rect 4856 40536 4862 40548
rect 4939 40545 4951 40579
rect 4985 40576 4997 40579
rect 5074 40576 5080 40588
rect 4985 40548 5080 40576
rect 4985 40545 4997 40548
rect 4939 40539 4997 40545
rect 5074 40536 5080 40548
rect 5132 40536 5138 40588
rect 5626 40536 5632 40588
rect 5684 40576 5690 40588
rect 6472 40585 6500 40616
rect 8294 40604 8300 40616
rect 8352 40604 8358 40656
rect 8662 40604 8668 40656
rect 8720 40644 8726 40656
rect 8720 40616 8800 40644
rect 8720 40604 8726 40616
rect 5813 40579 5871 40585
rect 5813 40576 5825 40579
rect 5684 40548 5825 40576
rect 5684 40536 5690 40548
rect 5813 40545 5825 40548
rect 5859 40545 5871 40579
rect 5813 40539 5871 40545
rect 6457 40579 6515 40585
rect 6457 40545 6469 40579
rect 6503 40545 6515 40579
rect 6457 40539 6515 40545
rect 6724 40579 6782 40585
rect 6724 40545 6736 40579
rect 6770 40576 6782 40579
rect 8478 40576 8484 40588
rect 6770 40548 8340 40576
rect 8439 40548 8484 40576
rect 6770 40545 6782 40548
rect 6724 40539 6782 40545
rect 8312 40517 8340 40548
rect 8478 40536 8484 40548
rect 8536 40536 8542 40588
rect 8772 40585 8800 40616
rect 10318 40604 10324 40656
rect 10376 40644 10382 40656
rect 10376 40616 10640 40644
rect 10376 40604 10382 40616
rect 8757 40579 8815 40585
rect 8757 40545 8769 40579
rect 8803 40545 8815 40579
rect 8757 40539 8815 40545
rect 8849 40579 8907 40585
rect 8849 40545 8861 40579
rect 8895 40576 8907 40579
rect 8938 40576 8944 40588
rect 8895 40548 8944 40576
rect 8895 40545 8907 40548
rect 8849 40539 8907 40545
rect 8938 40536 8944 40548
rect 8996 40536 9002 40588
rect 9033 40579 9091 40585
rect 9033 40545 9045 40579
rect 9079 40576 9091 40579
rect 9306 40576 9312 40588
rect 9079 40548 9312 40576
rect 9079 40545 9091 40548
rect 9033 40539 9091 40545
rect 9306 40536 9312 40548
rect 9364 40536 9370 40588
rect 9493 40579 9551 40585
rect 9493 40545 9505 40579
rect 9539 40545 9551 40579
rect 9493 40539 9551 40545
rect 9677 40579 9735 40585
rect 9677 40545 9689 40579
rect 9723 40576 9735 40579
rect 10134 40576 10140 40588
rect 9723 40548 10140 40576
rect 9723 40545 9735 40548
rect 9677 40539 9735 40545
rect 4120 40480 4752 40508
rect 8297 40511 8355 40517
rect 4120 40468 4126 40480
rect 8297 40477 8309 40511
rect 8343 40477 8355 40511
rect 8297 40471 8355 40477
rect 8665 40511 8723 40517
rect 8665 40477 8677 40511
rect 8711 40508 8723 40511
rect 9508 40508 9536 40539
rect 10134 40536 10140 40548
rect 10192 40536 10198 40588
rect 10612 40585 10640 40616
rect 12452 40585 12480 40684
rect 13814 40672 13820 40684
rect 13872 40672 13878 40724
rect 14734 40672 14740 40724
rect 14792 40712 14798 40724
rect 14829 40715 14887 40721
rect 14829 40712 14841 40715
rect 14792 40684 14841 40712
rect 14792 40672 14798 40684
rect 14829 40681 14841 40684
rect 14875 40681 14887 40715
rect 17218 40712 17224 40724
rect 14829 40675 14887 40681
rect 15948 40684 17224 40712
rect 13722 40653 13728 40656
rect 13716 40644 13728 40653
rect 13683 40616 13728 40644
rect 13716 40607 13728 40616
rect 13722 40604 13728 40607
rect 13780 40604 13786 40656
rect 15948 40653 15976 40684
rect 17218 40672 17224 40684
rect 17276 40672 17282 40724
rect 17402 40672 17408 40724
rect 17460 40672 17466 40724
rect 19242 40672 19248 40724
rect 19300 40712 19306 40724
rect 20717 40715 20775 40721
rect 20717 40712 20729 40715
rect 19300 40684 20729 40712
rect 19300 40672 19306 40684
rect 20717 40681 20729 40684
rect 20763 40681 20775 40715
rect 20717 40675 20775 40681
rect 21174 40672 21180 40724
rect 21232 40712 21238 40724
rect 21232 40684 22416 40712
rect 21232 40672 21238 40684
rect 15933 40647 15991 40653
rect 15933 40613 15945 40647
rect 15979 40613 15991 40647
rect 16114 40644 16120 40656
rect 16075 40616 16120 40644
rect 15933 40607 15991 40613
rect 16114 40604 16120 40616
rect 16172 40604 16178 40656
rect 17126 40604 17132 40656
rect 17184 40604 17190 40656
rect 17420 40644 17448 40672
rect 17236 40616 17448 40644
rect 10597 40579 10655 40585
rect 10597 40545 10609 40579
rect 10643 40576 10655 40579
rect 11701 40579 11759 40585
rect 11701 40576 11713 40579
rect 10643 40548 11713 40576
rect 10643 40545 10655 40548
rect 10597 40539 10655 40545
rect 11701 40545 11713 40548
rect 11747 40576 11759 40579
rect 12437 40579 12495 40585
rect 11747 40548 12112 40576
rect 11747 40545 11759 40548
rect 11701 40539 11759 40545
rect 9858 40508 9864 40520
rect 8711 40480 8892 40508
rect 9508 40480 9864 40508
rect 8711 40477 8723 40480
rect 8665 40471 8723 40477
rect 8864 40452 8892 40480
rect 9858 40468 9864 40480
rect 9916 40468 9922 40520
rect 10318 40508 10324 40520
rect 10279 40480 10324 40508
rect 10318 40468 10324 40480
rect 10376 40468 10382 40520
rect 10413 40511 10471 40517
rect 10413 40477 10425 40511
rect 10459 40508 10471 40511
rect 10962 40508 10968 40520
rect 10459 40480 10968 40508
rect 10459 40477 10471 40480
rect 10413 40471 10471 40477
rect 10962 40468 10968 40480
rect 11020 40468 11026 40520
rect 12084 40452 12112 40548
rect 12437 40545 12449 40579
rect 12483 40545 12495 40579
rect 12802 40576 12808 40588
rect 12763 40548 12808 40576
rect 12437 40539 12495 40545
rect 12802 40536 12808 40548
rect 12860 40536 12866 40588
rect 12986 40536 12992 40588
rect 13044 40576 13050 40588
rect 13538 40576 13544 40588
rect 13044 40548 13544 40576
rect 13044 40536 13050 40548
rect 13538 40536 13544 40548
rect 13596 40536 13602 40588
rect 16850 40576 16856 40588
rect 16811 40548 16856 40576
rect 16850 40536 16856 40548
rect 16908 40536 16914 40588
rect 17037 40579 17095 40585
rect 17037 40545 17049 40579
rect 17083 40576 17095 40579
rect 17144 40576 17172 40604
rect 17236 40585 17264 40616
rect 18046 40604 18052 40656
rect 18104 40644 18110 40656
rect 19582 40647 19640 40653
rect 19582 40644 19594 40647
rect 18104 40616 19594 40644
rect 18104 40604 18110 40616
rect 19582 40613 19594 40616
rect 19628 40613 19640 40647
rect 19582 40607 19640 40613
rect 21821 40647 21879 40653
rect 21821 40613 21833 40647
rect 21867 40644 21879 40647
rect 22094 40644 22100 40656
rect 21867 40616 22100 40644
rect 21867 40613 21879 40616
rect 21821 40607 21879 40613
rect 22094 40604 22100 40616
rect 22152 40604 22158 40656
rect 22388 40644 22416 40684
rect 22462 40672 22468 40724
rect 22520 40712 22526 40724
rect 22646 40712 22652 40724
rect 22520 40684 22652 40712
rect 22520 40672 22526 40684
rect 22646 40672 22652 40684
rect 22704 40672 22710 40724
rect 26329 40715 26387 40721
rect 26329 40681 26341 40715
rect 26375 40712 26387 40715
rect 27246 40712 27252 40724
rect 26375 40684 27252 40712
rect 26375 40681 26387 40684
rect 26329 40675 26387 40681
rect 27246 40672 27252 40684
rect 27304 40672 27310 40724
rect 23474 40644 23480 40656
rect 22388 40616 23480 40644
rect 23474 40604 23480 40616
rect 23532 40604 23538 40656
rect 24210 40604 24216 40656
rect 24268 40644 24274 40656
rect 24268 40616 24440 40644
rect 24268 40604 24274 40616
rect 17083 40548 17172 40576
rect 17221 40579 17279 40585
rect 17083 40545 17095 40548
rect 17037 40539 17095 40545
rect 17221 40545 17233 40579
rect 17267 40545 17279 40579
rect 17221 40539 17279 40545
rect 17310 40536 17316 40588
rect 17368 40576 17374 40588
rect 17405 40579 17463 40585
rect 17405 40576 17417 40579
rect 17368 40548 17417 40576
rect 17368 40536 17374 40548
rect 17405 40545 17417 40548
rect 17451 40545 17463 40579
rect 17405 40539 17463 40545
rect 18506 40536 18512 40588
rect 18564 40576 18570 40588
rect 19337 40579 19395 40585
rect 19337 40576 19349 40579
rect 18564 40548 19349 40576
rect 18564 40536 18570 40548
rect 19337 40545 19349 40548
rect 19383 40576 19395 40579
rect 19426 40576 19432 40588
rect 19383 40548 19432 40576
rect 19383 40545 19395 40548
rect 19337 40539 19395 40545
rect 19426 40536 19432 40548
rect 19484 40536 19490 40588
rect 22002 40576 22008 40588
rect 21963 40548 22008 40576
rect 22002 40536 22008 40548
rect 22060 40536 22066 40588
rect 22186 40576 22192 40588
rect 22147 40548 22192 40576
rect 22186 40536 22192 40548
rect 22244 40536 22250 40588
rect 22278 40536 22284 40588
rect 22336 40576 22342 40588
rect 22336 40548 22381 40576
rect 22336 40536 22342 40548
rect 22462 40536 22468 40588
rect 22520 40576 22526 40588
rect 22520 40548 22565 40576
rect 22520 40536 22526 40548
rect 23106 40536 23112 40588
rect 23164 40576 23170 40588
rect 24314 40579 24372 40585
rect 24314 40576 24326 40579
rect 23164 40548 24326 40576
rect 23164 40536 23170 40548
rect 24314 40545 24326 40548
rect 24360 40545 24372 40579
rect 24412 40576 24440 40616
rect 26050 40604 26056 40656
rect 26108 40644 26114 40656
rect 27338 40644 27344 40656
rect 26108 40616 26280 40644
rect 26108 40604 26114 40616
rect 25041 40579 25099 40585
rect 25041 40576 25053 40579
rect 24412 40548 25053 40576
rect 24314 40539 24372 40545
rect 25041 40545 25053 40548
rect 25087 40545 25099 40579
rect 25225 40579 25283 40585
rect 25225 40576 25237 40579
rect 25041 40539 25099 40545
rect 25148 40548 25237 40576
rect 12618 40508 12624 40520
rect 12579 40480 12624 40508
rect 12618 40468 12624 40480
rect 12676 40468 12682 40520
rect 12713 40511 12771 40517
rect 12713 40477 12725 40511
rect 12759 40477 12771 40511
rect 12713 40471 12771 40477
rect 8846 40400 8852 40452
rect 8904 40400 8910 40452
rect 10505 40443 10563 40449
rect 10505 40409 10517 40443
rect 10551 40409 10563 40443
rect 10505 40403 10563 40409
rect 1946 40372 1952 40384
rect 1907 40344 1952 40372
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 5169 40375 5227 40381
rect 5169 40341 5181 40375
rect 5215 40372 5227 40375
rect 5258 40372 5264 40384
rect 5215 40344 5264 40372
rect 5215 40341 5227 40344
rect 5169 40335 5227 40341
rect 5258 40332 5264 40344
rect 5316 40332 5322 40384
rect 5534 40332 5540 40384
rect 5592 40372 5598 40384
rect 5721 40375 5779 40381
rect 5721 40372 5733 40375
rect 5592 40344 5733 40372
rect 5592 40332 5598 40344
rect 5721 40341 5733 40344
rect 5767 40341 5779 40375
rect 5721 40335 5779 40341
rect 9677 40375 9735 40381
rect 9677 40341 9689 40375
rect 9723 40372 9735 40375
rect 10226 40372 10232 40384
rect 9723 40344 10232 40372
rect 9723 40341 9735 40344
rect 9677 40335 9735 40341
rect 10226 40332 10232 40344
rect 10284 40332 10290 40384
rect 10520 40372 10548 40403
rect 10686 40400 10692 40452
rect 10744 40440 10750 40452
rect 11609 40443 11667 40449
rect 11609 40440 11621 40443
rect 10744 40412 11621 40440
rect 10744 40400 10750 40412
rect 11609 40409 11621 40412
rect 11655 40409 11667 40443
rect 11609 40403 11667 40409
rect 12066 40400 12072 40452
rect 12124 40440 12130 40452
rect 12526 40440 12532 40452
rect 12124 40412 12532 40440
rect 12124 40400 12130 40412
rect 12526 40400 12532 40412
rect 12584 40400 12590 40452
rect 10594 40372 10600 40384
rect 10507 40344 10600 40372
rect 10594 40332 10600 40344
rect 10652 40372 10658 40384
rect 11422 40372 11428 40384
rect 10652 40344 11428 40372
rect 10652 40332 10658 40344
rect 11422 40332 11428 40344
rect 11480 40332 11486 40384
rect 12728 40372 12756 40471
rect 13078 40468 13084 40520
rect 13136 40508 13142 40520
rect 13449 40511 13507 40517
rect 13449 40508 13461 40511
rect 13136 40480 13461 40508
rect 13136 40468 13142 40480
rect 13449 40477 13461 40480
rect 13495 40477 13507 40511
rect 13449 40471 13507 40477
rect 17129 40511 17187 40517
rect 17129 40477 17141 40511
rect 17175 40508 17187 40511
rect 17770 40508 17776 40520
rect 17175 40480 17776 40508
rect 17175 40477 17187 40480
rect 17129 40471 17187 40477
rect 17770 40468 17776 40480
rect 17828 40508 17834 40520
rect 18601 40511 18659 40517
rect 18601 40508 18613 40511
rect 17828 40480 18613 40508
rect 17828 40468 17834 40480
rect 18601 40477 18613 40480
rect 18647 40477 18659 40511
rect 18601 40471 18659 40477
rect 18877 40511 18935 40517
rect 18877 40477 18889 40511
rect 18923 40508 18935 40511
rect 22097 40511 22155 40517
rect 18923 40480 19380 40508
rect 18923 40477 18935 40480
rect 18877 40471 18935 40477
rect 14550 40372 14556 40384
rect 12728 40344 14556 40372
rect 14550 40332 14556 40344
rect 14608 40332 14614 40384
rect 15749 40375 15807 40381
rect 15749 40341 15761 40375
rect 15795 40372 15807 40375
rect 16022 40372 16028 40384
rect 15795 40344 16028 40372
rect 15795 40341 15807 40344
rect 15749 40335 15807 40341
rect 16022 40332 16028 40344
rect 16080 40372 16086 40384
rect 16206 40372 16212 40384
rect 16080 40344 16212 40372
rect 16080 40332 16086 40344
rect 16206 40332 16212 40344
rect 16264 40332 16270 40384
rect 17589 40375 17647 40381
rect 17589 40341 17601 40375
rect 17635 40372 17647 40375
rect 17954 40372 17960 40384
rect 17635 40344 17960 40372
rect 17635 40341 17647 40344
rect 17589 40335 17647 40341
rect 17954 40332 17960 40344
rect 18012 40332 18018 40384
rect 19352 40372 19380 40480
rect 22097 40477 22109 40511
rect 22143 40508 22155 40511
rect 23198 40508 23204 40520
rect 22143 40480 23204 40508
rect 22143 40477 22155 40480
rect 22097 40471 22155 40477
rect 23198 40468 23204 40480
rect 23256 40468 23262 40520
rect 24581 40511 24639 40517
rect 24581 40477 24593 40511
rect 24627 40508 24639 40511
rect 24854 40508 24860 40520
rect 24627 40480 24860 40508
rect 24627 40477 24639 40480
rect 24581 40471 24639 40477
rect 24854 40468 24860 40480
rect 24912 40468 24918 40520
rect 24946 40468 24952 40520
rect 25004 40508 25010 40520
rect 25148 40508 25176 40548
rect 25225 40545 25237 40548
rect 25271 40576 25283 40579
rect 25498 40576 25504 40588
rect 25271 40548 25504 40576
rect 25271 40545 25283 40548
rect 25225 40539 25283 40545
rect 25498 40536 25504 40548
rect 25556 40536 25562 40588
rect 26252 40585 26280 40616
rect 27172 40616 27344 40644
rect 27172 40585 27200 40616
rect 27338 40604 27344 40616
rect 27396 40604 27402 40656
rect 25593 40579 25651 40585
rect 25593 40545 25605 40579
rect 25639 40576 25651 40579
rect 26237 40579 26295 40585
rect 25639 40548 26188 40576
rect 25639 40545 25651 40548
rect 25593 40539 25651 40545
rect 25314 40508 25320 40520
rect 25004 40480 25176 40508
rect 25275 40480 25320 40508
rect 25004 40468 25010 40480
rect 25314 40468 25320 40480
rect 25372 40468 25378 40520
rect 25409 40511 25467 40517
rect 25409 40477 25421 40511
rect 25455 40508 25467 40511
rect 26050 40508 26056 40520
rect 25455 40480 26056 40508
rect 25455 40477 25467 40480
rect 25409 40471 25467 40477
rect 26050 40468 26056 40480
rect 26108 40468 26114 40520
rect 26160 40508 26188 40548
rect 26237 40545 26249 40579
rect 26283 40545 26295 40579
rect 26237 40539 26295 40545
rect 27157 40579 27215 40585
rect 27157 40545 27169 40579
rect 27203 40545 27215 40579
rect 27157 40539 27215 40545
rect 27246 40536 27252 40588
rect 27304 40576 27310 40588
rect 27304 40548 27349 40576
rect 27304 40536 27310 40548
rect 27430 40536 27436 40588
rect 27488 40576 27494 40588
rect 27525 40579 27583 40585
rect 27525 40576 27537 40579
rect 27488 40548 27537 40576
rect 27488 40536 27494 40548
rect 27525 40545 27537 40548
rect 27571 40545 27583 40579
rect 27525 40539 27583 40545
rect 28626 40536 28632 40588
rect 28684 40576 28690 40588
rect 29549 40579 29607 40585
rect 29549 40576 29561 40579
rect 28684 40548 29561 40576
rect 28684 40536 28690 40548
rect 29549 40545 29561 40548
rect 29595 40545 29607 40579
rect 29549 40539 29607 40545
rect 29816 40579 29874 40585
rect 29816 40545 29828 40579
rect 29862 40576 29874 40579
rect 30282 40576 30288 40588
rect 29862 40548 30288 40576
rect 29862 40545 29874 40548
rect 29816 40539 29874 40545
rect 30282 40536 30288 40548
rect 30340 40536 30346 40588
rect 26326 40508 26332 40520
rect 26160 40480 26332 40508
rect 26326 40468 26332 40480
rect 26384 40468 26390 40520
rect 28166 40508 28172 40520
rect 28127 40480 28172 40508
rect 28166 40468 28172 40480
rect 28224 40468 28230 40520
rect 28445 40511 28503 40517
rect 28445 40477 28457 40511
rect 28491 40508 28503 40511
rect 28534 40508 28540 40520
rect 28491 40480 28540 40508
rect 28491 40477 28503 40480
rect 28445 40471 28503 40477
rect 28534 40468 28540 40480
rect 28592 40508 28598 40520
rect 28902 40508 28908 40520
rect 28592 40480 28908 40508
rect 28592 40468 28598 40480
rect 28902 40468 28908 40480
rect 28960 40468 28966 40520
rect 26973 40443 27031 40449
rect 26973 40409 26985 40443
rect 27019 40440 27031 40443
rect 27614 40440 27620 40452
rect 27019 40412 27620 40440
rect 27019 40409 27031 40412
rect 26973 40403 27031 40409
rect 27614 40400 27620 40412
rect 27672 40400 27678 40452
rect 20070 40372 20076 40384
rect 19352 40344 20076 40372
rect 20070 40332 20076 40344
rect 20128 40332 20134 40384
rect 21174 40372 21180 40384
rect 21135 40344 21180 40372
rect 21174 40332 21180 40344
rect 21232 40332 21238 40384
rect 22002 40332 22008 40384
rect 22060 40372 22066 40384
rect 22278 40372 22284 40384
rect 22060 40344 22284 40372
rect 22060 40332 22066 40344
rect 22278 40332 22284 40344
rect 22336 40332 22342 40384
rect 23201 40375 23259 40381
rect 23201 40341 23213 40375
rect 23247 40372 23259 40375
rect 23290 40372 23296 40384
rect 23247 40344 23296 40372
rect 23247 40341 23259 40344
rect 23201 40335 23259 40341
rect 23290 40332 23296 40344
rect 23348 40332 23354 40384
rect 25774 40372 25780 40384
rect 25735 40344 25780 40372
rect 25774 40332 25780 40344
rect 25832 40332 25838 40384
rect 27338 40332 27344 40384
rect 27396 40372 27402 40384
rect 27433 40375 27491 40381
rect 27433 40372 27445 40375
rect 27396 40344 27445 40372
rect 27396 40332 27402 40344
rect 27433 40341 27445 40344
rect 27479 40341 27491 40375
rect 27433 40335 27491 40341
rect 30558 40332 30564 40384
rect 30616 40372 30622 40384
rect 30929 40375 30987 40381
rect 30929 40372 30941 40375
rect 30616 40344 30941 40372
rect 30616 40332 30622 40344
rect 30929 40341 30941 40344
rect 30975 40341 30987 40375
rect 30929 40335 30987 40341
rect 1104 40282 32016 40304
rect 1104 40230 6102 40282
rect 6154 40230 6166 40282
rect 6218 40230 6230 40282
rect 6282 40230 6294 40282
rect 6346 40230 6358 40282
rect 6410 40230 16405 40282
rect 16457 40230 16469 40282
rect 16521 40230 16533 40282
rect 16585 40230 16597 40282
rect 16649 40230 16661 40282
rect 16713 40230 26709 40282
rect 26761 40230 26773 40282
rect 26825 40230 26837 40282
rect 26889 40230 26901 40282
rect 26953 40230 26965 40282
rect 27017 40230 32016 40282
rect 1104 40208 32016 40230
rect 3145 40171 3203 40177
rect 3145 40137 3157 40171
rect 3191 40168 3203 40171
rect 4062 40168 4068 40180
rect 3191 40140 4068 40168
rect 3191 40137 3203 40140
rect 3145 40131 3203 40137
rect 4062 40128 4068 40140
rect 4120 40128 4126 40180
rect 9953 40171 10011 40177
rect 9232 40140 9674 40168
rect 4338 40060 4344 40112
rect 4396 40100 4402 40112
rect 4982 40100 4988 40112
rect 4396 40072 4988 40100
rect 4396 40060 4402 40072
rect 4982 40060 4988 40072
rect 5040 40060 5046 40112
rect 2133 40035 2191 40041
rect 2133 40001 2145 40035
rect 2179 40032 2191 40035
rect 2498 40032 2504 40044
rect 2179 40004 2504 40032
rect 2179 40001 2191 40004
rect 2133 39995 2191 40001
rect 2498 39992 2504 40004
rect 2556 39992 2562 40044
rect 4062 40032 4068 40044
rect 2746 40004 3832 40032
rect 4023 40004 4068 40032
rect 1857 39967 1915 39973
rect 1857 39933 1869 39967
rect 1903 39933 1915 39967
rect 1857 39927 1915 39933
rect 2041 39967 2099 39973
rect 2041 39933 2053 39967
rect 2087 39933 2099 39967
rect 2222 39964 2228 39976
rect 2183 39936 2228 39964
rect 2041 39927 2099 39933
rect 0 39828 800 39842
rect 1394 39828 1400 39840
rect 0 39800 1400 39828
rect 0 39786 800 39800
rect 1394 39788 1400 39800
rect 1452 39788 1458 39840
rect 1670 39828 1676 39840
rect 1631 39800 1676 39828
rect 1670 39788 1676 39800
rect 1728 39788 1734 39840
rect 1872 39828 1900 39927
rect 2056 39896 2084 39927
rect 2222 39924 2228 39936
rect 2280 39924 2286 39976
rect 2406 39964 2412 39976
rect 2367 39936 2412 39964
rect 2406 39924 2412 39936
rect 2464 39964 2470 39976
rect 2746 39964 2774 40004
rect 2464 39936 2774 39964
rect 3237 39967 3295 39973
rect 2464 39924 2470 39936
rect 3237 39933 3249 39967
rect 3283 39964 3295 39967
rect 3418 39964 3424 39976
rect 3283 39936 3424 39964
rect 3283 39933 3295 39936
rect 3237 39927 3295 39933
rect 3418 39924 3424 39936
rect 3476 39964 3482 39976
rect 3694 39964 3700 39976
rect 3476 39936 3700 39964
rect 3476 39924 3482 39936
rect 3694 39924 3700 39936
rect 3752 39924 3758 39976
rect 3804 39973 3832 40004
rect 4062 39992 4068 40004
rect 4120 39992 4126 40044
rect 4522 40032 4528 40044
rect 4483 40004 4528 40032
rect 4522 39992 4528 40004
rect 4580 39992 4586 40044
rect 5445 40035 5503 40041
rect 5445 40001 5457 40035
rect 5491 40032 5503 40035
rect 5626 40032 5632 40044
rect 5491 40004 5632 40032
rect 5491 40001 5503 40004
rect 5445 39995 5503 40001
rect 5626 39992 5632 40004
rect 5684 40032 5690 40044
rect 6638 40032 6644 40044
rect 5684 40004 6644 40032
rect 5684 39992 5690 40004
rect 6638 39992 6644 40004
rect 6696 39992 6702 40044
rect 3789 39967 3847 39973
rect 3789 39933 3801 39967
rect 3835 39964 3847 39967
rect 3878 39964 3884 39976
rect 3835 39936 3884 39964
rect 3835 39933 3847 39936
rect 3789 39927 3847 39933
rect 3878 39924 3884 39936
rect 3936 39924 3942 39976
rect 3970 39924 3976 39976
rect 4028 39964 4034 39976
rect 4157 39967 4215 39973
rect 4028 39936 4073 39964
rect 4028 39924 4034 39936
rect 4157 39933 4169 39967
rect 4203 39933 4215 39967
rect 4338 39964 4344 39976
rect 4299 39936 4344 39964
rect 4157 39927 4215 39933
rect 4172 39896 4200 39927
rect 4338 39924 4344 39936
rect 4396 39924 4402 39976
rect 4982 39924 4988 39976
rect 5040 39964 5046 39976
rect 5537 39967 5595 39973
rect 5537 39964 5549 39967
rect 5040 39936 5549 39964
rect 5040 39924 5046 39936
rect 5537 39933 5549 39936
rect 5583 39933 5595 39967
rect 7193 39967 7251 39973
rect 7193 39964 7205 39967
rect 5537 39927 5595 39933
rect 6012 39936 7205 39964
rect 2056 39868 2728 39896
rect 2700 39840 2728 39868
rect 3068 39868 4200 39896
rect 2590 39828 2596 39840
rect 1872 39800 2596 39828
rect 2590 39788 2596 39800
rect 2648 39788 2654 39840
rect 2682 39788 2688 39840
rect 2740 39828 2746 39840
rect 3068 39828 3096 39868
rect 2740 39800 3096 39828
rect 2740 39788 2746 39800
rect 5626 39788 5632 39840
rect 5684 39828 5690 39840
rect 6012 39837 6040 39936
rect 7193 39933 7205 39936
rect 7239 39933 7251 39967
rect 7193 39927 7251 39933
rect 7834 39924 7840 39976
rect 7892 39964 7898 39976
rect 9232 39973 9260 40140
rect 9398 40060 9404 40112
rect 9456 40060 9462 40112
rect 9416 39973 9444 40060
rect 9646 40044 9674 40140
rect 9953 40137 9965 40171
rect 9999 40168 10011 40171
rect 10318 40168 10324 40180
rect 9999 40140 10324 40168
rect 9999 40137 10011 40140
rect 9953 40131 10011 40137
rect 10318 40128 10324 40140
rect 10376 40128 10382 40180
rect 15749 40171 15807 40177
rect 15749 40137 15761 40171
rect 15795 40168 15807 40171
rect 16298 40168 16304 40180
rect 15795 40140 16304 40168
rect 15795 40137 15807 40140
rect 15749 40131 15807 40137
rect 16298 40128 16304 40140
rect 16356 40128 16362 40180
rect 16853 40171 16911 40177
rect 16853 40137 16865 40171
rect 16899 40168 16911 40171
rect 17310 40168 17316 40180
rect 16899 40140 17316 40168
rect 16899 40137 16911 40140
rect 16853 40131 16911 40137
rect 17310 40128 17316 40140
rect 17368 40128 17374 40180
rect 23106 40168 23112 40180
rect 23067 40140 23112 40168
rect 23106 40128 23112 40140
rect 23164 40128 23170 40180
rect 24762 40168 24768 40180
rect 23207 40140 24768 40168
rect 10134 40060 10140 40112
rect 10192 40100 10198 40112
rect 10413 40103 10471 40109
rect 10413 40100 10425 40103
rect 10192 40072 10425 40100
rect 10192 40060 10198 40072
rect 10413 40069 10425 40072
rect 10459 40069 10471 40103
rect 10413 40063 10471 40069
rect 14016 40072 14504 40100
rect 9646 40004 9680 40044
rect 9674 39992 9680 40004
rect 9732 39992 9738 40044
rect 12434 39992 12440 40044
rect 12492 40032 12498 40044
rect 12492 40004 12537 40032
rect 12492 39992 12498 40004
rect 12618 39992 12624 40044
rect 12676 40032 12682 40044
rect 14016 40032 14044 40072
rect 12676 40004 14044 40032
rect 14093 40035 14151 40041
rect 12676 39992 12682 40004
rect 14093 40001 14105 40035
rect 14139 40032 14151 40035
rect 14366 40032 14372 40044
rect 14139 40004 14372 40032
rect 14139 40001 14151 40004
rect 14093 39995 14151 40001
rect 14366 39992 14372 40004
rect 14424 39992 14430 40044
rect 8205 39967 8263 39973
rect 8205 39964 8217 39967
rect 7892 39936 8217 39964
rect 7892 39924 7898 39936
rect 8205 39933 8217 39936
rect 8251 39933 8263 39967
rect 8205 39927 8263 39933
rect 9217 39967 9275 39973
rect 9217 39933 9229 39967
rect 9263 39933 9275 39967
rect 9217 39927 9275 39933
rect 9401 39967 9459 39973
rect 9401 39933 9413 39967
rect 9447 39933 9459 39967
rect 9401 39927 9459 39933
rect 9487 39967 9545 39973
rect 9487 39954 9499 39967
rect 9533 39954 9545 39967
rect 9585 39967 9643 39973
rect 9585 39954 9597 39967
rect 9631 39954 9643 39967
rect 9769 39967 9827 39973
rect 9487 39927 9496 39954
rect 6638 39896 6644 39908
rect 6599 39868 6644 39896
rect 6638 39856 6644 39868
rect 6696 39856 6702 39908
rect 9490 39902 9496 39927
rect 9548 39902 9554 39954
rect 9582 39902 9588 39954
rect 9640 39902 9646 39954
rect 9769 39933 9781 39967
rect 9815 39933 9827 39967
rect 10778 39964 10784 39976
rect 10739 39936 10784 39964
rect 9769 39927 9827 39933
rect 9784 39896 9812 39927
rect 10778 39924 10784 39936
rect 10836 39964 10842 39976
rect 11333 39967 11391 39973
rect 11333 39964 11345 39967
rect 10836 39936 11345 39964
rect 10836 39924 10842 39936
rect 11333 39933 11345 39936
rect 11379 39933 11391 39967
rect 11333 39927 11391 39933
rect 11422 39924 11428 39976
rect 11480 39964 11486 39976
rect 11974 39964 11980 39976
rect 11480 39936 11980 39964
rect 11480 39924 11486 39936
rect 11974 39924 11980 39936
rect 12032 39924 12038 39976
rect 12713 39967 12771 39973
rect 12713 39933 12725 39967
rect 12759 39964 12771 39967
rect 12986 39964 12992 39976
rect 12759 39936 12992 39964
rect 12759 39933 12771 39936
rect 12713 39927 12771 39933
rect 12986 39924 12992 39936
rect 13044 39924 13050 39976
rect 13265 39967 13323 39973
rect 13265 39933 13277 39967
rect 13311 39964 13323 39967
rect 13998 39964 14004 39976
rect 13311 39936 14004 39964
rect 13311 39933 13323 39936
rect 13265 39927 13323 39933
rect 13998 39924 14004 39936
rect 14056 39924 14062 39976
rect 14274 39964 14280 39976
rect 14235 39936 14280 39964
rect 14274 39924 14280 39936
rect 14332 39924 14338 39976
rect 14476 39973 14504 40072
rect 14550 40060 14556 40112
rect 14608 40060 14614 40112
rect 21450 40060 21456 40112
rect 21508 40100 21514 40112
rect 23207 40100 23235 40140
rect 24762 40128 24768 40140
rect 24820 40128 24826 40180
rect 30282 40168 30288 40180
rect 30243 40140 30288 40168
rect 30282 40128 30288 40140
rect 30340 40128 30346 40180
rect 30374 40128 30380 40180
rect 30432 40168 30438 40180
rect 30650 40168 30656 40180
rect 30432 40140 30656 40168
rect 30432 40128 30438 40140
rect 30650 40128 30656 40140
rect 30708 40128 30714 40180
rect 21508 40072 23235 40100
rect 21508 40060 21514 40072
rect 23566 40060 23572 40112
rect 23624 40060 23630 40112
rect 14568 39973 14596 40060
rect 22097 40035 22155 40041
rect 22097 40001 22109 40035
rect 22143 40032 22155 40035
rect 22554 40032 22560 40044
rect 22143 40004 22560 40032
rect 22143 40001 22155 40004
rect 22097 39995 22155 40001
rect 14461 39967 14519 39973
rect 14461 39933 14473 39967
rect 14507 39933 14519 39967
rect 14461 39927 14519 39933
rect 14550 39967 14608 39973
rect 14550 39933 14562 39967
rect 14596 39933 14608 39967
rect 14550 39927 14608 39933
rect 14645 39967 14703 39973
rect 14645 39933 14657 39967
rect 14691 39964 14703 39967
rect 14734 39964 14740 39976
rect 14691 39936 14740 39964
rect 14691 39933 14703 39936
rect 14645 39927 14703 39933
rect 14734 39924 14740 39936
rect 14792 39924 14798 39976
rect 14829 39967 14887 39973
rect 14829 39933 14841 39967
rect 14875 39933 14887 39967
rect 14829 39927 14887 39933
rect 15933 39967 15991 39973
rect 15933 39933 15945 39967
rect 15979 39964 15991 39967
rect 16942 39964 16948 39976
rect 15979 39936 16948 39964
rect 15979 39933 15991 39936
rect 15933 39927 15991 39933
rect 9692 39868 9812 39896
rect 10597 39899 10655 39905
rect 5997 39831 6055 39837
rect 5684 39800 5729 39828
rect 5684 39788 5690 39800
rect 5997 39797 6009 39831
rect 6043 39797 6055 39831
rect 5997 39791 6055 39797
rect 6362 39788 6368 39840
rect 6420 39828 6426 39840
rect 6549 39831 6607 39837
rect 6549 39828 6561 39831
rect 6420 39800 6561 39828
rect 6420 39788 6426 39800
rect 6549 39797 6561 39800
rect 6595 39797 6607 39831
rect 6549 39791 6607 39797
rect 7006 39788 7012 39840
rect 7064 39828 7070 39840
rect 7285 39831 7343 39837
rect 7285 39828 7297 39831
rect 7064 39800 7297 39828
rect 7064 39788 7070 39800
rect 7285 39797 7297 39800
rect 7331 39797 7343 39831
rect 7285 39791 7343 39797
rect 8297 39831 8355 39837
rect 8297 39797 8309 39831
rect 8343 39828 8355 39831
rect 9692 39828 9720 39868
rect 10597 39865 10609 39899
rect 10643 39896 10655 39899
rect 10686 39896 10692 39908
rect 10643 39868 10692 39896
rect 10643 39865 10655 39868
rect 10597 39859 10655 39865
rect 10686 39856 10692 39868
rect 10744 39856 10750 39908
rect 13538 39856 13544 39908
rect 13596 39896 13602 39908
rect 14844 39896 14872 39927
rect 16942 39924 16948 39936
rect 17000 39964 17006 39976
rect 17586 39964 17592 39976
rect 17000 39936 17592 39964
rect 17000 39924 17006 39936
rect 17586 39924 17592 39936
rect 17644 39924 17650 39976
rect 17954 39924 17960 39976
rect 18012 39973 18018 39976
rect 18012 39964 18024 39973
rect 18233 39967 18291 39973
rect 18012 39936 18057 39964
rect 18012 39927 18024 39936
rect 18233 39933 18245 39967
rect 18279 39964 18291 39967
rect 19518 39964 19524 39976
rect 18279 39936 19524 39964
rect 18279 39933 18291 39936
rect 18233 39927 18291 39933
rect 18012 39924 18018 39927
rect 19518 39924 19524 39936
rect 19576 39924 19582 39976
rect 21174 39964 21180 39976
rect 20548 39936 21180 39964
rect 13596 39868 14872 39896
rect 16117 39899 16175 39905
rect 13596 39856 13602 39868
rect 16117 39865 16129 39899
rect 16163 39896 16175 39899
rect 17678 39896 17684 39908
rect 16163 39868 17684 39896
rect 16163 39865 16175 39868
rect 16117 39859 16175 39865
rect 17678 39856 17684 39868
rect 17736 39856 17742 39908
rect 19334 39856 19340 39908
rect 19392 39896 19398 39908
rect 19610 39896 19616 39908
rect 19392 39868 19616 39896
rect 19392 39856 19398 39868
rect 19610 39856 19616 39868
rect 19668 39856 19674 39908
rect 8343 39800 9720 39828
rect 13357 39831 13415 39837
rect 8343 39797 8355 39800
rect 8297 39791 8355 39797
rect 13357 39797 13369 39831
rect 13403 39828 13415 39831
rect 13446 39828 13452 39840
rect 13403 39800 13452 39828
rect 13403 39797 13415 39800
rect 13357 39791 13415 39797
rect 13446 39788 13452 39800
rect 13504 39828 13510 39840
rect 13722 39828 13728 39840
rect 13504 39800 13728 39828
rect 13504 39788 13510 39800
rect 13722 39788 13728 39800
rect 13780 39788 13786 39840
rect 13998 39788 14004 39840
rect 14056 39828 14062 39840
rect 20548 39828 20576 39936
rect 21174 39924 21180 39936
rect 21232 39924 21238 39976
rect 21821 39967 21879 39973
rect 21821 39933 21833 39967
rect 21867 39964 21879 39967
rect 21910 39964 21916 39976
rect 21867 39936 21916 39964
rect 21867 39933 21879 39936
rect 21821 39927 21879 39933
rect 21910 39924 21916 39936
rect 21968 39924 21974 39976
rect 22005 39967 22063 39973
rect 22005 39933 22017 39967
rect 22051 39933 22063 39967
rect 22005 39927 22063 39933
rect 20714 39856 20720 39908
rect 20772 39896 20778 39908
rect 22020 39896 22048 39927
rect 20772 39868 22048 39896
rect 20772 39856 20778 39868
rect 14056 39800 20576 39828
rect 14056 39788 14062 39800
rect 20622 39788 20628 39840
rect 20680 39828 20686 39840
rect 20901 39831 20959 39837
rect 20901 39828 20913 39831
rect 20680 39800 20913 39828
rect 20680 39788 20686 39800
rect 20901 39797 20913 39800
rect 20947 39797 20959 39831
rect 20901 39791 20959 39797
rect 22002 39788 22008 39840
rect 22060 39828 22066 39840
rect 22112 39828 22140 39995
rect 22554 39992 22560 40004
rect 22612 39992 22618 40044
rect 23477 40035 23535 40041
rect 23477 40001 23489 40035
rect 23523 40032 23535 40035
rect 23584 40032 23612 40060
rect 23523 40004 23612 40032
rect 23523 40001 23535 40004
rect 23477 39995 23535 40001
rect 23934 39992 23940 40044
rect 23992 40032 23998 40044
rect 23992 40004 24440 40032
rect 23992 39992 23998 40004
rect 22186 39924 22192 39976
rect 22244 39964 22250 39976
rect 22373 39967 22431 39973
rect 22244 39936 22289 39964
rect 22244 39924 22250 39936
rect 22373 39933 22385 39967
rect 22419 39964 22431 39967
rect 23106 39964 23112 39976
rect 22419 39936 23112 39964
rect 22419 39933 22431 39936
rect 22373 39927 22431 39933
rect 23106 39924 23112 39936
rect 23164 39924 23170 39976
rect 23290 39964 23296 39976
rect 23251 39936 23296 39964
rect 23290 39924 23296 39936
rect 23348 39924 23354 39976
rect 23569 39967 23627 39973
rect 23569 39933 23581 39967
rect 23615 39933 23627 39967
rect 23569 39927 23627 39933
rect 22204 39896 22232 39924
rect 22922 39896 22928 39908
rect 22204 39868 22928 39896
rect 22922 39856 22928 39868
rect 22980 39856 22986 39908
rect 23584 39896 23612 39927
rect 23658 39924 23664 39976
rect 23716 39964 23722 39976
rect 23845 39967 23903 39973
rect 23716 39936 23761 39964
rect 23716 39924 23722 39936
rect 23845 39933 23857 39967
rect 23891 39964 23903 39967
rect 24210 39964 24216 39976
rect 23891 39936 24216 39964
rect 23891 39933 23903 39936
rect 23845 39927 23903 39933
rect 24210 39924 24216 39936
rect 24268 39924 24274 39976
rect 24412 39973 24440 40004
rect 26234 39992 26240 40044
rect 26292 40032 26298 40044
rect 27617 40035 27675 40041
rect 27617 40032 27629 40035
rect 26292 40004 27629 40032
rect 26292 39992 26298 40004
rect 27617 40001 27629 40004
rect 27663 40001 27675 40035
rect 27617 39995 27675 40001
rect 27893 40035 27951 40041
rect 27893 40001 27905 40035
rect 27939 40032 27951 40035
rect 28166 40032 28172 40044
rect 27939 40004 28172 40032
rect 27939 40001 27951 40004
rect 27893 39995 27951 40001
rect 28166 39992 28172 40004
rect 28224 39992 28230 40044
rect 29454 40032 29460 40044
rect 28368 40004 29460 40032
rect 24397 39967 24455 39973
rect 24397 39933 24409 39967
rect 24443 39933 24455 39967
rect 24578 39964 24584 39976
rect 24539 39936 24584 39964
rect 24397 39927 24455 39933
rect 24578 39924 24584 39936
rect 24636 39924 24642 39976
rect 24854 39924 24860 39976
rect 24912 39964 24918 39976
rect 25041 39967 25099 39973
rect 25041 39964 25053 39967
rect 24912 39936 25053 39964
rect 24912 39924 24918 39936
rect 25041 39933 25053 39936
rect 25087 39933 25099 39967
rect 25041 39927 25099 39933
rect 25308 39967 25366 39973
rect 25308 39933 25320 39967
rect 25354 39964 25366 39967
rect 25774 39964 25780 39976
rect 25354 39936 25780 39964
rect 25354 39933 25366 39936
rect 25308 39927 25366 39933
rect 25774 39924 25780 39936
rect 25832 39924 25838 39976
rect 26510 39924 26516 39976
rect 26568 39964 26574 39976
rect 28368 39964 28396 40004
rect 29454 39992 29460 40004
rect 29512 39992 29518 40044
rect 31018 40032 31024 40044
rect 29748 40004 31024 40032
rect 26568 39936 28396 39964
rect 26568 39924 26574 39936
rect 28442 39924 28448 39976
rect 28500 39964 28506 39976
rect 28537 39967 28595 39973
rect 28537 39964 28549 39967
rect 28500 39936 28549 39964
rect 28500 39924 28506 39936
rect 28537 39933 28549 39936
rect 28583 39933 28595 39967
rect 28537 39927 28595 39933
rect 29270 39924 29276 39976
rect 29328 39964 29334 39976
rect 29748 39973 29776 40004
rect 31018 39992 31024 40004
rect 31076 39992 31082 40044
rect 29549 39967 29607 39973
rect 29549 39964 29561 39967
rect 29328 39936 29561 39964
rect 29328 39924 29334 39936
rect 29549 39933 29561 39936
rect 29595 39933 29607 39967
rect 29549 39927 29607 39933
rect 29733 39967 29791 39973
rect 29733 39933 29745 39967
rect 29779 39933 29791 39967
rect 29733 39927 29791 39933
rect 29825 39967 29883 39973
rect 29825 39933 29837 39967
rect 29871 39933 29883 39967
rect 29825 39927 29883 39933
rect 23584 39868 25360 39896
rect 25332 39840 25360 39868
rect 28626 39856 28632 39908
rect 28684 39896 28690 39908
rect 29840 39896 29868 39927
rect 29914 39924 29920 39976
rect 29972 39964 29978 39976
rect 30101 39967 30159 39973
rect 29972 39936 30017 39964
rect 29972 39924 29978 39936
rect 30101 39933 30113 39967
rect 30147 39964 30159 39967
rect 30466 39964 30472 39976
rect 30147 39936 30472 39964
rect 30147 39933 30159 39936
rect 30101 39927 30159 39933
rect 30466 39924 30472 39936
rect 30524 39924 30530 39976
rect 31113 39967 31171 39973
rect 31113 39933 31125 39967
rect 31159 39964 31171 39967
rect 31294 39964 31300 39976
rect 31159 39936 31300 39964
rect 31159 39933 31171 39936
rect 31113 39927 31171 39933
rect 31294 39924 31300 39936
rect 31352 39924 31358 39976
rect 28684 39868 29868 39896
rect 28684 39856 28690 39868
rect 22554 39828 22560 39840
rect 22060 39800 22140 39828
rect 22515 39800 22560 39828
rect 22060 39788 22066 39800
rect 22554 39788 22560 39800
rect 22612 39788 22618 39840
rect 22830 39788 22836 39840
rect 22888 39828 22894 39840
rect 24397 39831 24455 39837
rect 24397 39828 24409 39831
rect 22888 39800 24409 39828
rect 22888 39788 22894 39800
rect 24397 39797 24409 39800
rect 24443 39797 24455 39831
rect 24397 39791 24455 39797
rect 25314 39788 25320 39840
rect 25372 39788 25378 39840
rect 26326 39788 26332 39840
rect 26384 39828 26390 39840
rect 26421 39831 26479 39837
rect 26421 39828 26433 39831
rect 26384 39800 26433 39828
rect 26384 39788 26390 39800
rect 26421 39797 26433 39800
rect 26467 39797 26479 39831
rect 26421 39791 26479 39797
rect 27430 39788 27436 39840
rect 27488 39828 27494 39840
rect 28445 39831 28503 39837
rect 28445 39828 28457 39831
rect 27488 39800 28457 39828
rect 27488 39788 27494 39800
rect 28445 39797 28457 39800
rect 28491 39828 28503 39831
rect 29638 39828 29644 39840
rect 28491 39800 29644 39828
rect 28491 39797 28503 39800
rect 28445 39791 28503 39797
rect 29638 39788 29644 39800
rect 29696 39788 29702 39840
rect 31297 39831 31355 39837
rect 31297 39797 31309 39831
rect 31343 39828 31355 39831
rect 32320 39828 33120 39842
rect 31343 39800 33120 39828
rect 31343 39797 31355 39800
rect 31297 39791 31355 39797
rect 32320 39786 33120 39800
rect 1104 39738 32016 39760
rect 1104 39686 11253 39738
rect 11305 39686 11317 39738
rect 11369 39686 11381 39738
rect 11433 39686 11445 39738
rect 11497 39686 11509 39738
rect 11561 39686 21557 39738
rect 21609 39686 21621 39738
rect 21673 39686 21685 39738
rect 21737 39686 21749 39738
rect 21801 39686 21813 39738
rect 21865 39686 32016 39738
rect 1104 39664 32016 39686
rect 3234 39624 3240 39636
rect 3195 39596 3240 39624
rect 3234 39584 3240 39596
rect 3292 39584 3298 39636
rect 4246 39584 4252 39636
rect 4304 39624 4310 39636
rect 4522 39624 4528 39636
rect 4304 39596 4528 39624
rect 4304 39584 4310 39596
rect 4522 39584 4528 39596
rect 4580 39584 4586 39636
rect 9582 39584 9588 39636
rect 9640 39624 9646 39636
rect 10137 39627 10195 39633
rect 10137 39624 10149 39627
rect 9640 39596 10149 39624
rect 9640 39584 9646 39596
rect 10137 39593 10149 39596
rect 10183 39593 10195 39627
rect 10137 39587 10195 39593
rect 14461 39627 14519 39633
rect 14461 39593 14473 39627
rect 14507 39624 14519 39627
rect 15194 39624 15200 39636
rect 14507 39596 15200 39624
rect 14507 39593 14519 39596
rect 14461 39587 14519 39593
rect 15194 39584 15200 39596
rect 15252 39584 15258 39636
rect 22097 39627 22155 39633
rect 22097 39593 22109 39627
rect 22143 39624 22155 39627
rect 22462 39624 22468 39636
rect 22143 39596 22468 39624
rect 22143 39593 22155 39596
rect 22097 39587 22155 39593
rect 22462 39584 22468 39596
rect 22520 39584 22526 39636
rect 22646 39584 22652 39636
rect 22704 39624 22710 39636
rect 23934 39624 23940 39636
rect 22704 39596 23940 39624
rect 22704 39584 22710 39596
rect 23934 39584 23940 39596
rect 23992 39584 23998 39636
rect 24302 39624 24308 39636
rect 24263 39596 24308 39624
rect 24302 39584 24308 39596
rect 24360 39584 24366 39636
rect 28166 39624 28172 39636
rect 26252 39596 28172 39624
rect 2774 39556 2780 39568
rect 1412 39528 2780 39556
rect 1412 39500 1440 39528
rect 2774 39516 2780 39528
rect 2832 39516 2838 39568
rect 3142 39516 3148 39568
rect 3200 39556 3206 39568
rect 3326 39556 3332 39568
rect 3200 39528 3332 39556
rect 3200 39516 3206 39528
rect 3326 39516 3332 39528
rect 3384 39556 3390 39568
rect 3384 39528 3832 39556
rect 3384 39516 3390 39528
rect 1394 39488 1400 39500
rect 1307 39460 1400 39488
rect 1394 39448 1400 39460
rect 1452 39448 1458 39500
rect 1670 39497 1676 39500
rect 1664 39488 1676 39497
rect 1631 39460 1676 39488
rect 1664 39451 1676 39460
rect 1670 39448 1676 39451
rect 1728 39448 1734 39500
rect 2130 39448 2136 39500
rect 2188 39488 2194 39500
rect 2682 39488 2688 39500
rect 2188 39460 2688 39488
rect 2188 39448 2194 39460
rect 2682 39448 2688 39460
rect 2740 39488 2746 39500
rect 3418 39488 3424 39500
rect 2740 39448 2774 39488
rect 3379 39460 3424 39488
rect 3418 39448 3424 39460
rect 3476 39448 3482 39500
rect 3804 39497 3832 39528
rect 4338 39516 4344 39568
rect 4396 39556 4402 39568
rect 5074 39556 5080 39568
rect 4396 39528 5080 39556
rect 4396 39516 4402 39528
rect 5074 39516 5080 39528
rect 5132 39556 5138 39568
rect 6362 39556 6368 39568
rect 5132 39528 6368 39556
rect 5132 39516 5138 39528
rect 3789 39491 3847 39497
rect 3789 39457 3801 39491
rect 3835 39457 3847 39491
rect 3789 39451 3847 39457
rect 3878 39448 3884 39500
rect 3936 39488 3942 39500
rect 3973 39491 4031 39497
rect 3973 39488 3985 39491
rect 3936 39460 3985 39488
rect 3936 39448 3942 39460
rect 3973 39457 3985 39460
rect 4019 39457 4031 39491
rect 4982 39488 4988 39500
rect 4943 39460 4988 39488
rect 3973 39451 4031 39457
rect 4982 39448 4988 39460
rect 5040 39448 5046 39500
rect 5368 39497 5396 39528
rect 6362 39516 6368 39528
rect 6420 39516 6426 39568
rect 12434 39556 12440 39568
rect 12406 39516 12440 39556
rect 12492 39516 12498 39568
rect 17126 39516 17132 39568
rect 17184 39556 17190 39568
rect 18322 39556 18328 39568
rect 17184 39528 18328 39556
rect 17184 39516 17190 39528
rect 18322 39516 18328 39528
rect 18380 39516 18386 39568
rect 19702 39516 19708 39568
rect 19760 39556 19766 39568
rect 23382 39556 23388 39568
rect 19760 39528 23244 39556
rect 23343 39528 23388 39556
rect 19760 39516 19766 39528
rect 5353 39491 5411 39497
rect 5353 39457 5365 39491
rect 5399 39457 5411 39491
rect 5353 39451 5411 39457
rect 5629 39491 5687 39497
rect 5629 39457 5641 39491
rect 5675 39488 5687 39491
rect 6733 39491 6791 39497
rect 6733 39488 6745 39491
rect 5675 39460 6745 39488
rect 5675 39457 5687 39460
rect 5629 39451 5687 39457
rect 6733 39457 6745 39460
rect 6779 39457 6791 39491
rect 7006 39488 7012 39500
rect 6967 39460 7012 39488
rect 6733 39451 6791 39457
rect 7006 39448 7012 39460
rect 7064 39448 7070 39500
rect 7466 39488 7472 39500
rect 7427 39460 7472 39488
rect 7466 39448 7472 39460
rect 7524 39448 7530 39500
rect 8294 39488 8300 39500
rect 8255 39460 8300 39488
rect 8294 39448 8300 39460
rect 8352 39448 8358 39500
rect 8386 39448 8392 39500
rect 8444 39488 8450 39500
rect 8553 39491 8611 39497
rect 8553 39488 8565 39491
rect 8444 39460 8565 39488
rect 8444 39448 8450 39460
rect 8553 39457 8565 39460
rect 8599 39457 8611 39491
rect 8553 39451 8611 39457
rect 10321 39491 10379 39497
rect 10321 39457 10333 39491
rect 10367 39488 10379 39491
rect 10410 39488 10416 39500
rect 10367 39460 10416 39488
rect 10367 39457 10379 39460
rect 10321 39451 10379 39457
rect 10410 39448 10416 39460
rect 10468 39448 10474 39500
rect 10505 39491 10563 39497
rect 10505 39457 10517 39491
rect 10551 39488 10563 39491
rect 11146 39488 11152 39500
rect 10551 39460 11152 39488
rect 10551 39457 10563 39460
rect 10505 39451 10563 39457
rect 11146 39448 11152 39460
rect 11204 39448 11210 39500
rect 11793 39491 11851 39497
rect 11793 39457 11805 39491
rect 11839 39488 11851 39491
rect 12406 39488 12434 39516
rect 11839 39460 12434 39488
rect 11839 39457 11851 39460
rect 11793 39451 11851 39457
rect 13814 39448 13820 39500
rect 13872 39488 13878 39500
rect 14369 39491 14427 39497
rect 14369 39488 14381 39491
rect 13872 39460 14381 39488
rect 13872 39448 13878 39460
rect 14369 39457 14381 39460
rect 14415 39457 14427 39491
rect 14369 39451 14427 39457
rect 15102 39448 15108 39500
rect 15160 39488 15166 39500
rect 15657 39491 15715 39497
rect 15657 39488 15669 39491
rect 15160 39460 15669 39488
rect 15160 39448 15166 39460
rect 15657 39457 15669 39460
rect 15703 39457 15715 39491
rect 15657 39451 15715 39457
rect 15841 39491 15899 39497
rect 15841 39457 15853 39491
rect 15887 39488 15899 39491
rect 15930 39488 15936 39500
rect 15887 39460 15936 39488
rect 15887 39457 15899 39460
rect 15841 39451 15899 39457
rect 15930 39448 15936 39460
rect 15988 39448 15994 39500
rect 18230 39488 18236 39500
rect 18288 39497 18294 39500
rect 18200 39460 18236 39488
rect 18230 39448 18236 39460
rect 18288 39451 18300 39497
rect 20530 39488 20536 39500
rect 20588 39497 20594 39500
rect 20500 39460 20536 39488
rect 18288 39448 18294 39451
rect 20530 39448 20536 39460
rect 20588 39451 20600 39497
rect 22281 39491 22339 39497
rect 22281 39457 22293 39491
rect 22327 39457 22339 39491
rect 22281 39451 22339 39457
rect 20588 39448 20594 39451
rect 2746 39420 2774 39448
rect 3605 39423 3663 39429
rect 3605 39420 3617 39423
rect 2746 39392 3617 39420
rect 3605 39389 3617 39392
rect 3651 39389 3663 39423
rect 3605 39383 3663 39389
rect 3697 39423 3755 39429
rect 3697 39389 3709 39423
rect 3743 39420 3755 39423
rect 4246 39420 4252 39432
rect 3743 39392 4252 39420
rect 3743 39389 3755 39392
rect 3697 39383 3755 39389
rect 4246 39380 4252 39392
rect 4304 39380 4310 39432
rect 5169 39423 5227 39429
rect 5169 39389 5181 39423
rect 5215 39389 5227 39423
rect 5169 39383 5227 39389
rect 5813 39423 5871 39429
rect 5813 39389 5825 39423
rect 5859 39420 5871 39423
rect 6454 39420 6460 39432
rect 5859 39392 6460 39420
rect 5859 39389 5871 39392
rect 5813 39383 5871 39389
rect 4982 39312 4988 39364
rect 5040 39352 5046 39364
rect 5184 39352 5212 39383
rect 6454 39380 6460 39392
rect 6512 39380 6518 39432
rect 7190 39420 7196 39432
rect 7151 39392 7196 39420
rect 7190 39380 7196 39392
rect 7248 39380 7254 39432
rect 12069 39423 12127 39429
rect 12069 39389 12081 39423
rect 12115 39420 12127 39423
rect 12434 39420 12440 39432
rect 12115 39392 12440 39420
rect 12115 39389 12127 39392
rect 12069 39383 12127 39389
rect 12434 39380 12440 39392
rect 12492 39380 12498 39432
rect 13446 39380 13452 39432
rect 13504 39420 13510 39432
rect 13633 39423 13691 39429
rect 13633 39420 13645 39423
rect 13504 39392 13645 39420
rect 13504 39380 13510 39392
rect 13633 39389 13645 39392
rect 13679 39389 13691 39423
rect 13633 39383 13691 39389
rect 13722 39380 13728 39432
rect 13780 39420 13786 39432
rect 13909 39423 13967 39429
rect 13909 39420 13921 39423
rect 13780 39392 13921 39420
rect 13780 39380 13786 39392
rect 13909 39389 13921 39392
rect 13955 39420 13967 39423
rect 15562 39420 15568 39432
rect 13955 39392 15568 39420
rect 13955 39389 13967 39392
rect 13909 39383 13967 39389
rect 15562 39380 15568 39392
rect 15620 39380 15626 39432
rect 18509 39423 18567 39429
rect 18509 39389 18521 39423
rect 18555 39420 18567 39423
rect 19610 39420 19616 39432
rect 18555 39392 19616 39420
rect 18555 39389 18567 39392
rect 18509 39383 18567 39389
rect 19610 39380 19616 39392
rect 19668 39380 19674 39432
rect 20809 39423 20867 39429
rect 20809 39389 20821 39423
rect 20855 39389 20867 39423
rect 20809 39383 20867 39389
rect 5040 39324 5212 39352
rect 7837 39355 7895 39361
rect 5040 39312 5046 39324
rect 7837 39321 7849 39355
rect 7883 39352 7895 39355
rect 8202 39352 8208 39364
rect 7883 39324 8208 39352
rect 7883 39321 7895 39324
rect 7837 39315 7895 39321
rect 8202 39312 8208 39324
rect 8260 39312 8266 39364
rect 14826 39312 14832 39364
rect 14884 39352 14890 39364
rect 15378 39352 15384 39364
rect 14884 39324 15384 39352
rect 14884 39312 14890 39324
rect 15378 39312 15384 39324
rect 15436 39312 15442 39364
rect 2682 39244 2688 39296
rect 2740 39284 2746 39296
rect 2777 39287 2835 39293
rect 2777 39284 2789 39287
rect 2740 39256 2789 39284
rect 2740 39244 2746 39256
rect 2777 39253 2789 39256
rect 2823 39253 2835 39287
rect 2777 39247 2835 39253
rect 3786 39244 3792 39296
rect 3844 39284 3850 39296
rect 4062 39284 4068 39296
rect 3844 39256 4068 39284
rect 3844 39244 3850 39256
rect 4062 39244 4068 39256
rect 4120 39284 4126 39296
rect 4433 39287 4491 39293
rect 4433 39284 4445 39287
rect 4120 39256 4445 39284
rect 4120 39244 4126 39256
rect 4433 39253 4445 39256
rect 4479 39253 4491 39287
rect 4433 39247 4491 39253
rect 8938 39244 8944 39296
rect 8996 39284 9002 39296
rect 9677 39287 9735 39293
rect 9677 39284 9689 39287
rect 8996 39256 9689 39284
rect 8996 39244 9002 39256
rect 9677 39253 9689 39256
rect 9723 39253 9735 39287
rect 9677 39247 9735 39253
rect 15194 39244 15200 39296
rect 15252 39284 15258 39296
rect 15473 39287 15531 39293
rect 15473 39284 15485 39287
rect 15252 39256 15485 39284
rect 15252 39244 15258 39256
rect 15473 39253 15485 39256
rect 15519 39253 15531 39287
rect 15654 39284 15660 39296
rect 15615 39256 15660 39284
rect 15473 39247 15531 39253
rect 15654 39244 15660 39256
rect 15712 39244 15718 39296
rect 17129 39287 17187 39293
rect 17129 39253 17141 39287
rect 17175 39284 17187 39287
rect 18138 39284 18144 39296
rect 17175 39256 18144 39284
rect 17175 39253 17187 39256
rect 17129 39247 17187 39253
rect 18138 39244 18144 39256
rect 18196 39244 18202 39296
rect 18506 39244 18512 39296
rect 18564 39284 18570 39296
rect 19429 39287 19487 39293
rect 19429 39284 19441 39287
rect 18564 39256 19441 39284
rect 18564 39244 18570 39256
rect 19429 39253 19441 39256
rect 19475 39253 19487 39287
rect 19429 39247 19487 39253
rect 19610 39244 19616 39296
rect 19668 39284 19674 39296
rect 20622 39284 20628 39296
rect 19668 39256 20628 39284
rect 19668 39244 19674 39256
rect 20622 39244 20628 39256
rect 20680 39284 20686 39296
rect 20824 39284 20852 39383
rect 20680 39256 20852 39284
rect 22296 39284 22324 39451
rect 22370 39448 22376 39500
rect 22428 39448 22434 39500
rect 22554 39488 22560 39500
rect 22515 39460 22560 39488
rect 22554 39448 22560 39460
rect 22612 39448 22618 39500
rect 22738 39488 22744 39500
rect 22699 39460 22744 39488
rect 22738 39448 22744 39460
rect 22796 39448 22802 39500
rect 23216 39488 23244 39528
rect 23382 39516 23388 39528
rect 23440 39516 23446 39568
rect 23474 39516 23480 39568
rect 23532 39556 23538 39568
rect 23569 39559 23627 39565
rect 23569 39556 23581 39559
rect 23532 39528 23581 39556
rect 23532 39516 23538 39528
rect 23569 39525 23581 39528
rect 23615 39556 23627 39559
rect 24946 39556 24952 39568
rect 23615 39528 24952 39556
rect 23615 39525 23627 39528
rect 23569 39519 23627 39525
rect 24946 39516 24952 39528
rect 25004 39516 25010 39568
rect 26142 39556 26148 39568
rect 26103 39528 26148 39556
rect 26142 39516 26148 39528
rect 26200 39516 26206 39568
rect 23658 39488 23664 39500
rect 23216 39460 23664 39488
rect 23658 39448 23664 39460
rect 23716 39448 23722 39500
rect 24213 39491 24271 39497
rect 24213 39457 24225 39491
rect 24259 39457 24271 39491
rect 24213 39451 24271 39457
rect 22388 39420 22416 39448
rect 22465 39423 22523 39429
rect 22465 39420 22477 39423
rect 22388 39392 22477 39420
rect 22465 39389 22477 39392
rect 22511 39389 22523 39423
rect 23198 39420 23204 39432
rect 22465 39383 22523 39389
rect 22572 39392 23204 39420
rect 22572 39364 22600 39392
rect 23198 39380 23204 39392
rect 23256 39420 23262 39432
rect 24228 39420 24256 39451
rect 25314 39448 25320 39500
rect 25372 39488 25378 39500
rect 25409 39491 25467 39497
rect 25409 39488 25421 39491
rect 25372 39460 25421 39488
rect 25372 39448 25378 39460
rect 25409 39457 25421 39460
rect 25455 39457 25467 39491
rect 25409 39451 25467 39457
rect 25685 39491 25743 39497
rect 25685 39457 25697 39491
rect 25731 39488 25743 39491
rect 26252 39488 26280 39596
rect 28166 39584 28172 39596
rect 28224 39624 28230 39636
rect 28350 39624 28356 39636
rect 28224 39596 28356 39624
rect 28224 39584 28230 39596
rect 28350 39584 28356 39596
rect 28408 39584 28414 39636
rect 28994 39624 29000 39636
rect 28955 39596 29000 39624
rect 28994 39584 29000 39596
rect 29052 39584 29058 39636
rect 29454 39584 29460 39636
rect 29512 39624 29518 39636
rect 29512 39596 29868 39624
rect 29512 39584 29518 39596
rect 27246 39516 27252 39568
rect 27304 39556 27310 39568
rect 29178 39556 29184 39568
rect 27304 39528 28120 39556
rect 27304 39516 27310 39528
rect 25731 39460 26280 39488
rect 26329 39491 26387 39497
rect 25731 39457 25743 39460
rect 25685 39451 25743 39457
rect 26329 39457 26341 39491
rect 26375 39488 26387 39491
rect 26418 39488 26424 39500
rect 26375 39460 26424 39488
rect 26375 39457 26387 39460
rect 26329 39451 26387 39457
rect 26418 39448 26424 39460
rect 26476 39448 26482 39500
rect 27154 39488 27160 39500
rect 27115 39460 27160 39488
rect 27154 39448 27160 39460
rect 27212 39448 27218 39500
rect 27522 39488 27528 39500
rect 27483 39460 27528 39488
rect 27522 39448 27528 39460
rect 27580 39448 27586 39500
rect 27706 39488 27712 39500
rect 27667 39460 27712 39488
rect 27706 39448 27712 39460
rect 27764 39448 27770 39500
rect 23256 39392 24256 39420
rect 27341 39423 27399 39429
rect 23256 39380 23262 39392
rect 27341 39389 27353 39423
rect 27387 39389 27399 39423
rect 27341 39383 27399 39389
rect 27433 39423 27491 39429
rect 27433 39389 27445 39423
rect 27479 39420 27491 39423
rect 27982 39420 27988 39432
rect 27479 39392 27988 39420
rect 27479 39389 27491 39392
rect 27433 39383 27491 39389
rect 22373 39355 22431 39361
rect 22373 39321 22385 39355
rect 22419 39352 22431 39355
rect 22554 39352 22560 39364
rect 22419 39324 22560 39352
rect 22419 39321 22431 39324
rect 22373 39315 22431 39321
rect 22554 39312 22560 39324
rect 22612 39312 22618 39364
rect 23106 39312 23112 39364
rect 23164 39352 23170 39364
rect 24394 39352 24400 39364
rect 23164 39324 24400 39352
rect 23164 39312 23170 39324
rect 24394 39312 24400 39324
rect 24452 39312 24458 39364
rect 27356 39352 27384 39383
rect 27982 39380 27988 39392
rect 28040 39380 28046 39432
rect 27798 39352 27804 39364
rect 27356 39324 27804 39352
rect 27798 39312 27804 39324
rect 27856 39312 27862 39364
rect 22462 39284 22468 39296
rect 22296 39256 22468 39284
rect 20680 39244 20686 39256
rect 22462 39244 22468 39256
rect 22520 39284 22526 39296
rect 23014 39284 23020 39296
rect 22520 39256 23020 39284
rect 22520 39244 22526 39256
rect 23014 39244 23020 39256
rect 23072 39244 23078 39296
rect 26973 39287 27031 39293
rect 26973 39253 26985 39287
rect 27019 39284 27031 39287
rect 27430 39284 27436 39296
rect 27019 39256 27436 39284
rect 27019 39253 27031 39256
rect 26973 39247 27031 39253
rect 27430 39244 27436 39256
rect 27488 39244 27494 39296
rect 28092 39284 28120 39528
rect 28460 39528 29184 39556
rect 28460 39497 28488 39528
rect 29178 39516 29184 39528
rect 29236 39516 29242 39568
rect 29638 39556 29644 39568
rect 29599 39528 29644 39556
rect 29638 39516 29644 39528
rect 29696 39516 29702 39568
rect 29840 39565 29868 39596
rect 29825 39559 29883 39565
rect 29825 39525 29837 39559
rect 29871 39556 29883 39559
rect 30558 39556 30564 39568
rect 29871 39528 30564 39556
rect 29871 39525 29883 39528
rect 29825 39519 29883 39525
rect 30558 39516 30564 39528
rect 30616 39556 30622 39568
rect 30837 39559 30895 39565
rect 30837 39556 30849 39559
rect 30616 39528 30849 39556
rect 30616 39516 30622 39528
rect 30837 39525 30849 39528
rect 30883 39525 30895 39559
rect 30837 39519 30895 39525
rect 28261 39491 28319 39497
rect 28261 39457 28273 39491
rect 28307 39457 28319 39491
rect 28261 39451 28319 39457
rect 28445 39491 28503 39497
rect 28445 39457 28457 39491
rect 28491 39457 28503 39491
rect 28445 39451 28503 39457
rect 28166 39312 28172 39364
rect 28224 39352 28230 39364
rect 28276 39352 28304 39451
rect 28534 39448 28540 39500
rect 28592 39488 28598 39500
rect 28813 39491 28871 39497
rect 28592 39460 28637 39488
rect 28592 39448 28598 39460
rect 28813 39457 28825 39491
rect 28859 39488 28871 39491
rect 29086 39488 29092 39500
rect 28859 39460 29092 39488
rect 28859 39457 28871 39460
rect 28813 39451 28871 39457
rect 29086 39448 29092 39460
rect 29144 39448 29150 39500
rect 28626 39380 28632 39432
rect 28684 39420 28690 39432
rect 29914 39420 29920 39432
rect 28684 39392 29920 39420
rect 28684 39380 28690 39392
rect 29914 39380 29920 39392
rect 29972 39380 29978 39432
rect 29270 39352 29276 39364
rect 28224 39324 29276 39352
rect 28224 39312 28230 39324
rect 29270 39312 29276 39324
rect 29328 39312 29334 39364
rect 29086 39284 29092 39296
rect 28092 39256 29092 39284
rect 29086 39244 29092 39256
rect 29144 39284 29150 39296
rect 29457 39287 29515 39293
rect 29457 39284 29469 39287
rect 29144 39256 29469 39284
rect 29144 39244 29150 39256
rect 29457 39253 29469 39256
rect 29503 39253 29515 39287
rect 30374 39284 30380 39296
rect 30335 39256 30380 39284
rect 29457 39247 29515 39253
rect 30374 39244 30380 39256
rect 30432 39244 30438 39296
rect 1104 39194 32016 39216
rect 1104 39142 6102 39194
rect 6154 39142 6166 39194
rect 6218 39142 6230 39194
rect 6282 39142 6294 39194
rect 6346 39142 6358 39194
rect 6410 39142 16405 39194
rect 16457 39142 16469 39194
rect 16521 39142 16533 39194
rect 16585 39142 16597 39194
rect 16649 39142 16661 39194
rect 16713 39142 26709 39194
rect 26761 39142 26773 39194
rect 26825 39142 26837 39194
rect 26889 39142 26901 39194
rect 26953 39142 26965 39194
rect 27017 39142 32016 39194
rect 1104 39120 32016 39142
rect 5810 39080 5816 39092
rect 5771 39052 5816 39080
rect 5810 39040 5816 39052
rect 5868 39040 5874 39092
rect 6454 39040 6460 39092
rect 6512 39080 6518 39092
rect 6733 39083 6791 39089
rect 6733 39080 6745 39083
rect 6512 39052 6745 39080
rect 6512 39040 6518 39052
rect 6733 39049 6745 39052
rect 6779 39049 6791 39083
rect 6733 39043 6791 39049
rect 6822 39040 6828 39092
rect 6880 39080 6886 39092
rect 6917 39083 6975 39089
rect 6917 39080 6929 39083
rect 6880 39052 6929 39080
rect 6880 39040 6886 39052
rect 6917 39049 6929 39052
rect 6963 39080 6975 39083
rect 7374 39080 7380 39092
rect 6963 39052 7380 39080
rect 6963 39049 6975 39052
rect 6917 39043 6975 39049
rect 7374 39040 7380 39052
rect 7432 39040 7438 39092
rect 8386 39080 8392 39092
rect 8347 39052 8392 39080
rect 8386 39040 8392 39052
rect 8444 39040 8450 39092
rect 9033 39083 9091 39089
rect 9033 39049 9045 39083
rect 9079 39080 9091 39083
rect 9766 39080 9772 39092
rect 9079 39052 9772 39080
rect 9079 39049 9091 39052
rect 9033 39043 9091 39049
rect 9766 39040 9772 39052
rect 9824 39040 9830 39092
rect 14461 39083 14519 39089
rect 14461 39049 14473 39083
rect 14507 39080 14519 39083
rect 15654 39080 15660 39092
rect 14507 39052 15660 39080
rect 14507 39049 14519 39052
rect 14461 39043 14519 39049
rect 15654 39040 15660 39052
rect 15712 39040 15718 39092
rect 17957 39083 18015 39089
rect 17957 39049 17969 39083
rect 18003 39080 18015 39083
rect 18046 39080 18052 39092
rect 18003 39052 18052 39080
rect 18003 39049 18015 39052
rect 17957 39043 18015 39049
rect 18046 39040 18052 39052
rect 18104 39040 18110 39092
rect 19242 39080 19248 39092
rect 18340 39052 19248 39080
rect 5350 38972 5356 39024
rect 5408 39012 5414 39024
rect 6270 39012 6276 39024
rect 5408 38984 6276 39012
rect 5408 38972 5414 38984
rect 6270 38972 6276 38984
rect 6328 38972 6334 39024
rect 9858 39012 9864 39024
rect 9819 38984 9864 39012
rect 9858 38972 9864 38984
rect 9916 38972 9922 39024
rect 13078 39012 13084 39024
rect 12360 38984 13084 39012
rect 1394 38944 1400 38956
rect 1355 38916 1400 38944
rect 1394 38904 1400 38916
rect 1452 38904 1458 38956
rect 7929 38947 7987 38953
rect 7929 38913 7941 38947
rect 7975 38944 7987 38947
rect 8662 38944 8668 38956
rect 7975 38916 8668 38944
rect 7975 38913 7987 38916
rect 7929 38907 7987 38913
rect 8662 38904 8668 38916
rect 8720 38904 8726 38956
rect 12360 38953 12388 38984
rect 13078 38972 13084 38984
rect 13136 38972 13142 39024
rect 15286 39012 15292 39024
rect 15247 38984 15292 39012
rect 15286 38972 15292 38984
rect 15344 38972 15350 39024
rect 12345 38947 12403 38953
rect 12345 38913 12357 38947
rect 12391 38913 12403 38947
rect 12345 38907 12403 38913
rect 12434 38904 12440 38956
rect 12492 38944 12498 38956
rect 13265 38947 13323 38953
rect 13265 38944 13277 38947
rect 12492 38916 13277 38944
rect 12492 38904 12498 38916
rect 13265 38913 13277 38916
rect 13311 38913 13323 38947
rect 13265 38907 13323 38913
rect 14568 38916 15424 38944
rect 3786 38876 3792 38888
rect 2746 38848 3792 38876
rect 1664 38811 1722 38817
rect 1664 38777 1676 38811
rect 1710 38808 1722 38811
rect 1762 38808 1768 38820
rect 1710 38780 1768 38808
rect 1710 38777 1722 38780
rect 1664 38771 1722 38777
rect 1762 38768 1768 38780
rect 1820 38768 1826 38820
rect 2498 38768 2504 38820
rect 2556 38808 2562 38820
rect 2746 38808 2774 38848
rect 3786 38836 3792 38848
rect 3844 38836 3850 38888
rect 4154 38836 4160 38888
rect 4212 38876 4218 38888
rect 4525 38879 4583 38885
rect 4525 38876 4537 38879
rect 4212 38848 4537 38876
rect 4212 38836 4218 38848
rect 4525 38845 4537 38848
rect 4571 38845 4583 38879
rect 4525 38839 4583 38845
rect 7653 38879 7711 38885
rect 7653 38845 7665 38879
rect 7699 38845 7711 38879
rect 7834 38876 7840 38888
rect 7795 38848 7840 38876
rect 7653 38839 7711 38845
rect 2556 38780 2774 38808
rect 2556 38768 2562 38780
rect 3510 38768 3516 38820
rect 3568 38808 3574 38820
rect 4614 38808 4620 38820
rect 3568 38780 4620 38808
rect 3568 38768 3574 38780
rect 4614 38768 4620 38780
rect 4672 38768 4678 38820
rect 5626 38768 5632 38820
rect 5684 38808 5690 38820
rect 6885 38811 6943 38817
rect 6885 38808 6897 38811
rect 5684 38780 6897 38808
rect 5684 38768 5690 38780
rect 6885 38777 6897 38780
rect 6931 38777 6943 38811
rect 6885 38771 6943 38777
rect 7006 38768 7012 38820
rect 7064 38808 7070 38820
rect 7101 38811 7159 38817
rect 7101 38808 7113 38811
rect 7064 38780 7113 38808
rect 7064 38768 7070 38780
rect 7101 38777 7113 38780
rect 7147 38777 7159 38811
rect 7668 38808 7696 38839
rect 7834 38836 7840 38848
rect 7892 38836 7898 38888
rect 8021 38879 8079 38885
rect 8021 38845 8033 38879
rect 8067 38876 8079 38879
rect 8110 38876 8116 38888
rect 8067 38848 8116 38876
rect 8067 38845 8079 38848
rect 8021 38839 8079 38845
rect 8110 38836 8116 38848
rect 8168 38836 8174 38888
rect 8205 38879 8263 38885
rect 8205 38845 8217 38879
rect 8251 38876 8263 38879
rect 8938 38876 8944 38888
rect 8251 38848 8944 38876
rect 8251 38845 8263 38848
rect 8205 38839 8263 38845
rect 8938 38836 8944 38848
rect 8996 38836 9002 38888
rect 9217 38879 9275 38885
rect 9217 38845 9229 38879
rect 9263 38876 9275 38879
rect 10042 38876 10048 38888
rect 9263 38848 10048 38876
rect 9263 38845 9275 38848
rect 9217 38839 9275 38845
rect 10042 38836 10048 38848
rect 10100 38836 10106 38888
rect 12989 38879 13047 38885
rect 12989 38845 13001 38879
rect 13035 38845 13047 38879
rect 13170 38876 13176 38888
rect 13131 38848 13176 38876
rect 12989 38839 13047 38845
rect 9306 38808 9312 38820
rect 7668 38780 9312 38808
rect 7101 38771 7159 38777
rect 9306 38768 9312 38780
rect 9364 38768 9370 38820
rect 9401 38811 9459 38817
rect 9401 38777 9413 38811
rect 9447 38808 9459 38811
rect 9950 38808 9956 38820
rect 9447 38780 9956 38808
rect 9447 38777 9459 38780
rect 9401 38771 9459 38777
rect 9950 38768 9956 38780
rect 10008 38768 10014 38820
rect 10229 38811 10287 38817
rect 10229 38777 10241 38811
rect 10275 38808 10287 38811
rect 11146 38808 11152 38820
rect 10275 38780 11152 38808
rect 10275 38777 10287 38780
rect 10229 38771 10287 38777
rect 11146 38768 11152 38780
rect 11204 38768 11210 38820
rect 12100 38811 12158 38817
rect 12100 38777 12112 38811
rect 12146 38808 12158 38811
rect 12805 38811 12863 38817
rect 12805 38808 12817 38811
rect 12146 38780 12817 38808
rect 12146 38777 12158 38780
rect 12100 38771 12158 38777
rect 12805 38777 12817 38780
rect 12851 38777 12863 38811
rect 12805 38771 12863 38777
rect 2222 38700 2228 38752
rect 2280 38740 2286 38752
rect 2777 38743 2835 38749
rect 2777 38740 2789 38743
rect 2280 38712 2789 38740
rect 2280 38700 2286 38712
rect 2777 38709 2789 38712
rect 2823 38709 2835 38743
rect 2777 38703 2835 38709
rect 10965 38743 11023 38749
rect 10965 38709 10977 38743
rect 11011 38740 11023 38743
rect 11790 38740 11796 38752
rect 11011 38712 11796 38740
rect 11011 38709 11023 38712
rect 10965 38703 11023 38709
rect 11790 38700 11796 38712
rect 11848 38740 11854 38752
rect 13004 38740 13032 38839
rect 13170 38836 13176 38848
rect 13228 38836 13234 38888
rect 13354 38836 13360 38888
rect 13412 38876 13418 38888
rect 14568 38885 14596 38916
rect 15396 38888 15424 38916
rect 15562 38904 15568 38956
rect 15620 38944 15626 38956
rect 16485 38947 16543 38953
rect 16485 38944 16497 38947
rect 15620 38916 16497 38944
rect 15620 38904 15626 38916
rect 16485 38913 16497 38916
rect 16531 38913 16543 38947
rect 16485 38907 16543 38913
rect 16761 38947 16819 38953
rect 16761 38913 16773 38947
rect 16807 38944 16819 38947
rect 16850 38944 16856 38956
rect 16807 38916 16856 38944
rect 16807 38913 16819 38916
rect 16761 38907 16819 38913
rect 16850 38904 16856 38916
rect 16908 38944 16914 38956
rect 17494 38944 17500 38956
rect 16908 38916 17500 38944
rect 16908 38904 16914 38916
rect 17494 38904 17500 38916
rect 17552 38904 17558 38956
rect 18340 38944 18368 39052
rect 19242 39040 19248 39052
rect 19300 39040 19306 39092
rect 20530 39080 20536 39092
rect 20491 39052 20536 39080
rect 20530 39040 20536 39052
rect 20588 39040 20594 39092
rect 22278 39080 22284 39092
rect 22239 39052 22284 39080
rect 22278 39040 22284 39052
rect 22336 39040 22342 39092
rect 23382 39040 23388 39092
rect 23440 39080 23446 39092
rect 25314 39080 25320 39092
rect 23440 39052 25320 39080
rect 23440 39040 23446 39052
rect 25314 39040 25320 39052
rect 25372 39040 25378 39092
rect 25774 39040 25780 39092
rect 25832 39080 25838 39092
rect 26510 39080 26516 39092
rect 25832 39052 26516 39080
rect 25832 39040 25838 39052
rect 26510 39040 26516 39052
rect 26568 39080 26574 39092
rect 26697 39083 26755 39089
rect 26697 39080 26709 39083
rect 26568 39052 26709 39080
rect 26568 39040 26574 39052
rect 26697 39049 26709 39052
rect 26743 39049 26755 39083
rect 26697 39043 26755 39049
rect 27157 39083 27215 39089
rect 27157 39049 27169 39083
rect 27203 39080 27215 39083
rect 27706 39080 27712 39092
rect 27203 39052 27712 39080
rect 27203 39049 27215 39052
rect 27157 39043 27215 39049
rect 27706 39040 27712 39052
rect 27764 39040 27770 39092
rect 29733 39083 29791 39089
rect 29733 39049 29745 39083
rect 29779 39080 29791 39083
rect 29914 39080 29920 39092
rect 29779 39052 29920 39080
rect 29779 39049 29791 39052
rect 29733 39043 29791 39049
rect 29914 39040 29920 39052
rect 29972 39040 29978 39092
rect 31294 39080 31300 39092
rect 31255 39052 31300 39080
rect 31294 39040 31300 39052
rect 31352 39040 31358 39092
rect 19794 39012 19800 39024
rect 18432 38984 19800 39012
rect 18432 38953 18460 38984
rect 19794 38972 19800 38984
rect 19852 39012 19858 39024
rect 20438 39012 20444 39024
rect 19852 38984 20444 39012
rect 19852 38972 19858 38984
rect 20438 38972 20444 38984
rect 20496 39012 20502 39024
rect 20496 38984 21036 39012
rect 20496 38972 20502 38984
rect 18156 38916 18368 38944
rect 18417 38947 18475 38953
rect 13541 38879 13599 38885
rect 13412 38848 13457 38876
rect 13412 38836 13418 38848
rect 13541 38845 13553 38879
rect 13587 38845 13599 38879
rect 13541 38839 13599 38845
rect 14553 38879 14611 38885
rect 14553 38845 14565 38879
rect 14599 38845 14611 38879
rect 14553 38839 14611 38845
rect 15013 38879 15071 38885
rect 15013 38845 15025 38879
rect 15059 38845 15071 38879
rect 15194 38876 15200 38888
rect 15155 38848 15200 38876
rect 15013 38839 15071 38845
rect 13446 38768 13452 38820
rect 13504 38808 13510 38820
rect 13556 38808 13584 38839
rect 13504 38780 13584 38808
rect 15028 38808 15056 38839
rect 15194 38836 15200 38848
rect 15252 38836 15258 38888
rect 15378 38876 15384 38888
rect 15339 38848 15384 38876
rect 15378 38836 15384 38848
rect 15436 38836 15442 38888
rect 15470 38836 15476 38888
rect 15528 38876 15534 38888
rect 18156 38885 18184 38916
rect 18417 38913 18429 38947
rect 18463 38913 18475 38947
rect 20898 38944 20904 38956
rect 18417 38907 18475 38913
rect 18524 38916 20760 38944
rect 20859 38916 20904 38944
rect 18524 38888 18552 38916
rect 18141 38879 18199 38885
rect 15528 38848 15573 38876
rect 15528 38836 15534 38848
rect 18141 38845 18153 38879
rect 18187 38845 18199 38879
rect 18141 38839 18199 38845
rect 18325 38879 18383 38885
rect 18325 38845 18337 38879
rect 18371 38845 18383 38879
rect 18325 38839 18383 38845
rect 15286 38808 15292 38820
rect 15028 38780 15292 38808
rect 13504 38768 13510 38780
rect 15286 38768 15292 38780
rect 15344 38768 15350 38820
rect 16206 38768 16212 38820
rect 16264 38808 16270 38820
rect 17862 38808 17868 38820
rect 16264 38780 17868 38808
rect 16264 38768 16270 38780
rect 17862 38768 17868 38780
rect 17920 38768 17926 38820
rect 11848 38712 13032 38740
rect 15657 38743 15715 38749
rect 11848 38700 11854 38712
rect 15657 38709 15669 38743
rect 15703 38740 15715 38743
rect 16850 38740 16856 38752
rect 15703 38712 16856 38740
rect 15703 38709 15715 38712
rect 15657 38703 15715 38709
rect 16850 38700 16856 38712
rect 16908 38700 16914 38752
rect 18340 38740 18368 38839
rect 18506 38836 18512 38888
rect 18564 38876 18570 38888
rect 18693 38879 18751 38885
rect 18564 38848 18609 38876
rect 18564 38836 18570 38848
rect 18693 38845 18705 38879
rect 18739 38876 18751 38879
rect 19426 38876 19432 38888
rect 18739 38848 19432 38876
rect 18739 38845 18751 38848
rect 18693 38839 18751 38845
rect 19426 38836 19432 38848
rect 19484 38876 19490 38888
rect 19797 38879 19855 38885
rect 19484 38848 19748 38876
rect 19484 38836 19490 38848
rect 19720 38808 19748 38848
rect 19797 38845 19809 38879
rect 19843 38876 19855 38879
rect 19978 38876 19984 38888
rect 19843 38848 19984 38876
rect 19843 38845 19855 38848
rect 19797 38839 19855 38845
rect 19978 38836 19984 38848
rect 20036 38836 20042 38888
rect 20073 38879 20131 38885
rect 20073 38845 20085 38879
rect 20119 38876 20131 38879
rect 20530 38876 20536 38888
rect 20119 38848 20536 38876
rect 20119 38845 20131 38848
rect 20073 38839 20131 38845
rect 20530 38836 20536 38848
rect 20588 38836 20594 38888
rect 20732 38885 20760 38916
rect 20898 38904 20904 38916
rect 20956 38904 20962 38956
rect 21008 38953 21036 38984
rect 21358 38972 21364 39024
rect 21416 39012 21422 39024
rect 24578 39012 24584 39024
rect 21416 38984 24584 39012
rect 21416 38972 21422 38984
rect 24578 38972 24584 38984
rect 24636 39012 24642 39024
rect 25406 39012 25412 39024
rect 24636 38984 25412 39012
rect 24636 38972 24642 38984
rect 25406 38972 25412 38984
rect 25464 38972 25470 39024
rect 28442 39012 28448 39024
rect 26252 38984 28448 39012
rect 20993 38947 21051 38953
rect 20993 38913 21005 38947
rect 21039 38913 21051 38947
rect 20993 38907 21051 38913
rect 23198 38904 23204 38956
rect 23256 38944 23262 38956
rect 23382 38944 23388 38956
rect 23256 38916 23388 38944
rect 23256 38904 23262 38916
rect 23382 38904 23388 38916
rect 23440 38904 23446 38956
rect 23474 38904 23480 38956
rect 23532 38944 23538 38956
rect 24762 38944 24768 38956
rect 23532 38916 24768 38944
rect 23532 38904 23538 38916
rect 24762 38904 24768 38916
rect 24820 38944 24826 38956
rect 25041 38947 25099 38953
rect 25041 38944 25053 38947
rect 24820 38916 25053 38944
rect 24820 38904 24826 38916
rect 25041 38913 25053 38916
rect 25087 38913 25099 38947
rect 25041 38907 25099 38913
rect 26252 38888 26280 38984
rect 28442 38972 28448 38984
rect 28500 39012 28506 39024
rect 28905 39015 28963 39021
rect 28905 39012 28917 39015
rect 28500 38984 28917 39012
rect 28500 38972 28506 38984
rect 28905 38981 28917 38984
rect 28951 39012 28963 39015
rect 30374 39012 30380 39024
rect 28951 38984 30380 39012
rect 28951 38981 28963 38984
rect 28905 38975 28963 38981
rect 30374 38972 30380 38984
rect 30432 39012 30438 39024
rect 31110 39012 31116 39024
rect 30432 38984 31116 39012
rect 30432 38972 30438 38984
rect 31110 38972 31116 38984
rect 31168 38972 31174 39024
rect 27798 38904 27804 38956
rect 27856 38944 27862 38956
rect 28077 38947 28135 38953
rect 28077 38944 28089 38947
rect 27856 38916 28089 38944
rect 27856 38904 27862 38916
rect 28077 38913 28089 38916
rect 28123 38913 28135 38947
rect 28077 38907 28135 38913
rect 20717 38879 20775 38885
rect 20717 38845 20729 38879
rect 20763 38845 20775 38879
rect 20717 38839 20775 38845
rect 21085 38879 21143 38885
rect 21085 38845 21097 38879
rect 21131 38876 21143 38879
rect 21174 38876 21180 38888
rect 21131 38848 21180 38876
rect 21131 38845 21143 38848
rect 21085 38839 21143 38845
rect 21174 38836 21180 38848
rect 21232 38836 21238 38888
rect 21269 38879 21327 38885
rect 21269 38845 21281 38879
rect 21315 38845 21327 38879
rect 22370 38876 22376 38888
rect 22331 38848 22376 38876
rect 21269 38839 21327 38845
rect 20346 38808 20352 38820
rect 19720 38780 20352 38808
rect 20346 38768 20352 38780
rect 20404 38808 20410 38820
rect 21284 38808 21312 38839
rect 22370 38836 22376 38848
rect 22428 38836 22434 38888
rect 23106 38876 23112 38888
rect 23067 38848 23112 38876
rect 23106 38836 23112 38848
rect 23164 38836 23170 38888
rect 23290 38876 23296 38888
rect 23251 38848 23296 38876
rect 23290 38836 23296 38848
rect 23348 38836 23354 38888
rect 23566 38836 23572 38888
rect 23624 38876 23630 38888
rect 23661 38879 23719 38885
rect 23661 38876 23673 38879
rect 23624 38848 23673 38876
rect 23624 38836 23630 38848
rect 23661 38845 23673 38848
rect 23707 38845 23719 38879
rect 25961 38879 26019 38885
rect 25961 38876 25973 38879
rect 23661 38839 23719 38845
rect 24504 38848 25973 38876
rect 24504 38808 24532 38848
rect 25961 38845 25973 38848
rect 26007 38876 26019 38879
rect 26234 38876 26240 38888
rect 26007 38848 26240 38876
rect 26007 38845 26019 38848
rect 25961 38839 26019 38845
rect 26234 38836 26240 38848
rect 26292 38836 26298 38888
rect 26602 38876 26608 38888
rect 26563 38848 26608 38876
rect 26602 38836 26608 38848
rect 26660 38836 26666 38888
rect 26973 38879 27031 38885
rect 26973 38845 26985 38879
rect 27019 38876 27031 38879
rect 27522 38876 27528 38888
rect 27019 38848 27528 38876
rect 27019 38845 27031 38848
rect 26973 38839 27031 38845
rect 27522 38836 27528 38848
rect 27580 38836 27586 38888
rect 27614 38836 27620 38888
rect 27672 38876 27678 38888
rect 27709 38879 27767 38885
rect 27709 38876 27721 38879
rect 27672 38848 27721 38876
rect 27672 38836 27678 38848
rect 27709 38845 27721 38848
rect 27755 38845 27767 38879
rect 27890 38876 27896 38888
rect 27851 38848 27896 38876
rect 27709 38839 27767 38845
rect 27890 38836 27896 38848
rect 27948 38836 27954 38888
rect 27982 38836 27988 38888
rect 28040 38876 28046 38888
rect 28258 38876 28264 38888
rect 28040 38848 28085 38876
rect 28219 38848 28264 38876
rect 28040 38836 28046 38848
rect 28258 38836 28264 38848
rect 28316 38836 28322 38888
rect 30466 38876 30472 38888
rect 30427 38848 30472 38876
rect 30466 38836 30472 38848
rect 30524 38836 30530 38888
rect 31018 38836 31024 38888
rect 31076 38876 31082 38888
rect 31113 38879 31171 38885
rect 31113 38876 31125 38879
rect 31076 38848 31125 38876
rect 31076 38836 31082 38848
rect 31113 38845 31125 38848
rect 31159 38845 31171 38879
rect 31113 38839 31171 38845
rect 20404 38780 21312 38808
rect 23676 38780 24532 38808
rect 24857 38811 24915 38817
rect 20404 38768 20410 38780
rect 23676 38752 23704 38780
rect 24857 38777 24869 38811
rect 24903 38808 24915 38811
rect 24903 38780 25728 38808
rect 24903 38777 24915 38780
rect 24857 38771 24915 38777
rect 19702 38740 19708 38752
rect 18340 38712 19708 38740
rect 19702 38700 19708 38712
rect 19760 38740 19766 38752
rect 20898 38740 20904 38752
rect 19760 38712 20904 38740
rect 19760 38700 19766 38712
rect 20898 38700 20904 38712
rect 20956 38700 20962 38752
rect 22002 38700 22008 38752
rect 22060 38740 22066 38752
rect 22278 38740 22284 38752
rect 22060 38712 22284 38740
rect 22060 38700 22066 38712
rect 22278 38700 22284 38712
rect 22336 38700 22342 38752
rect 23658 38700 23664 38752
rect 23716 38700 23722 38752
rect 23842 38740 23848 38752
rect 23803 38712 23848 38740
rect 23842 38700 23848 38712
rect 23900 38700 23906 38752
rect 24302 38700 24308 38752
rect 24360 38740 24366 38752
rect 25038 38740 25044 38752
rect 24360 38712 25044 38740
rect 24360 38700 24366 38712
rect 25038 38700 25044 38712
rect 25096 38700 25102 38752
rect 25700 38740 25728 38780
rect 25774 38768 25780 38820
rect 25832 38808 25838 38820
rect 26145 38811 26203 38817
rect 25832 38780 25877 38808
rect 25832 38768 25838 38780
rect 26145 38777 26157 38811
rect 26191 38808 26203 38811
rect 28000 38808 28028 38836
rect 29641 38811 29699 38817
rect 29641 38808 29653 38811
rect 26191 38780 28028 38808
rect 28092 38780 29653 38808
rect 26191 38777 26203 38780
rect 26145 38771 26203 38777
rect 26418 38740 26424 38752
rect 25700 38712 26424 38740
rect 26418 38700 26424 38712
rect 26476 38740 26482 38752
rect 28092 38740 28120 38780
rect 29641 38777 29653 38780
rect 29687 38777 29699 38811
rect 29641 38771 29699 38777
rect 28442 38740 28448 38752
rect 26476 38712 28120 38740
rect 28403 38712 28448 38740
rect 26476 38700 26482 38712
rect 28442 38700 28448 38712
rect 28500 38700 28506 38752
rect 30374 38740 30380 38752
rect 30335 38712 30380 38740
rect 30374 38700 30380 38712
rect 30432 38700 30438 38752
rect 1104 38650 32016 38672
rect 1104 38598 11253 38650
rect 11305 38598 11317 38650
rect 11369 38598 11381 38650
rect 11433 38598 11445 38650
rect 11497 38598 11509 38650
rect 11561 38598 21557 38650
rect 21609 38598 21621 38650
rect 21673 38598 21685 38650
rect 21737 38598 21749 38650
rect 21801 38598 21813 38650
rect 21865 38598 32016 38650
rect 1104 38576 32016 38598
rect 1762 38536 1768 38548
rect 1723 38508 1768 38536
rect 1762 38496 1768 38508
rect 1820 38496 1826 38548
rect 2222 38536 2228 38548
rect 1964 38508 2228 38536
rect 1762 38360 1768 38412
rect 1820 38400 1826 38412
rect 1964 38409 1992 38508
rect 2222 38496 2228 38508
rect 2280 38496 2286 38548
rect 2498 38496 2504 38548
rect 2556 38496 2562 38548
rect 4338 38536 4344 38548
rect 4080 38508 4344 38536
rect 2516 38468 2544 38496
rect 2240 38440 2544 38468
rect 2240 38409 2268 38440
rect 1949 38403 2007 38409
rect 1949 38400 1961 38403
rect 1820 38372 1961 38400
rect 1820 38360 1826 38372
rect 1949 38369 1961 38372
rect 1995 38369 2007 38403
rect 1949 38363 2007 38369
rect 2225 38403 2283 38409
rect 2225 38369 2237 38403
rect 2271 38369 2283 38403
rect 2225 38363 2283 38369
rect 2317 38403 2375 38409
rect 2317 38369 2329 38403
rect 2363 38369 2375 38403
rect 2317 38363 2375 38369
rect 2130 38332 2136 38344
rect 2091 38304 2136 38332
rect 2130 38292 2136 38304
rect 2188 38292 2194 38344
rect 2332 38332 2360 38363
rect 2406 38360 2412 38412
rect 2464 38400 2470 38412
rect 2501 38403 2559 38409
rect 2501 38400 2513 38403
rect 2464 38372 2513 38400
rect 2464 38360 2470 38372
rect 2501 38369 2513 38372
rect 2547 38369 2559 38403
rect 2501 38363 2559 38369
rect 3142 38360 3148 38412
rect 3200 38400 3206 38412
rect 3237 38403 3295 38409
rect 3237 38400 3249 38403
rect 3200 38372 3249 38400
rect 3200 38360 3206 38372
rect 3237 38369 3249 38372
rect 3283 38369 3295 38403
rect 3878 38400 3884 38412
rect 3839 38372 3884 38400
rect 3237 38363 3295 38369
rect 3878 38360 3884 38372
rect 3936 38360 3942 38412
rect 4080 38409 4108 38508
rect 4338 38496 4344 38508
rect 4396 38496 4402 38548
rect 5261 38539 5319 38545
rect 5261 38505 5273 38539
rect 5307 38536 5319 38539
rect 7190 38536 7196 38548
rect 5307 38508 7196 38536
rect 5307 38505 5319 38508
rect 5261 38499 5319 38505
rect 7190 38496 7196 38508
rect 7248 38496 7254 38548
rect 7834 38496 7840 38548
rect 7892 38536 7898 38548
rect 8113 38539 8171 38545
rect 8113 38536 8125 38539
rect 7892 38508 8125 38536
rect 7892 38496 7898 38508
rect 8113 38505 8125 38508
rect 8159 38505 8171 38539
rect 8113 38499 8171 38505
rect 4246 38468 4252 38480
rect 4172 38440 4252 38468
rect 4172 38409 4200 38440
rect 4246 38428 4252 38440
rect 4304 38428 4310 38480
rect 6914 38468 6920 38480
rect 5552 38440 6920 38468
rect 5552 38412 5580 38440
rect 6914 38428 6920 38440
rect 6972 38428 6978 38480
rect 8128 38468 8156 38499
rect 8662 38496 8668 38548
rect 8720 38536 8726 38548
rect 8720 38508 9076 38536
rect 8720 38496 8726 38508
rect 9048 38468 9076 38508
rect 9674 38496 9680 38548
rect 9732 38536 9738 38548
rect 9769 38539 9827 38545
rect 9769 38536 9781 38539
rect 9732 38508 9781 38536
rect 9732 38496 9738 38508
rect 9769 38505 9781 38508
rect 9815 38505 9827 38539
rect 9769 38499 9827 38505
rect 11146 38496 11152 38548
rect 11204 38536 11210 38548
rect 11609 38539 11667 38545
rect 11609 38536 11621 38539
rect 11204 38508 11621 38536
rect 11204 38496 11210 38508
rect 11609 38505 11621 38508
rect 11655 38505 11667 38539
rect 12526 38536 12532 38548
rect 11609 38499 11667 38505
rect 12406 38508 12532 38536
rect 9214 38468 9220 38480
rect 8128 38440 8800 38468
rect 4065 38403 4123 38409
rect 4065 38369 4077 38403
rect 4111 38369 4123 38403
rect 4065 38363 4123 38369
rect 4157 38403 4215 38409
rect 4157 38369 4169 38403
rect 4203 38369 4215 38403
rect 4157 38363 4215 38369
rect 4433 38403 4491 38409
rect 4433 38369 4445 38403
rect 4479 38400 4491 38403
rect 5534 38400 5540 38412
rect 4479 38372 5396 38400
rect 5495 38372 5540 38400
rect 4479 38369 4491 38372
rect 4433 38363 4491 38369
rect 2590 38332 2596 38344
rect 2332 38304 2596 38332
rect 2590 38292 2596 38304
rect 2648 38292 2654 38344
rect 4249 38335 4307 38341
rect 4249 38301 4261 38335
rect 4295 38332 4307 38335
rect 5258 38332 5264 38344
rect 4295 38304 4568 38332
rect 5219 38304 5264 38332
rect 4295 38301 4307 38304
rect 4249 38295 4307 38301
rect 3329 38267 3387 38273
rect 3329 38233 3341 38267
rect 3375 38264 3387 38267
rect 4430 38264 4436 38276
rect 3375 38236 4436 38264
rect 3375 38233 3387 38236
rect 3329 38227 3387 38233
rect 4430 38224 4436 38236
rect 4488 38224 4494 38276
rect 4154 38156 4160 38208
rect 4212 38196 4218 38208
rect 4540 38196 4568 38304
rect 5258 38292 5264 38304
rect 5316 38292 5322 38344
rect 5368 38332 5396 38372
rect 5534 38360 5540 38372
rect 5592 38360 5598 38412
rect 5810 38360 5816 38412
rect 5868 38400 5874 38412
rect 6638 38400 6644 38412
rect 5868 38372 6644 38400
rect 5868 38360 5874 38372
rect 6638 38360 6644 38372
rect 6696 38400 6702 38412
rect 8772 38409 8800 38440
rect 9048 38440 9220 38468
rect 9048 38409 9076 38440
rect 9214 38428 9220 38440
rect 9272 38428 9278 38480
rect 10873 38471 10931 38477
rect 10873 38468 10885 38471
rect 10060 38440 10885 38468
rect 10060 38412 10088 38440
rect 10873 38437 10885 38440
rect 10919 38437 10931 38471
rect 12406 38468 12434 38508
rect 12526 38496 12532 38508
rect 12584 38536 12590 38548
rect 13446 38536 13452 38548
rect 12584 38508 13452 38536
rect 12584 38496 12590 38508
rect 13446 38496 13452 38508
rect 13504 38496 13510 38548
rect 14642 38496 14648 38548
rect 14700 38536 14706 38548
rect 14737 38539 14795 38545
rect 14737 38536 14749 38539
rect 14700 38508 14749 38536
rect 14700 38496 14706 38508
rect 14737 38505 14749 38508
rect 14783 38536 14795 38539
rect 15565 38539 15623 38545
rect 15565 38536 15577 38539
rect 14783 38508 15577 38536
rect 14783 38505 14795 38508
rect 14737 38499 14795 38505
rect 15565 38505 15577 38508
rect 15611 38505 15623 38539
rect 15565 38499 15623 38505
rect 16025 38539 16083 38545
rect 16025 38505 16037 38539
rect 16071 38536 16083 38539
rect 16827 38539 16885 38545
rect 16827 38536 16839 38539
rect 16071 38508 16839 38536
rect 16071 38505 16083 38508
rect 16025 38499 16083 38505
rect 16827 38505 16839 38508
rect 16873 38505 16885 38539
rect 16827 38499 16885 38505
rect 17402 38496 17408 38548
rect 17460 38536 17466 38548
rect 17460 38508 17816 38536
rect 17460 38496 17466 38508
rect 10873 38431 10931 38437
rect 12176 38440 12434 38468
rect 12897 38471 12955 38477
rect 6733 38403 6791 38409
rect 6733 38400 6745 38403
rect 6696 38372 6745 38400
rect 6696 38360 6702 38372
rect 6733 38369 6745 38372
rect 6779 38369 6791 38403
rect 6733 38363 6791 38369
rect 7000 38403 7058 38409
rect 7000 38369 7012 38403
rect 7046 38400 7058 38403
rect 8573 38403 8631 38409
rect 8573 38400 8585 38403
rect 7046 38372 8585 38400
rect 7046 38369 7058 38372
rect 7000 38363 7058 38369
rect 8573 38369 8585 38372
rect 8619 38369 8631 38403
rect 8573 38363 8631 38369
rect 8757 38403 8815 38409
rect 8757 38369 8769 38403
rect 8803 38369 8815 38403
rect 8757 38363 8815 38369
rect 9033 38403 9091 38409
rect 9033 38369 9045 38403
rect 9079 38369 9091 38403
rect 9033 38363 9091 38369
rect 9122 38360 9128 38412
rect 9180 38400 9186 38412
rect 9180 38372 9273 38400
rect 9180 38360 9186 38372
rect 5718 38332 5724 38344
rect 5368 38304 5724 38332
rect 5718 38292 5724 38304
rect 5776 38292 5782 38344
rect 8110 38292 8116 38344
rect 8168 38332 8174 38344
rect 8846 38332 8852 38344
rect 8168 38304 8852 38332
rect 8168 38292 8174 38304
rect 8846 38292 8852 38304
rect 8904 38332 8910 38344
rect 8941 38335 8999 38341
rect 8941 38332 8953 38335
rect 8904 38304 8953 38332
rect 8904 38292 8910 38304
rect 8941 38301 8953 38304
rect 8987 38301 8999 38335
rect 9226 38332 9254 38372
rect 9306 38360 9312 38412
rect 9364 38400 9370 38412
rect 10042 38400 10048 38412
rect 9364 38372 9409 38400
rect 10003 38372 10048 38400
rect 9364 38360 9370 38372
rect 10042 38360 10048 38372
rect 10100 38360 10106 38412
rect 10321 38403 10379 38409
rect 10321 38369 10333 38403
rect 10367 38369 10379 38403
rect 10321 38363 10379 38369
rect 10336 38332 10364 38363
rect 10410 38360 10416 38412
rect 10468 38400 10474 38412
rect 10962 38400 10968 38412
rect 10468 38372 10968 38400
rect 10468 38360 10474 38372
rect 10962 38360 10968 38372
rect 11020 38360 11026 38412
rect 11517 38403 11575 38409
rect 11517 38369 11529 38403
rect 11563 38369 11575 38403
rect 11517 38363 11575 38369
rect 9226 38304 10364 38332
rect 8941 38295 8999 38301
rect 4890 38224 4896 38276
rect 4948 38264 4954 38276
rect 5350 38264 5356 38276
rect 4948 38236 5356 38264
rect 4948 38224 4954 38236
rect 5350 38224 5356 38236
rect 5408 38264 5414 38276
rect 5445 38267 5503 38273
rect 5445 38264 5457 38267
rect 5408 38236 5457 38264
rect 5408 38224 5414 38236
rect 5445 38233 5457 38236
rect 5491 38233 5503 38267
rect 8956 38264 8984 38295
rect 9582 38264 9588 38276
rect 8956 38236 9588 38264
rect 5445 38227 5503 38233
rect 4212 38168 4568 38196
rect 4617 38199 4675 38205
rect 4212 38156 4218 38168
rect 4617 38165 4629 38199
rect 4663 38196 4675 38199
rect 4706 38196 4712 38208
rect 4663 38168 4712 38196
rect 4663 38165 4675 38168
rect 4617 38159 4675 38165
rect 4706 38156 4712 38168
rect 4764 38156 4770 38208
rect 5460 38196 5488 38227
rect 9582 38224 9588 38236
rect 9640 38224 9646 38276
rect 11532 38264 11560 38363
rect 11698 38360 11704 38412
rect 11756 38400 11762 38412
rect 12176 38409 12204 38440
rect 12897 38437 12909 38471
rect 12943 38468 12955 38471
rect 13602 38471 13660 38477
rect 13602 38468 13614 38471
rect 12943 38440 13614 38468
rect 12943 38437 12955 38440
rect 12897 38431 12955 38437
rect 13602 38437 13614 38440
rect 13648 38437 13660 38471
rect 13602 38431 13660 38437
rect 12161 38403 12219 38409
rect 12161 38400 12173 38403
rect 11756 38372 12173 38400
rect 11756 38360 11762 38372
rect 12161 38369 12173 38372
rect 12207 38369 12219 38403
rect 12161 38363 12219 38369
rect 12345 38403 12403 38409
rect 12345 38369 12357 38403
rect 12391 38369 12403 38403
rect 12345 38363 12403 38369
rect 12529 38403 12587 38409
rect 12529 38369 12541 38403
rect 12575 38400 12587 38403
rect 12618 38400 12624 38412
rect 12575 38372 12624 38400
rect 12575 38369 12587 38372
rect 12529 38363 12587 38369
rect 10060 38236 11560 38264
rect 10060 38208 10088 38236
rect 7650 38196 7656 38208
rect 5460 38168 7656 38196
rect 7650 38156 7656 38168
rect 7708 38156 7714 38208
rect 10042 38196 10048 38208
rect 10003 38168 10048 38196
rect 10042 38156 10048 38168
rect 10100 38156 10106 38208
rect 12360 38196 12388 38363
rect 12618 38360 12624 38372
rect 12676 38360 12682 38412
rect 12713 38403 12771 38409
rect 12713 38369 12725 38403
rect 12759 38400 12771 38403
rect 14660 38400 14688 38496
rect 15657 38471 15715 38477
rect 15657 38437 15669 38471
rect 15703 38468 15715 38471
rect 16942 38468 16948 38480
rect 15703 38440 16948 38468
rect 15703 38437 15715 38440
rect 15657 38431 15715 38437
rect 16942 38428 16948 38440
rect 17000 38428 17006 38480
rect 17037 38471 17095 38477
rect 17037 38437 17049 38471
rect 17083 38468 17095 38471
rect 17310 38468 17316 38480
rect 17083 38440 17316 38468
rect 17083 38437 17095 38440
rect 17037 38431 17095 38437
rect 17310 38428 17316 38440
rect 17368 38468 17374 38480
rect 17368 38440 17724 38468
rect 17368 38428 17374 38440
rect 12759 38372 14688 38400
rect 12759 38369 12771 38372
rect 12713 38363 12771 38369
rect 16666 38360 16672 38412
rect 16724 38400 16730 38412
rect 17218 38400 17224 38412
rect 16724 38372 17224 38400
rect 16724 38360 16730 38372
rect 17218 38360 17224 38372
rect 17276 38360 17282 38412
rect 17494 38400 17500 38412
rect 17455 38372 17500 38400
rect 17494 38360 17500 38372
rect 17552 38360 17558 38412
rect 17696 38409 17724 38440
rect 17681 38403 17739 38409
rect 17681 38369 17693 38403
rect 17727 38369 17739 38403
rect 17788 38400 17816 38508
rect 17862 38496 17868 38548
rect 17920 38496 17926 38548
rect 18230 38536 18236 38548
rect 18191 38508 18236 38536
rect 18230 38496 18236 38508
rect 18288 38496 18294 38548
rect 19058 38496 19064 38548
rect 19116 38536 19122 38548
rect 20346 38536 20352 38548
rect 19116 38508 20352 38536
rect 19116 38496 19122 38508
rect 20346 38496 20352 38508
rect 20404 38496 20410 38548
rect 22002 38496 22008 38548
rect 22060 38536 22066 38548
rect 22060 38508 23060 38536
rect 22060 38496 22066 38508
rect 17880 38468 17908 38496
rect 22738 38468 22744 38480
rect 17880 38440 18920 38468
rect 17865 38403 17923 38409
rect 17865 38400 17877 38403
rect 17788 38372 17877 38400
rect 17681 38363 17739 38369
rect 17865 38369 17877 38372
rect 17911 38369 17923 38403
rect 17865 38363 17923 38369
rect 18049 38403 18107 38409
rect 18049 38369 18061 38403
rect 18095 38400 18107 38403
rect 18138 38400 18144 38412
rect 18095 38372 18144 38400
rect 18095 38369 18107 38372
rect 18049 38363 18107 38369
rect 18138 38360 18144 38372
rect 18196 38360 18202 38412
rect 18690 38400 18696 38412
rect 18651 38372 18696 38400
rect 18690 38360 18696 38372
rect 18748 38360 18754 38412
rect 18892 38409 18920 38440
rect 19306 38440 22744 38468
rect 18877 38403 18935 38409
rect 18877 38369 18889 38403
rect 18923 38369 18935 38403
rect 18877 38363 18935 38369
rect 12434 38292 12440 38344
rect 12492 38332 12498 38344
rect 12492 38304 12537 38332
rect 12492 38292 12498 38304
rect 13078 38292 13084 38344
rect 13136 38332 13142 38344
rect 13357 38335 13415 38341
rect 13357 38332 13369 38335
rect 13136 38304 13369 38332
rect 13136 38292 13142 38304
rect 13357 38301 13369 38304
rect 13403 38301 13415 38335
rect 13357 38295 13415 38301
rect 15473 38335 15531 38341
rect 15473 38301 15485 38335
rect 15519 38332 15531 38335
rect 17770 38332 17776 38344
rect 15519 38304 17080 38332
rect 17731 38304 17776 38332
rect 15519 38301 15531 38304
rect 15473 38295 15531 38301
rect 16666 38264 16672 38276
rect 16627 38236 16672 38264
rect 16666 38224 16672 38236
rect 16724 38224 16730 38276
rect 17052 38264 17080 38304
rect 17770 38292 17776 38304
rect 17828 38292 17834 38344
rect 18693 38267 18751 38273
rect 18693 38264 18705 38267
rect 17052 38236 18705 38264
rect 18693 38233 18705 38236
rect 18739 38233 18751 38267
rect 18693 38227 18751 38233
rect 16298 38196 16304 38208
rect 12360 38168 16304 38196
rect 16298 38156 16304 38168
rect 16356 38156 16362 38208
rect 16853 38199 16911 38205
rect 16853 38165 16865 38199
rect 16899 38196 16911 38199
rect 16942 38196 16948 38208
rect 16899 38168 16948 38196
rect 16899 38165 16911 38168
rect 16853 38159 16911 38165
rect 16942 38156 16948 38168
rect 17000 38196 17006 38208
rect 19306 38196 19334 38440
rect 22738 38428 22744 38440
rect 22796 38428 22802 38480
rect 23032 38468 23060 38508
rect 23106 38496 23112 38548
rect 23164 38536 23170 38548
rect 24210 38536 24216 38548
rect 23164 38508 24216 38536
rect 23164 38496 23170 38508
rect 24210 38496 24216 38508
rect 24268 38496 24274 38548
rect 24486 38496 24492 38548
rect 24544 38536 24550 38548
rect 24544 38508 24900 38536
rect 24544 38496 24550 38508
rect 23658 38468 23664 38480
rect 23032 38440 23664 38468
rect 23658 38428 23664 38440
rect 23716 38428 23722 38480
rect 23842 38428 23848 38480
rect 23900 38468 23906 38480
rect 23946 38471 24004 38477
rect 23946 38468 23958 38471
rect 23900 38440 23958 38468
rect 23900 38428 23906 38440
rect 23946 38437 23958 38440
rect 23992 38437 24004 38471
rect 24228 38468 24256 38496
rect 24228 38440 24696 38468
rect 23946 38431 24004 38437
rect 20070 38409 20076 38412
rect 20064 38363 20076 38409
rect 20128 38400 20134 38412
rect 20128 38372 20164 38400
rect 20070 38360 20076 38363
rect 20128 38360 20134 38372
rect 22094 38360 22100 38412
rect 22152 38400 22158 38412
rect 24668 38409 24696 38440
rect 24872 38409 24900 38508
rect 27338 38496 27344 38548
rect 27396 38536 27402 38548
rect 30466 38536 30472 38548
rect 27396 38508 27752 38536
rect 27396 38496 27402 38508
rect 25314 38468 25320 38480
rect 24964 38440 25320 38468
rect 24964 38409 24992 38440
rect 25314 38428 25320 38440
rect 25372 38428 25378 38480
rect 26234 38468 26240 38480
rect 26195 38440 26240 38468
rect 26234 38428 26240 38440
rect 26292 38428 26298 38480
rect 27522 38468 27528 38480
rect 27483 38440 27528 38468
rect 27522 38428 27528 38440
rect 27580 38428 27586 38480
rect 27724 38477 27752 38508
rect 28368 38508 30472 38536
rect 27709 38471 27767 38477
rect 27709 38437 27721 38471
rect 27755 38437 27767 38471
rect 28258 38468 28264 38480
rect 27709 38431 27767 38437
rect 27816 38440 28264 38468
rect 24668 38403 24731 38409
rect 22152 38372 22197 38400
rect 24668 38374 24685 38403
rect 22152 38360 22158 38372
rect 24673 38369 24685 38374
rect 24719 38369 24731 38403
rect 24673 38363 24731 38369
rect 24857 38403 24915 38409
rect 24857 38369 24869 38403
rect 24903 38369 24915 38403
rect 24857 38363 24915 38369
rect 24949 38403 25007 38409
rect 24949 38369 24961 38403
rect 24995 38369 25007 38403
rect 25222 38400 25228 38412
rect 25183 38372 25228 38400
rect 24949 38363 25007 38369
rect 25222 38360 25228 38372
rect 25280 38360 25286 38412
rect 26421 38403 26479 38409
rect 26421 38369 26433 38403
rect 26467 38400 26479 38403
rect 26602 38400 26608 38412
rect 26467 38372 26608 38400
rect 26467 38369 26479 38372
rect 26421 38363 26479 38369
rect 26602 38360 26608 38372
rect 26660 38400 26666 38412
rect 27341 38403 27399 38409
rect 27341 38400 27353 38403
rect 26660 38372 27353 38400
rect 26660 38360 26666 38372
rect 27341 38369 27353 38372
rect 27387 38369 27399 38403
rect 27341 38363 27399 38369
rect 19610 38292 19616 38344
rect 19668 38332 19674 38344
rect 19797 38335 19855 38341
rect 19797 38332 19809 38335
rect 19668 38304 19809 38332
rect 19668 38292 19674 38304
rect 19797 38301 19809 38304
rect 19843 38301 19855 38335
rect 19797 38295 19855 38301
rect 24213 38335 24271 38341
rect 24213 38301 24225 38335
rect 24259 38332 24271 38335
rect 25041 38335 25099 38341
rect 24259 38304 24900 38332
rect 24259 38301 24271 38304
rect 24213 38295 24271 38301
rect 24872 38276 24900 38304
rect 25041 38301 25053 38335
rect 25087 38301 25099 38335
rect 25041 38295 25099 38301
rect 24854 38224 24860 38276
rect 24912 38224 24918 38276
rect 21174 38196 21180 38208
rect 17000 38168 19334 38196
rect 21135 38168 21180 38196
rect 17000 38156 17006 38168
rect 21174 38156 21180 38168
rect 21232 38156 21238 38208
rect 22094 38156 22100 38208
rect 22152 38196 22158 38208
rect 22189 38199 22247 38205
rect 22189 38196 22201 38199
rect 22152 38168 22201 38196
rect 22152 38156 22158 38168
rect 22189 38165 22201 38168
rect 22235 38165 22247 38199
rect 22189 38159 22247 38165
rect 22833 38199 22891 38205
rect 22833 38165 22845 38199
rect 22879 38196 22891 38199
rect 23566 38196 23572 38208
rect 22879 38168 23572 38196
rect 22879 38165 22891 38168
rect 22833 38159 22891 38165
rect 23566 38156 23572 38168
rect 23624 38156 23630 38208
rect 23842 38156 23848 38208
rect 23900 38196 23906 38208
rect 24394 38196 24400 38208
rect 23900 38168 24400 38196
rect 23900 38156 23906 38168
rect 24394 38156 24400 38168
rect 24452 38156 24458 38208
rect 24762 38156 24768 38208
rect 24820 38196 24826 38208
rect 25056 38196 25084 38295
rect 27706 38292 27712 38344
rect 27764 38332 27770 38344
rect 27816 38332 27844 38440
rect 28258 38428 28264 38440
rect 28316 38428 28322 38480
rect 28166 38400 28172 38412
rect 28127 38372 28172 38400
rect 28166 38360 28172 38372
rect 28224 38360 28230 38412
rect 28368 38409 28396 38508
rect 30466 38496 30472 38508
rect 30524 38496 30530 38548
rect 31110 38496 31116 38548
rect 31168 38536 31174 38548
rect 31205 38539 31263 38545
rect 31205 38536 31217 38539
rect 31168 38508 31217 38536
rect 31168 38496 31174 38508
rect 31205 38505 31217 38508
rect 31251 38505 31263 38539
rect 31205 38499 31263 38505
rect 28534 38468 28540 38480
rect 28460 38440 28540 38468
rect 28460 38409 28488 38440
rect 28534 38428 28540 38440
rect 28592 38428 28598 38480
rect 28905 38471 28963 38477
rect 28905 38437 28917 38471
rect 28951 38468 28963 38471
rect 29610 38471 29668 38477
rect 29610 38468 29622 38471
rect 28951 38440 29622 38468
rect 28951 38437 28963 38440
rect 28905 38431 28963 38437
rect 29610 38437 29622 38440
rect 29656 38437 29668 38471
rect 29610 38431 29668 38437
rect 28353 38403 28411 38409
rect 28353 38369 28365 38403
rect 28399 38369 28411 38403
rect 28353 38363 28411 38369
rect 28445 38403 28503 38409
rect 28445 38369 28457 38403
rect 28491 38369 28503 38403
rect 28445 38363 28503 38369
rect 27764 38304 27844 38332
rect 27764 38292 27770 38304
rect 27890 38292 27896 38344
rect 27948 38332 27954 38344
rect 28460 38332 28488 38363
rect 28718 38360 28724 38412
rect 28776 38400 28782 38412
rect 28776 38372 30788 38400
rect 28776 38360 28782 38372
rect 27948 38304 28488 38332
rect 28537 38335 28595 38341
rect 27948 38292 27954 38304
rect 28537 38301 28549 38335
rect 28583 38332 28595 38335
rect 28626 38332 28632 38344
rect 28583 38304 28632 38332
rect 28583 38301 28595 38304
rect 28537 38295 28595 38301
rect 28626 38292 28632 38304
rect 28684 38292 28690 38344
rect 29362 38332 29368 38344
rect 28966 38304 29368 38332
rect 25130 38224 25136 38276
rect 25188 38264 25194 38276
rect 25314 38264 25320 38276
rect 25188 38236 25320 38264
rect 25188 38224 25194 38236
rect 25314 38224 25320 38236
rect 25372 38224 25378 38276
rect 26234 38224 26240 38276
rect 26292 38264 26298 38276
rect 28966 38264 28994 38304
rect 29362 38292 29368 38304
rect 29420 38292 29426 38344
rect 26292 38236 28994 38264
rect 26292 38224 26298 38236
rect 30760 38208 30788 38372
rect 25406 38196 25412 38208
rect 24820 38168 25084 38196
rect 25367 38168 25412 38196
rect 24820 38156 24826 38168
rect 25406 38156 25412 38168
rect 25464 38156 25470 38208
rect 26053 38199 26111 38205
rect 26053 38165 26065 38199
rect 26099 38196 26111 38199
rect 27798 38196 27804 38208
rect 26099 38168 27804 38196
rect 26099 38165 26111 38168
rect 26053 38159 26111 38165
rect 27798 38156 27804 38168
rect 27856 38156 27862 38208
rect 28074 38156 28080 38208
rect 28132 38196 28138 38208
rect 28902 38196 28908 38208
rect 28132 38168 28908 38196
rect 28132 38156 28138 38168
rect 28902 38156 28908 38168
rect 28960 38156 28966 38208
rect 30742 38196 30748 38208
rect 30703 38168 30748 38196
rect 30742 38156 30748 38168
rect 30800 38156 30806 38208
rect 1104 38106 32016 38128
rect 1104 38054 6102 38106
rect 6154 38054 6166 38106
rect 6218 38054 6230 38106
rect 6282 38054 6294 38106
rect 6346 38054 6358 38106
rect 6410 38054 16405 38106
rect 16457 38054 16469 38106
rect 16521 38054 16533 38106
rect 16585 38054 16597 38106
rect 16649 38054 16661 38106
rect 16713 38054 26709 38106
rect 26761 38054 26773 38106
rect 26825 38054 26837 38106
rect 26889 38054 26901 38106
rect 26953 38054 26965 38106
rect 27017 38054 32016 38106
rect 1104 38032 32016 38054
rect 5350 37952 5356 38004
rect 5408 37992 5414 38004
rect 5537 37995 5595 38001
rect 5537 37992 5549 37995
rect 5408 37964 5549 37992
rect 5408 37952 5414 37964
rect 5537 37961 5549 37964
rect 5583 37961 5595 37995
rect 5537 37955 5595 37961
rect 7009 37995 7067 38001
rect 7009 37961 7021 37995
rect 7055 37992 7067 37995
rect 7466 37992 7472 38004
rect 7055 37964 7472 37992
rect 7055 37961 7067 37964
rect 7009 37955 7067 37961
rect 7466 37952 7472 37964
rect 7524 37952 7530 38004
rect 9033 37995 9091 38001
rect 9033 37961 9045 37995
rect 9079 37992 9091 37995
rect 9398 37992 9404 38004
rect 9079 37964 9404 37992
rect 9079 37961 9091 37964
rect 9033 37955 9091 37961
rect 9398 37952 9404 37964
rect 9456 37952 9462 38004
rect 9490 37952 9496 38004
rect 9548 37992 9554 38004
rect 9677 37995 9735 38001
rect 9677 37992 9689 37995
rect 9548 37964 9689 37992
rect 9548 37952 9554 37964
rect 9677 37961 9689 37964
rect 9723 37961 9735 37995
rect 15286 37992 15292 38004
rect 9677 37955 9735 37961
rect 10980 37964 11928 37992
rect 15247 37964 15292 37992
rect 3878 37884 3884 37936
rect 3936 37924 3942 37936
rect 10980 37924 11008 37964
rect 11900 37936 11928 37964
rect 15286 37952 15292 37964
rect 15344 37952 15350 38004
rect 18690 37992 18696 38004
rect 16776 37964 18696 37992
rect 3936 37896 4476 37924
rect 3936 37884 3942 37896
rect 4246 37856 4252 37868
rect 4207 37828 4252 37856
rect 4246 37816 4252 37828
rect 4304 37816 4310 37868
rect 0 37788 800 37802
rect 4448 37800 4476 37896
rect 10888 37896 11008 37924
rect 5902 37816 5908 37868
rect 5960 37856 5966 37868
rect 10888 37865 10916 37896
rect 11146 37884 11152 37936
rect 11204 37924 11210 37936
rect 11790 37924 11796 37936
rect 11204 37896 11796 37924
rect 11204 37884 11210 37896
rect 11790 37884 11796 37896
rect 11848 37884 11854 37936
rect 11882 37884 11888 37936
rect 11940 37924 11946 37936
rect 12066 37924 12072 37936
rect 11940 37896 12072 37924
rect 11940 37884 11946 37896
rect 12066 37884 12072 37896
rect 12124 37924 12130 37936
rect 12802 37924 12808 37936
rect 12124 37896 12808 37924
rect 12124 37884 12130 37896
rect 12802 37884 12808 37896
rect 12860 37924 12866 37936
rect 13170 37924 13176 37936
rect 12860 37896 13176 37924
rect 12860 37884 12866 37896
rect 13170 37884 13176 37896
rect 13228 37884 13234 37936
rect 14737 37927 14795 37933
rect 14737 37893 14749 37927
rect 14783 37924 14795 37927
rect 15470 37924 15476 37936
rect 14783 37896 15476 37924
rect 14783 37893 14795 37896
rect 14737 37887 14795 37893
rect 15470 37884 15476 37896
rect 15528 37884 15534 37936
rect 7101 37859 7159 37865
rect 7101 37856 7113 37859
rect 5960 37828 7113 37856
rect 5960 37816 5966 37828
rect 7101 37825 7113 37828
rect 7147 37825 7159 37859
rect 7101 37819 7159 37825
rect 10873 37859 10931 37865
rect 10873 37825 10885 37859
rect 10919 37825 10931 37859
rect 10873 37819 10931 37825
rect 10965 37859 11023 37865
rect 10965 37825 10977 37859
rect 11011 37856 11023 37859
rect 11977 37859 12035 37865
rect 11977 37856 11989 37859
rect 11011 37828 11989 37856
rect 11011 37825 11023 37828
rect 10965 37819 11023 37825
rect 11977 37825 11989 37828
rect 12023 37856 12035 37859
rect 12434 37856 12440 37868
rect 12023 37828 12440 37856
rect 12023 37825 12035 37828
rect 11977 37819 12035 37825
rect 12434 37816 12440 37828
rect 12492 37856 12498 37868
rect 12710 37856 12716 37868
rect 12492 37828 12716 37856
rect 12492 37816 12498 37828
rect 12710 37816 12716 37828
rect 12768 37816 12774 37868
rect 15746 37856 15752 37868
rect 15707 37828 15752 37856
rect 15746 37816 15752 37828
rect 15804 37816 15810 37868
rect 1857 37791 1915 37797
rect 1857 37788 1869 37791
rect 0 37760 1869 37788
rect 0 37746 800 37760
rect 1857 37757 1869 37760
rect 1903 37788 1915 37791
rect 2038 37788 2044 37800
rect 1903 37760 2044 37788
rect 1903 37757 1915 37760
rect 1857 37751 1915 37757
rect 2038 37748 2044 37760
rect 2096 37748 2102 37800
rect 3142 37748 3148 37800
rect 3200 37788 3206 37800
rect 3973 37791 4031 37797
rect 3973 37788 3985 37791
rect 3200 37760 3985 37788
rect 3200 37748 3206 37760
rect 3973 37757 3985 37760
rect 4019 37757 4031 37791
rect 4154 37788 4160 37800
rect 4115 37760 4160 37788
rect 3973 37751 4031 37757
rect 4154 37748 4160 37760
rect 4212 37748 4218 37800
rect 4338 37788 4344 37800
rect 4299 37760 4344 37788
rect 4338 37748 4344 37760
rect 4396 37748 4402 37800
rect 4430 37748 4436 37800
rect 4488 37788 4494 37800
rect 4525 37791 4583 37797
rect 4525 37788 4537 37791
rect 4488 37760 4537 37788
rect 4488 37748 4494 37760
rect 4525 37757 4537 37760
rect 4571 37757 4583 37791
rect 6822 37788 6828 37800
rect 6783 37760 6828 37788
rect 4525 37751 4583 37757
rect 6822 37748 6828 37760
rect 6880 37748 6886 37800
rect 6917 37791 6975 37797
rect 6917 37757 6929 37791
rect 6963 37788 6975 37791
rect 7282 37788 7288 37800
rect 6963 37760 7288 37788
rect 6963 37757 6975 37760
rect 6917 37751 6975 37757
rect 7282 37748 7288 37760
rect 7340 37788 7346 37800
rect 7558 37788 7564 37800
rect 7340 37760 7564 37788
rect 7340 37748 7346 37760
rect 7558 37748 7564 37760
rect 7616 37748 7622 37800
rect 8938 37788 8944 37800
rect 8899 37760 8944 37788
rect 8938 37748 8944 37760
rect 8996 37748 9002 37800
rect 9861 37791 9919 37797
rect 9861 37757 9873 37791
rect 9907 37788 9919 37791
rect 10410 37788 10416 37800
rect 9907 37760 10416 37788
rect 9907 37757 9919 37760
rect 9861 37751 9919 37757
rect 10410 37748 10416 37760
rect 10468 37748 10474 37800
rect 10689 37791 10747 37797
rect 10689 37757 10701 37791
rect 10735 37757 10747 37791
rect 10689 37751 10747 37757
rect 11057 37791 11115 37797
rect 11057 37757 11069 37791
rect 11103 37788 11115 37791
rect 11146 37788 11152 37800
rect 11103 37760 11152 37788
rect 11103 37757 11115 37760
rect 11057 37751 11115 37757
rect 2225 37723 2283 37729
rect 2225 37689 2237 37723
rect 2271 37720 2283 37723
rect 7374 37720 7380 37732
rect 2271 37692 3188 37720
rect 2271 37689 2283 37692
rect 2225 37683 2283 37689
rect 2590 37612 2596 37664
rect 2648 37652 2654 37664
rect 2685 37655 2743 37661
rect 2685 37652 2697 37655
rect 2648 37624 2697 37652
rect 2648 37612 2654 37624
rect 2685 37621 2697 37624
rect 2731 37621 2743 37655
rect 3160 37652 3188 37692
rect 6840 37692 7380 37720
rect 6840 37664 6868 37692
rect 7374 37680 7380 37692
rect 7432 37680 7438 37732
rect 10042 37720 10048 37732
rect 10003 37692 10048 37720
rect 10042 37680 10048 37692
rect 10100 37680 10106 37732
rect 10704 37720 10732 37751
rect 11146 37748 11152 37760
rect 11204 37748 11210 37800
rect 11241 37791 11299 37797
rect 11241 37757 11253 37791
rect 11287 37788 11299 37791
rect 11698 37788 11704 37800
rect 11287 37760 11704 37788
rect 11287 37757 11299 37760
rect 11241 37751 11299 37757
rect 11698 37748 11704 37760
rect 11756 37748 11762 37800
rect 11882 37788 11888 37800
rect 11795 37760 11888 37788
rect 11808 37720 11836 37760
rect 11882 37748 11888 37760
rect 11940 37748 11946 37800
rect 12066 37788 12072 37800
rect 12027 37760 12072 37788
rect 12066 37748 12072 37760
rect 12124 37748 12130 37800
rect 12253 37791 12311 37797
rect 12253 37757 12265 37791
rect 12299 37788 12311 37791
rect 12618 37788 12624 37800
rect 12299 37760 12624 37788
rect 12299 37757 12311 37760
rect 12253 37751 12311 37757
rect 12618 37748 12624 37760
rect 12676 37748 12682 37800
rect 12986 37788 12992 37800
rect 12899 37760 12992 37788
rect 12986 37748 12992 37760
rect 13044 37788 13050 37800
rect 13170 37788 13176 37800
rect 13044 37760 13176 37788
rect 13044 37748 13050 37760
rect 13170 37748 13176 37760
rect 13228 37748 13234 37800
rect 14550 37748 14556 37800
rect 14608 37788 14614 37800
rect 14645 37791 14703 37797
rect 14645 37788 14657 37791
rect 14608 37760 14657 37788
rect 14608 37748 14614 37760
rect 14645 37757 14657 37760
rect 14691 37788 14703 37791
rect 15102 37788 15108 37800
rect 14691 37760 15108 37788
rect 14691 37757 14703 37760
rect 14645 37751 14703 37757
rect 15102 37748 15108 37760
rect 15160 37788 15166 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 15160 37760 15485 37788
rect 15160 37748 15166 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 15473 37751 15531 37757
rect 15565 37791 15623 37797
rect 15565 37757 15577 37791
rect 15611 37757 15623 37791
rect 15565 37751 15623 37757
rect 15657 37791 15715 37797
rect 15657 37757 15669 37791
rect 15703 37788 15715 37791
rect 15838 37788 15844 37800
rect 15703 37760 15844 37788
rect 15703 37757 15715 37760
rect 15657 37751 15715 37757
rect 10704 37692 11836 37720
rect 15378 37680 15384 37732
rect 15436 37720 15442 37732
rect 15580 37720 15608 37751
rect 15838 37748 15844 37760
rect 15896 37748 15902 37800
rect 15930 37748 15936 37800
rect 15988 37788 15994 37800
rect 16776 37788 16804 37964
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 20070 37992 20076 38004
rect 20031 37964 20076 37992
rect 20070 37952 20076 37964
rect 20128 37952 20134 38004
rect 20530 37952 20536 38004
rect 20588 37992 20594 38004
rect 20625 37995 20683 38001
rect 20625 37992 20637 37995
rect 20588 37964 20637 37992
rect 20588 37952 20594 37964
rect 20625 37961 20637 37964
rect 20671 37992 20683 37995
rect 22462 37992 22468 38004
rect 20671 37964 22324 37992
rect 22423 37964 22468 37992
rect 20671 37961 20683 37964
rect 20625 37955 20683 37961
rect 17402 37924 17408 37936
rect 17328 37896 17408 37924
rect 17328 37865 17356 37896
rect 17402 37884 17408 37896
rect 17460 37884 17466 37936
rect 17494 37884 17500 37936
rect 17552 37924 17558 37936
rect 18601 37927 18659 37933
rect 17552 37896 17908 37924
rect 17552 37884 17558 37896
rect 17313 37859 17371 37865
rect 17313 37825 17325 37859
rect 17359 37825 17371 37859
rect 17770 37856 17776 37868
rect 17313 37819 17371 37825
rect 17420 37828 17776 37856
rect 15988 37760 16804 37788
rect 15988 37748 15994 37760
rect 16942 37748 16948 37800
rect 17000 37748 17006 37800
rect 17420 37797 17448 37828
rect 17770 37816 17776 37828
rect 17828 37816 17834 37868
rect 17129 37791 17187 37797
rect 17129 37757 17141 37791
rect 17175 37757 17187 37791
rect 17129 37751 17187 37757
rect 17405 37791 17463 37797
rect 17405 37757 17417 37791
rect 17451 37757 17463 37791
rect 17405 37751 17463 37757
rect 17497 37791 17555 37797
rect 17497 37757 17509 37791
rect 17543 37757 17555 37791
rect 17497 37751 17555 37757
rect 17681 37791 17739 37797
rect 17681 37757 17693 37791
rect 17727 37788 17739 37791
rect 17880 37788 17908 37896
rect 18601 37893 18613 37927
rect 18647 37924 18659 37927
rect 20714 37924 20720 37936
rect 18647 37896 20720 37924
rect 18647 37893 18659 37896
rect 18601 37887 18659 37893
rect 20714 37884 20720 37896
rect 20772 37884 20778 37936
rect 21269 37927 21327 37933
rect 21269 37893 21281 37927
rect 21315 37924 21327 37927
rect 22296 37924 22324 37964
rect 22462 37952 22468 37964
rect 22520 37952 22526 38004
rect 23014 37952 23020 38004
rect 23072 37992 23078 38004
rect 24765 37995 24823 38001
rect 24765 37992 24777 37995
rect 23072 37964 24777 37992
rect 23072 37952 23078 37964
rect 24765 37961 24777 37964
rect 24811 37992 24823 37995
rect 25222 37992 25228 38004
rect 24811 37964 25228 37992
rect 24811 37961 24823 37964
rect 24765 37955 24823 37961
rect 25222 37952 25228 37964
rect 25280 37952 25286 38004
rect 26602 37952 26608 38004
rect 26660 37992 26666 38004
rect 26697 37995 26755 38001
rect 26697 37992 26709 37995
rect 26660 37964 26709 37992
rect 26660 37952 26666 37964
rect 26697 37961 26709 37964
rect 26743 37961 26755 37995
rect 27338 37992 27344 38004
rect 27299 37964 27344 37992
rect 26697 37955 26755 37961
rect 27338 37952 27344 37964
rect 27396 37952 27402 38004
rect 27522 37952 27528 38004
rect 27580 37992 27586 38004
rect 31110 37992 31116 38004
rect 27580 37964 31116 37992
rect 27580 37952 27586 37964
rect 31110 37952 31116 37964
rect 31168 37952 31174 38004
rect 25130 37924 25136 37936
rect 21315 37896 21864 37924
rect 22296 37896 25136 37924
rect 21315 37893 21327 37896
rect 21269 37887 21327 37893
rect 19613 37859 19671 37865
rect 19613 37825 19625 37859
rect 19659 37856 19671 37859
rect 19794 37856 19800 37868
rect 19659 37828 19800 37856
rect 19659 37825 19671 37828
rect 19613 37819 19671 37825
rect 19794 37816 19800 37828
rect 19852 37816 19858 37868
rect 21174 37856 21180 37868
rect 19904 37828 21180 37856
rect 18506 37788 18512 37800
rect 17727 37760 17908 37788
rect 18467 37760 18512 37788
rect 17727 37757 17739 37760
rect 17681 37751 17739 37757
rect 16485 37723 16543 37729
rect 15436 37692 15884 37720
rect 15436 37680 15442 37692
rect 15856 37664 15884 37692
rect 16485 37689 16497 37723
rect 16531 37720 16543 37723
rect 16960 37720 16988 37748
rect 16531 37692 16988 37720
rect 16531 37689 16543 37692
rect 16485 37683 16543 37689
rect 3510 37652 3516 37664
rect 3160 37624 3516 37652
rect 2685 37615 2743 37621
rect 3510 37612 3516 37624
rect 3568 37612 3574 37664
rect 3786 37652 3792 37664
rect 3747 37624 3792 37652
rect 3786 37612 3792 37624
rect 3844 37612 3850 37664
rect 4982 37612 4988 37664
rect 5040 37652 5046 37664
rect 5077 37655 5135 37661
rect 5077 37652 5089 37655
rect 5040 37624 5089 37652
rect 5040 37612 5046 37624
rect 5077 37621 5089 37624
rect 5123 37652 5135 37655
rect 5810 37652 5816 37664
rect 5123 37624 5816 37652
rect 5123 37621 5135 37624
rect 5077 37615 5135 37621
rect 5810 37612 5816 37624
rect 5868 37612 5874 37664
rect 6365 37655 6423 37661
rect 6365 37621 6377 37655
rect 6411 37652 6423 37655
rect 6822 37652 6828 37664
rect 6411 37624 6828 37652
rect 6411 37621 6423 37624
rect 6365 37615 6423 37621
rect 6822 37612 6828 37624
rect 6880 37612 6886 37664
rect 7190 37612 7196 37664
rect 7248 37652 7254 37664
rect 8113 37655 8171 37661
rect 8113 37652 8125 37655
rect 7248 37624 8125 37652
rect 7248 37612 7254 37624
rect 8113 37621 8125 37624
rect 8159 37621 8171 37655
rect 8113 37615 8171 37621
rect 10505 37655 10563 37661
rect 10505 37621 10517 37655
rect 10551 37652 10563 37655
rect 10778 37652 10784 37664
rect 10551 37624 10784 37652
rect 10551 37621 10563 37624
rect 10505 37615 10563 37621
rect 10778 37612 10784 37624
rect 10836 37612 10842 37664
rect 10962 37612 10968 37664
rect 11020 37652 11026 37664
rect 11698 37652 11704 37664
rect 11020 37624 11704 37652
rect 11020 37612 11026 37624
rect 11698 37612 11704 37624
rect 11756 37612 11762 37664
rect 12342 37612 12348 37664
rect 12400 37652 12406 37664
rect 12437 37655 12495 37661
rect 12437 37652 12449 37655
rect 12400 37624 12449 37652
rect 12400 37612 12406 37624
rect 12437 37621 12449 37624
rect 12483 37621 12495 37655
rect 12437 37615 12495 37621
rect 12986 37612 12992 37664
rect 13044 37652 13050 37664
rect 13449 37655 13507 37661
rect 13449 37652 13461 37655
rect 13044 37624 13461 37652
rect 13044 37612 13050 37624
rect 13449 37621 13461 37624
rect 13495 37621 13507 37655
rect 13449 37615 13507 37621
rect 13998 37612 14004 37664
rect 14056 37652 14062 37664
rect 14093 37655 14151 37661
rect 14093 37652 14105 37655
rect 14056 37624 14105 37652
rect 14056 37612 14062 37624
rect 14093 37621 14105 37624
rect 14139 37621 14151 37655
rect 14093 37615 14151 37621
rect 15838 37612 15844 37664
rect 15896 37612 15902 37664
rect 16942 37652 16948 37664
rect 16903 37624 16948 37652
rect 16942 37612 16948 37624
rect 17000 37612 17006 37664
rect 17144 37652 17172 37751
rect 17512 37720 17540 37751
rect 18506 37748 18512 37760
rect 18564 37748 18570 37800
rect 19337 37791 19395 37797
rect 19337 37757 19349 37791
rect 19383 37788 19395 37791
rect 19426 37788 19432 37800
rect 19383 37760 19432 37788
rect 19383 37757 19395 37760
rect 19337 37751 19395 37757
rect 19426 37748 19432 37760
rect 19484 37748 19490 37800
rect 19521 37791 19579 37797
rect 19521 37757 19533 37791
rect 19567 37757 19579 37791
rect 19702 37788 19708 37800
rect 19663 37760 19708 37788
rect 19521 37751 19579 37757
rect 17954 37720 17960 37732
rect 17512 37692 17960 37720
rect 17954 37680 17960 37692
rect 18012 37720 18018 37732
rect 19058 37720 19064 37732
rect 18012 37692 19064 37720
rect 18012 37680 18018 37692
rect 19058 37680 19064 37692
rect 19116 37680 19122 37732
rect 19536 37720 19564 37751
rect 19702 37748 19708 37760
rect 19760 37748 19766 37800
rect 19904 37797 19932 37828
rect 21174 37816 21180 37828
rect 21232 37816 21238 37868
rect 21836 37865 21864 37896
rect 25130 37884 25136 37896
rect 25188 37884 25194 37936
rect 27246 37884 27252 37936
rect 27304 37884 27310 37936
rect 28994 37924 29000 37936
rect 28690 37896 29000 37924
rect 21821 37859 21879 37865
rect 21821 37825 21833 37859
rect 21867 37825 21879 37859
rect 21821 37819 21879 37825
rect 21910 37816 21916 37868
rect 21968 37856 21974 37868
rect 22186 37856 22192 37868
rect 21968 37828 22192 37856
rect 21968 37816 21974 37828
rect 22186 37816 22192 37828
rect 22244 37816 22250 37868
rect 23198 37816 23204 37868
rect 23256 37856 23262 37868
rect 23394 37859 23452 37865
rect 23394 37856 23406 37859
rect 23256 37828 23406 37856
rect 23256 37816 23262 37828
rect 23394 37825 23406 37828
rect 23440 37825 23452 37859
rect 23394 37819 23452 37825
rect 23845 37859 23903 37865
rect 23845 37825 23857 37859
rect 23891 37856 23903 37859
rect 24394 37856 24400 37868
rect 23891 37828 24400 37856
rect 23891 37825 23903 37828
rect 23845 37819 23903 37825
rect 24394 37816 24400 37828
rect 24452 37816 24458 37868
rect 27264 37856 27292 37884
rect 27264 37828 27568 37856
rect 19889 37791 19947 37797
rect 19889 37757 19901 37791
rect 19935 37757 19947 37791
rect 21082 37788 21088 37800
rect 21043 37760 21088 37788
rect 19889 37751 19947 37757
rect 21082 37748 21088 37760
rect 21140 37748 21146 37800
rect 22094 37748 22100 37800
rect 22152 37788 22158 37800
rect 23106 37788 23112 37800
rect 22152 37760 22197 37788
rect 23067 37760 23112 37788
rect 22152 37748 22158 37760
rect 23106 37748 23112 37760
rect 23164 37748 23170 37800
rect 23293 37791 23351 37797
rect 23293 37757 23305 37791
rect 23339 37757 23351 37791
rect 23474 37788 23480 37800
rect 23435 37760 23480 37788
rect 23293 37751 23351 37757
rect 19794 37720 19800 37732
rect 19536 37692 19800 37720
rect 19794 37680 19800 37692
rect 19852 37720 19858 37732
rect 19852 37692 21036 37720
rect 19852 37680 19858 37692
rect 21008 37664 21036 37692
rect 21358 37680 21364 37732
rect 21416 37720 21422 37732
rect 23308 37720 23336 37751
rect 23474 37748 23480 37760
rect 23532 37748 23538 37800
rect 23658 37788 23664 37800
rect 23619 37760 23664 37788
rect 23658 37748 23664 37760
rect 23716 37788 23722 37800
rect 24486 37788 24492 37800
rect 23716 37760 24492 37788
rect 23716 37748 23722 37760
rect 24486 37748 24492 37760
rect 24544 37748 24550 37800
rect 25406 37748 25412 37800
rect 25464 37788 25470 37800
rect 25878 37791 25936 37797
rect 25878 37788 25890 37791
rect 25464 37760 25890 37788
rect 25464 37748 25470 37760
rect 25878 37757 25890 37760
rect 25924 37757 25936 37791
rect 25878 37751 25936 37757
rect 26145 37791 26203 37797
rect 26145 37757 26157 37791
rect 26191 37788 26203 37791
rect 26234 37788 26240 37800
rect 26191 37760 26240 37788
rect 26191 37757 26203 37760
rect 26145 37751 26203 37757
rect 26234 37748 26240 37760
rect 26292 37748 26298 37800
rect 27540 37797 27568 37828
rect 27890 37816 27896 37868
rect 27948 37856 27954 37868
rect 27948 37828 28589 37856
rect 27948 37816 27954 37828
rect 26789 37791 26847 37797
rect 26789 37757 26801 37791
rect 26835 37757 26847 37791
rect 26789 37751 26847 37757
rect 27249 37791 27307 37797
rect 27249 37757 27261 37791
rect 27295 37757 27307 37791
rect 27249 37751 27307 37757
rect 27525 37791 27583 37797
rect 27525 37757 27537 37791
rect 27571 37757 27583 37791
rect 27525 37751 27583 37757
rect 23566 37720 23572 37732
rect 21416 37692 23244 37720
rect 23308 37692 23572 37720
rect 21416 37680 21422 37692
rect 17862 37652 17868 37664
rect 17144 37624 17868 37652
rect 17862 37612 17868 37624
rect 17920 37612 17926 37664
rect 20990 37612 20996 37664
rect 21048 37652 21054 37664
rect 22005 37655 22063 37661
rect 22005 37652 22017 37655
rect 21048 37624 22017 37652
rect 21048 37612 21054 37624
rect 22005 37621 22017 37624
rect 22051 37621 22063 37655
rect 23216 37652 23244 37692
rect 23566 37680 23572 37692
rect 23624 37720 23630 37732
rect 23750 37720 23756 37732
rect 23624 37692 23756 37720
rect 23624 37680 23630 37692
rect 23750 37680 23756 37692
rect 23808 37680 23814 37732
rect 25774 37720 25780 37732
rect 24688 37692 25780 37720
rect 24688 37652 24716 37692
rect 25774 37680 25780 37692
rect 25832 37720 25838 37732
rect 26418 37720 26424 37732
rect 25832 37692 26424 37720
rect 25832 37680 25838 37692
rect 26418 37680 26424 37692
rect 26476 37720 26482 37732
rect 26804 37720 26832 37751
rect 26476 37692 26832 37720
rect 27264 37720 27292 37751
rect 27614 37748 27620 37800
rect 27672 37788 27678 37800
rect 27672 37760 27717 37788
rect 27672 37748 27678 37760
rect 28166 37748 28172 37800
rect 28224 37788 28230 37800
rect 28561 37797 28589 37828
rect 28690 37797 28718 37896
rect 28994 37884 29000 37896
rect 29052 37884 29058 37936
rect 29178 37856 29184 37868
rect 28828 37828 29184 37856
rect 28828 37797 28856 37828
rect 29178 37816 29184 37828
rect 29236 37816 29242 37868
rect 29362 37816 29368 37868
rect 29420 37856 29426 37868
rect 29549 37859 29607 37865
rect 29549 37856 29561 37859
rect 29420 37828 29561 37856
rect 29420 37816 29426 37828
rect 29549 37825 29561 37828
rect 29595 37825 29607 37859
rect 29549 37819 29607 37825
rect 28261 37791 28319 37797
rect 28261 37788 28273 37791
rect 28224 37760 28273 37788
rect 28224 37748 28230 37760
rect 28261 37757 28273 37760
rect 28307 37757 28319 37791
rect 28261 37751 28319 37757
rect 28445 37791 28503 37797
rect 28445 37757 28457 37791
rect 28491 37757 28503 37791
rect 28445 37751 28503 37757
rect 28531 37791 28589 37797
rect 28531 37757 28543 37791
rect 28577 37757 28589 37791
rect 28531 37751 28589 37757
rect 28675 37791 28733 37797
rect 28675 37757 28687 37791
rect 28721 37757 28733 37791
rect 28675 37751 28733 37757
rect 28813 37791 28871 37797
rect 28813 37757 28825 37791
rect 28859 37757 28871 37791
rect 28813 37751 28871 37757
rect 28074 37720 28080 37732
rect 27264 37692 28080 37720
rect 26476 37680 26482 37692
rect 28074 37680 28080 37692
rect 28132 37680 28138 37732
rect 28460 37720 28488 37751
rect 28902 37748 28908 37800
rect 28960 37788 28966 37800
rect 30374 37788 30380 37800
rect 28960 37760 30380 37788
rect 28960 37748 28966 37760
rect 30374 37748 30380 37760
rect 30432 37748 30438 37800
rect 32320 37788 33120 37802
rect 32048 37760 33120 37788
rect 28997 37723 29055 37729
rect 28460 37692 28764 37720
rect 28736 37664 28764 37692
rect 28997 37689 29009 37723
rect 29043 37720 29055 37723
rect 29794 37723 29852 37729
rect 29794 37720 29806 37723
rect 29043 37692 29806 37720
rect 29043 37689 29055 37692
rect 28997 37683 29055 37689
rect 29794 37689 29806 37692
rect 29840 37689 29852 37723
rect 29794 37683 29852 37689
rect 23216 37624 24716 37652
rect 27801 37655 27859 37661
rect 22005 37615 22063 37621
rect 27801 37621 27813 37655
rect 27847 37652 27859 37655
rect 27890 37652 27896 37664
rect 27847 37624 27896 37652
rect 27847 37621 27859 37624
rect 27801 37615 27859 37621
rect 27890 37612 27896 37624
rect 27948 37612 27954 37664
rect 28718 37612 28724 37664
rect 28776 37612 28782 37664
rect 29178 37612 29184 37664
rect 29236 37652 29242 37664
rect 30929 37655 30987 37661
rect 30929 37652 30941 37655
rect 29236 37624 30941 37652
rect 29236 37612 29242 37624
rect 30929 37621 30941 37624
rect 30975 37621 30987 37655
rect 30929 37615 30987 37621
rect 1104 37562 32016 37584
rect 1104 37510 11253 37562
rect 11305 37510 11317 37562
rect 11369 37510 11381 37562
rect 11433 37510 11445 37562
rect 11497 37510 11509 37562
rect 11561 37510 21557 37562
rect 21609 37510 21621 37562
rect 21673 37510 21685 37562
rect 21737 37510 21749 37562
rect 21801 37510 21813 37562
rect 21865 37510 32016 37562
rect 1104 37488 32016 37510
rect 2501 37451 2559 37457
rect 2501 37417 2513 37451
rect 2547 37448 2559 37451
rect 3142 37448 3148 37460
rect 2547 37420 3148 37448
rect 2547 37417 2559 37420
rect 2501 37411 2559 37417
rect 3142 37408 3148 37420
rect 3200 37408 3206 37460
rect 5718 37408 5724 37460
rect 5776 37448 5782 37460
rect 5813 37451 5871 37457
rect 5813 37448 5825 37451
rect 5776 37420 5825 37448
rect 5776 37408 5782 37420
rect 5813 37417 5825 37420
rect 5859 37417 5871 37451
rect 5813 37411 5871 37417
rect 7282 37408 7288 37460
rect 7340 37448 7346 37460
rect 8021 37451 8079 37457
rect 8021 37448 8033 37451
rect 7340 37420 8033 37448
rect 7340 37408 7346 37420
rect 8021 37417 8033 37420
rect 8067 37448 8079 37451
rect 8386 37448 8392 37460
rect 8067 37420 8392 37448
rect 8067 37417 8079 37420
rect 8021 37411 8079 37417
rect 8386 37408 8392 37420
rect 8444 37408 8450 37460
rect 8481 37451 8539 37457
rect 8481 37417 8493 37451
rect 8527 37448 8539 37451
rect 9122 37448 9128 37460
rect 8527 37420 9128 37448
rect 8527 37417 8539 37420
rect 8481 37411 8539 37417
rect 9122 37408 9128 37420
rect 9180 37448 9186 37460
rect 9398 37448 9404 37460
rect 9180 37420 9404 37448
rect 9180 37408 9186 37420
rect 9398 37408 9404 37420
rect 9456 37408 9462 37460
rect 9950 37448 9956 37460
rect 9646 37420 9956 37448
rect 3636 37383 3694 37389
rect 3636 37349 3648 37383
rect 3682 37380 3694 37383
rect 3786 37380 3792 37392
rect 3682 37352 3792 37380
rect 3682 37349 3694 37352
rect 3636 37343 3694 37349
rect 3786 37340 3792 37352
rect 3844 37340 3850 37392
rect 4448 37352 5304 37380
rect 2041 37315 2099 37321
rect 2041 37281 2053 37315
rect 2087 37312 2099 37315
rect 2130 37312 2136 37324
rect 2087 37284 2136 37312
rect 2087 37281 2099 37284
rect 2041 37275 2099 37281
rect 2130 37272 2136 37284
rect 2188 37312 2194 37324
rect 2498 37312 2504 37324
rect 2188 37284 2504 37312
rect 2188 37272 2194 37284
rect 2498 37272 2504 37284
rect 2556 37272 2562 37324
rect 3878 37312 3884 37324
rect 3791 37284 3884 37312
rect 3878 37272 3884 37284
rect 3936 37312 3942 37324
rect 4448 37321 4476 37352
rect 5276 37324 5304 37352
rect 6454 37340 6460 37392
rect 6512 37380 6518 37392
rect 9646 37380 9674 37420
rect 9950 37408 9956 37420
rect 10008 37408 10014 37460
rect 12618 37408 12624 37460
rect 12676 37448 12682 37460
rect 13449 37451 13507 37457
rect 13449 37448 13461 37451
rect 12676 37420 13461 37448
rect 12676 37408 12682 37420
rect 13449 37417 13461 37420
rect 13495 37417 13507 37451
rect 13449 37411 13507 37417
rect 14921 37451 14979 37457
rect 14921 37417 14933 37451
rect 14967 37448 14979 37451
rect 15749 37451 15807 37457
rect 14967 37420 15700 37448
rect 14967 37417 14979 37420
rect 14921 37411 14979 37417
rect 11054 37380 11060 37392
rect 6512 37352 9674 37380
rect 9876 37352 11060 37380
rect 6512 37340 6518 37352
rect 4706 37321 4712 37324
rect 4433 37315 4491 37321
rect 4433 37312 4445 37315
rect 3936 37284 4445 37312
rect 3936 37272 3942 37284
rect 4433 37281 4445 37284
rect 4479 37281 4491 37315
rect 4700 37312 4712 37321
rect 4667 37284 4712 37312
rect 4433 37275 4491 37281
rect 4700 37275 4712 37284
rect 4706 37272 4712 37275
rect 4764 37272 4770 37324
rect 5258 37272 5264 37324
rect 5316 37312 5322 37324
rect 6638 37312 6644 37324
rect 5316 37284 6644 37312
rect 5316 37272 5322 37284
rect 6638 37272 6644 37284
rect 6696 37272 6702 37324
rect 6914 37321 6920 37324
rect 6908 37275 6920 37321
rect 6972 37312 6978 37324
rect 9605 37315 9663 37321
rect 6972 37284 7008 37312
rect 6914 37272 6920 37275
rect 6972 37272 6978 37284
rect 9605 37281 9617 37315
rect 9651 37312 9663 37315
rect 9766 37312 9772 37324
rect 9651 37284 9772 37312
rect 9651 37281 9663 37284
rect 9605 37275 9663 37281
rect 9766 37272 9772 37284
rect 9824 37272 9830 37324
rect 9876 37321 9904 37352
rect 11054 37340 11060 37352
rect 11112 37340 11118 37392
rect 13078 37380 13084 37392
rect 12084 37352 13084 37380
rect 9861 37315 9919 37321
rect 9861 37281 9873 37315
rect 9907 37281 9919 37315
rect 9861 37275 9919 37281
rect 10505 37315 10563 37321
rect 10505 37281 10517 37315
rect 10551 37312 10563 37315
rect 10870 37312 10876 37324
rect 10551 37284 10876 37312
rect 10551 37281 10563 37284
rect 10505 37275 10563 37281
rect 10870 37272 10876 37284
rect 10928 37272 10934 37324
rect 11146 37272 11152 37324
rect 11204 37312 11210 37324
rect 12084 37321 12112 37352
rect 13078 37340 13084 37352
rect 13136 37340 13142 37392
rect 15470 37340 15476 37392
rect 15528 37380 15534 37392
rect 15565 37383 15623 37389
rect 15565 37380 15577 37383
rect 15528 37352 15577 37380
rect 15528 37340 15534 37352
rect 15565 37349 15577 37352
rect 15611 37349 15623 37383
rect 15672 37380 15700 37420
rect 15749 37417 15761 37451
rect 15795 37448 15807 37451
rect 15930 37448 15936 37460
rect 15795 37420 15936 37448
rect 15795 37417 15807 37420
rect 15749 37411 15807 37417
rect 15930 37408 15936 37420
rect 15988 37408 15994 37460
rect 16298 37408 16304 37460
rect 16356 37448 16362 37460
rect 20990 37448 20996 37460
rect 16356 37420 20116 37448
rect 20951 37420 20996 37448
rect 16356 37408 16362 37420
rect 16945 37383 17003 37389
rect 15672 37352 16712 37380
rect 15565 37343 15623 37349
rect 12342 37321 12348 37324
rect 11517 37315 11575 37321
rect 11517 37312 11529 37315
rect 11204 37284 11529 37312
rect 11204 37272 11210 37284
rect 11517 37281 11529 37284
rect 11563 37281 11575 37315
rect 11517 37275 11575 37281
rect 12069 37315 12127 37321
rect 12069 37281 12081 37315
rect 12115 37281 12127 37315
rect 12336 37312 12348 37321
rect 12303 37284 12348 37312
rect 12069 37275 12127 37281
rect 12336 37275 12348 37284
rect 12342 37272 12348 37275
rect 12400 37272 12406 37324
rect 15381 37315 15439 37321
rect 15381 37281 15393 37315
rect 15427 37312 15439 37315
rect 15654 37312 15660 37324
rect 15427 37284 15660 37312
rect 15427 37281 15439 37284
rect 15381 37275 15439 37281
rect 15654 37272 15660 37284
rect 15712 37272 15718 37324
rect 16684 37244 16712 37352
rect 16945 37349 16957 37383
rect 16991 37380 17003 37383
rect 17034 37380 17040 37392
rect 16991 37352 17040 37380
rect 16991 37349 17003 37352
rect 16945 37343 17003 37349
rect 17034 37340 17040 37352
rect 17092 37340 17098 37392
rect 17696 37352 19656 37380
rect 16850 37312 16856 37324
rect 16811 37284 16856 37312
rect 16850 37272 16856 37284
rect 16908 37272 16914 37324
rect 17696 37321 17724 37352
rect 19628 37324 19656 37352
rect 17681 37315 17739 37321
rect 16960 37284 17632 37312
rect 16960 37244 16988 37284
rect 16684 37216 16988 37244
rect 1489 37111 1547 37117
rect 1489 37077 1501 37111
rect 1535 37108 1547 37111
rect 2222 37108 2228 37120
rect 1535 37080 2228 37108
rect 1535 37077 1547 37080
rect 1489 37071 1547 37077
rect 2222 37068 2228 37080
rect 2280 37068 2286 37120
rect 10505 37111 10563 37117
rect 10505 37077 10517 37111
rect 10551 37108 10563 37111
rect 10594 37108 10600 37120
rect 10551 37080 10600 37108
rect 10551 37077 10563 37080
rect 10505 37071 10563 37077
rect 10594 37068 10600 37080
rect 10652 37068 10658 37120
rect 14090 37108 14096 37120
rect 14051 37080 14096 37108
rect 14090 37068 14096 37080
rect 14148 37068 14154 37120
rect 17604 37108 17632 37284
rect 17681 37281 17693 37315
rect 17727 37281 17739 37315
rect 17681 37275 17739 37281
rect 17948 37315 18006 37321
rect 17948 37281 17960 37315
rect 17994 37312 18006 37315
rect 18230 37312 18236 37324
rect 17994 37284 18236 37312
rect 17994 37281 18006 37284
rect 17948 37275 18006 37281
rect 18230 37272 18236 37284
rect 18288 37272 18294 37324
rect 19610 37312 19616 37324
rect 19571 37284 19616 37312
rect 19610 37272 19616 37284
rect 19668 37272 19674 37324
rect 19886 37321 19892 37324
rect 19880 37275 19892 37321
rect 19944 37312 19950 37324
rect 20088 37312 20116 37420
rect 20990 37408 20996 37420
rect 21048 37408 21054 37460
rect 21082 37408 21088 37460
rect 21140 37448 21146 37460
rect 21821 37451 21879 37457
rect 21821 37448 21833 37451
rect 21140 37420 21833 37448
rect 21140 37408 21146 37420
rect 21821 37417 21833 37420
rect 21867 37417 21879 37451
rect 21821 37411 21879 37417
rect 21910 37408 21916 37460
rect 21968 37448 21974 37460
rect 22005 37451 22063 37457
rect 22005 37448 22017 37451
rect 21968 37420 22017 37448
rect 21968 37408 21974 37420
rect 22005 37417 22017 37420
rect 22051 37417 22063 37451
rect 22186 37448 22192 37460
rect 22147 37420 22192 37448
rect 22005 37411 22063 37417
rect 22186 37408 22192 37420
rect 22244 37408 22250 37460
rect 22462 37408 22468 37460
rect 22520 37448 22526 37460
rect 23033 37451 23091 37457
rect 23033 37448 23045 37451
rect 22520 37420 23045 37448
rect 22520 37408 22526 37420
rect 23033 37417 23045 37420
rect 23079 37417 23091 37451
rect 23033 37411 23091 37417
rect 24486 37408 24492 37460
rect 24544 37448 24550 37460
rect 25777 37451 25835 37457
rect 25777 37448 25789 37451
rect 24544 37420 25789 37448
rect 24544 37408 24550 37420
rect 25777 37417 25789 37420
rect 25823 37417 25835 37451
rect 26418 37448 26424 37460
rect 26379 37420 26424 37448
rect 25777 37411 25835 37417
rect 26418 37408 26424 37420
rect 26476 37408 26482 37460
rect 27614 37408 27620 37460
rect 27672 37448 27678 37460
rect 29733 37451 29791 37457
rect 29733 37448 29745 37451
rect 27672 37420 29745 37448
rect 27672 37408 27678 37420
rect 29733 37417 29745 37420
rect 29779 37417 29791 37451
rect 29733 37411 29791 37417
rect 30377 37451 30435 37457
rect 30377 37417 30389 37451
rect 30423 37448 30435 37451
rect 30558 37448 30564 37460
rect 30423 37420 30564 37448
rect 30423 37417 30435 37420
rect 30377 37411 30435 37417
rect 30558 37408 30564 37420
rect 30616 37408 30622 37460
rect 31297 37451 31355 37457
rect 31297 37417 31309 37451
rect 31343 37448 31355 37451
rect 32048 37448 32076 37760
rect 32320 37746 33120 37760
rect 31343 37420 32076 37448
rect 31343 37417 31355 37420
rect 31297 37411 31355 37417
rect 21174 37340 21180 37392
rect 21232 37380 21238 37392
rect 22833 37383 22891 37389
rect 21232 37352 22784 37380
rect 21232 37340 21238 37352
rect 19944 37284 19980 37312
rect 20088 37284 21956 37312
rect 19886 37272 19892 37275
rect 19944 37272 19950 37284
rect 21928 37244 21956 37284
rect 22094 37272 22100 37324
rect 22152 37312 22158 37324
rect 22756 37312 22784 37352
rect 22833 37349 22845 37383
rect 22879 37380 22891 37383
rect 23290 37380 23296 37392
rect 22879 37352 23296 37380
rect 22879 37349 22891 37352
rect 22833 37343 22891 37349
rect 23290 37340 23296 37352
rect 23348 37340 23354 37392
rect 23842 37380 23848 37392
rect 23803 37352 23848 37380
rect 23842 37340 23848 37352
rect 23900 37340 23906 37392
rect 24854 37380 24860 37392
rect 24412 37352 24860 37380
rect 24412 37321 24440 37352
rect 24854 37340 24860 37352
rect 24912 37380 24918 37392
rect 26234 37380 26240 37392
rect 24912 37352 26240 37380
rect 24912 37340 24918 37352
rect 26234 37340 26240 37352
rect 26292 37340 26298 37392
rect 27065 37383 27123 37389
rect 27065 37349 27077 37383
rect 27111 37380 27123 37383
rect 27246 37380 27252 37392
rect 27111 37352 27252 37380
rect 27111 37349 27123 37352
rect 27065 37343 27123 37349
rect 27246 37340 27252 37352
rect 27304 37340 27310 37392
rect 27338 37340 27344 37392
rect 27396 37380 27402 37392
rect 27396 37352 27844 37380
rect 27396 37340 27402 37352
rect 23753 37315 23811 37321
rect 23753 37312 23765 37315
rect 22152 37284 22197 37312
rect 22756 37284 23765 37312
rect 22152 37272 22158 37284
rect 23753 37281 23765 37284
rect 23799 37281 23811 37315
rect 23753 37275 23811 37281
rect 24397 37315 24455 37321
rect 24397 37281 24409 37315
rect 24443 37281 24455 37315
rect 24397 37275 24455 37281
rect 24486 37272 24492 37324
rect 24544 37312 24550 37324
rect 24653 37315 24711 37321
rect 24653 37312 24665 37315
rect 24544 37284 24665 37312
rect 24544 37272 24550 37284
rect 24653 37281 24665 37284
rect 24699 37281 24711 37315
rect 24653 37275 24711 37281
rect 27157 37315 27215 37321
rect 27157 37281 27169 37315
rect 27203 37281 27215 37315
rect 27614 37312 27620 37324
rect 27575 37284 27620 37312
rect 27157 37275 27215 37281
rect 23014 37244 23020 37256
rect 21928 37216 23020 37244
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 27062 37204 27068 37256
rect 27120 37244 27126 37256
rect 27172 37244 27200 37275
rect 27614 37272 27620 37284
rect 27672 37272 27678 37324
rect 27816 37321 27844 37352
rect 28092 37352 28672 37380
rect 28092 37324 28120 37352
rect 27801 37315 27859 37321
rect 27801 37281 27813 37315
rect 27847 37281 27859 37315
rect 27801 37275 27859 37281
rect 28074 37272 28080 37324
rect 28132 37272 28138 37324
rect 28166 37272 28172 37324
rect 28224 37312 28230 37324
rect 28644 37321 28672 37352
rect 28353 37315 28411 37321
rect 28353 37312 28365 37315
rect 28224 37284 28365 37312
rect 28224 37272 28230 37284
rect 28353 37281 28365 37284
rect 28399 37281 28411 37315
rect 28353 37275 28411 37281
rect 28629 37315 28687 37321
rect 28629 37281 28641 37315
rect 28675 37281 28687 37315
rect 28629 37275 28687 37281
rect 29825 37315 29883 37321
rect 29825 37281 29837 37315
rect 29871 37312 29883 37315
rect 30742 37312 30748 37324
rect 29871 37284 30748 37312
rect 29871 37281 29883 37284
rect 29825 37275 29883 37281
rect 30742 37272 30748 37284
rect 30800 37272 30806 37324
rect 31110 37312 31116 37324
rect 31071 37284 31116 37312
rect 31110 37272 31116 37284
rect 31168 37272 31174 37324
rect 27120 37216 27200 37244
rect 27120 37204 27126 37216
rect 19058 37176 19064 37188
rect 19019 37148 19064 37176
rect 19058 37136 19064 37148
rect 19116 37136 19122 37188
rect 22370 37176 22376 37188
rect 22283 37148 22376 37176
rect 22370 37136 22376 37148
rect 22428 37176 22434 37188
rect 22922 37176 22928 37188
rect 22428 37148 22928 37176
rect 22428 37136 22434 37148
rect 22922 37136 22928 37148
rect 22980 37136 22986 37188
rect 27522 37176 27528 37188
rect 25332 37148 27528 37176
rect 18322 37108 18328 37120
rect 17604 37080 18328 37108
rect 18322 37068 18328 37080
rect 18380 37068 18386 37120
rect 22738 37068 22744 37120
rect 22796 37108 22802 37120
rect 23017 37111 23075 37117
rect 23017 37108 23029 37111
rect 22796 37080 23029 37108
rect 22796 37068 22802 37080
rect 23017 37077 23029 37080
rect 23063 37077 23075 37111
rect 23198 37108 23204 37120
rect 23159 37080 23204 37108
rect 23017 37071 23075 37077
rect 23198 37068 23204 37080
rect 23256 37068 23262 37120
rect 23382 37068 23388 37120
rect 23440 37108 23446 37120
rect 25332 37108 25360 37148
rect 27522 37136 27528 37148
rect 27580 37136 27586 37188
rect 23440 37080 25360 37108
rect 23440 37068 23446 37080
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27617 37111 27675 37117
rect 27617 37108 27629 37111
rect 26476 37080 27629 37108
rect 26476 37068 26482 37080
rect 27617 37077 27629 37080
rect 27663 37077 27675 37111
rect 27617 37071 27675 37077
rect 1104 37018 32016 37040
rect 1104 36966 6102 37018
rect 6154 36966 6166 37018
rect 6218 36966 6230 37018
rect 6282 36966 6294 37018
rect 6346 36966 6358 37018
rect 6410 36966 16405 37018
rect 16457 36966 16469 37018
rect 16521 36966 16533 37018
rect 16585 36966 16597 37018
rect 16649 36966 16661 37018
rect 16713 36966 26709 37018
rect 26761 36966 26773 37018
rect 26825 36966 26837 37018
rect 26889 36966 26901 37018
rect 26953 36966 26965 37018
rect 27017 36966 32016 37018
rect 1104 36944 32016 36966
rect 7190 36904 7196 36916
rect 7151 36876 7196 36904
rect 7190 36864 7196 36876
rect 7248 36864 7254 36916
rect 7650 36904 7656 36916
rect 7611 36876 7656 36904
rect 7650 36864 7656 36876
rect 7708 36864 7714 36916
rect 9306 36904 9312 36916
rect 8956 36876 9312 36904
rect 3234 36836 3240 36848
rect 1964 36808 3240 36836
rect 1762 36728 1768 36780
rect 1820 36728 1826 36780
rect 1780 36632 1808 36728
rect 1857 36703 1915 36709
rect 1857 36669 1869 36703
rect 1903 36700 1915 36703
rect 1964 36700 1992 36808
rect 3234 36796 3240 36808
rect 3292 36836 3298 36848
rect 4338 36836 4344 36848
rect 3292 36808 4344 36836
rect 3292 36796 3298 36808
rect 4338 36796 4344 36808
rect 4396 36796 4402 36848
rect 7208 36836 7236 36864
rect 7742 36836 7748 36848
rect 7208 36808 7748 36836
rect 7742 36796 7748 36808
rect 7800 36796 7806 36848
rect 2038 36728 2044 36780
rect 2096 36768 2102 36780
rect 4065 36771 4123 36777
rect 4065 36768 4077 36771
rect 2096 36740 4077 36768
rect 2096 36728 2102 36740
rect 4065 36737 4077 36740
rect 4111 36737 4123 36771
rect 5258 36768 5264 36780
rect 5219 36740 5264 36768
rect 4065 36731 4123 36737
rect 5258 36728 5264 36740
rect 5316 36728 5322 36780
rect 2130 36700 2136 36712
rect 1903 36672 1992 36700
rect 2091 36672 2136 36700
rect 1903 36669 1915 36672
rect 1857 36663 1915 36669
rect 2130 36660 2136 36672
rect 2188 36660 2194 36712
rect 2225 36703 2283 36709
rect 2225 36669 2237 36703
rect 2271 36669 2283 36703
rect 2406 36700 2412 36712
rect 2367 36672 2412 36700
rect 2225 36663 2283 36669
rect 2038 36632 2044 36644
rect 1780 36604 2044 36632
rect 2038 36592 2044 36604
rect 2096 36592 2102 36644
rect 2240 36632 2268 36663
rect 2406 36660 2412 36672
rect 2464 36660 2470 36712
rect 3789 36703 3847 36709
rect 3789 36669 3801 36703
rect 3835 36700 3847 36703
rect 3970 36700 3976 36712
rect 3835 36672 3976 36700
rect 3835 36669 3847 36672
rect 3789 36663 3847 36669
rect 3970 36660 3976 36672
rect 4028 36660 4034 36712
rect 8956 36709 8984 36876
rect 9306 36864 9312 36876
rect 9364 36864 9370 36916
rect 9677 36907 9735 36913
rect 9677 36873 9689 36907
rect 9723 36904 9735 36907
rect 9766 36904 9772 36916
rect 9723 36876 9772 36904
rect 9723 36873 9735 36876
rect 9677 36867 9735 36873
rect 9766 36864 9772 36876
rect 9824 36864 9830 36916
rect 11882 36904 11888 36916
rect 11843 36876 11888 36904
rect 11882 36864 11888 36876
rect 11940 36864 11946 36916
rect 19518 36904 19524 36916
rect 16316 36876 19524 36904
rect 9214 36796 9220 36848
rect 9272 36796 9278 36848
rect 9398 36796 9404 36848
rect 9456 36796 9462 36848
rect 12894 36796 12900 36848
rect 12952 36836 12958 36848
rect 14645 36839 14703 36845
rect 14645 36836 14657 36839
rect 12952 36808 14657 36836
rect 12952 36796 12958 36808
rect 14645 36805 14657 36808
rect 14691 36836 14703 36839
rect 16316 36836 16344 36876
rect 19518 36864 19524 36876
rect 19576 36864 19582 36916
rect 19886 36864 19892 36916
rect 19944 36904 19950 36916
rect 19981 36907 20039 36913
rect 19981 36904 19993 36907
rect 19944 36876 19993 36904
rect 19944 36864 19950 36876
rect 19981 36873 19993 36876
rect 20027 36873 20039 36907
rect 19981 36867 20039 36873
rect 20993 36907 21051 36913
rect 20993 36873 21005 36907
rect 21039 36904 21051 36907
rect 21910 36904 21916 36916
rect 21039 36876 21916 36904
rect 21039 36873 21051 36876
rect 20993 36867 21051 36873
rect 21910 36864 21916 36876
rect 21968 36864 21974 36916
rect 22094 36864 22100 36916
rect 22152 36904 22158 36916
rect 23290 36904 23296 36916
rect 22152 36876 22197 36904
rect 23251 36876 23296 36904
rect 22152 36864 22158 36876
rect 23290 36864 23296 36876
rect 23348 36904 23354 36916
rect 23658 36904 23664 36916
rect 23348 36876 23664 36904
rect 23348 36864 23354 36876
rect 23658 36864 23664 36876
rect 23716 36864 23722 36916
rect 25314 36864 25320 36916
rect 25372 36904 25378 36916
rect 30193 36907 30251 36913
rect 30193 36904 30205 36907
rect 25372 36876 30205 36904
rect 25372 36864 25378 36876
rect 30193 36873 30205 36876
rect 30239 36873 30251 36907
rect 30193 36867 30251 36873
rect 14691 36808 16344 36836
rect 14691 36805 14703 36808
rect 14645 36799 14703 36805
rect 17770 36796 17776 36848
rect 17828 36836 17834 36848
rect 19702 36836 19708 36848
rect 17828 36808 19564 36836
rect 17828 36796 17834 36808
rect 9232 36709 9260 36796
rect 9416 36768 9444 36796
rect 12526 36768 12532 36780
rect 9416 36740 9536 36768
rect 8941 36703 8999 36709
rect 8941 36669 8953 36703
rect 8987 36669 8999 36703
rect 8941 36663 8999 36669
rect 9125 36703 9183 36709
rect 9125 36669 9137 36703
rect 9171 36669 9183 36703
rect 9125 36663 9183 36669
rect 9211 36703 9269 36709
rect 9211 36669 9223 36703
rect 9257 36669 9269 36703
rect 9211 36663 9269 36669
rect 9309 36703 9367 36709
rect 9309 36669 9321 36703
rect 9355 36700 9367 36703
rect 9398 36700 9404 36712
rect 9355 36672 9404 36700
rect 9355 36669 9367 36672
rect 9309 36663 9367 36669
rect 2866 36632 2872 36644
rect 2240 36604 2872 36632
rect 2866 36592 2872 36604
rect 2924 36592 2930 36644
rect 5074 36592 5080 36644
rect 5132 36632 5138 36644
rect 5506 36635 5564 36641
rect 5506 36632 5518 36635
rect 5132 36604 5518 36632
rect 5132 36592 5138 36604
rect 5506 36601 5518 36604
rect 5552 36601 5564 36635
rect 5506 36595 5564 36601
rect 8202 36592 8208 36644
rect 8260 36632 8266 36644
rect 9140 36632 9168 36663
rect 9398 36660 9404 36672
rect 9456 36660 9462 36712
rect 9508 36709 9536 36740
rect 12452 36740 12532 36768
rect 9493 36703 9551 36709
rect 9493 36669 9505 36703
rect 9539 36669 9551 36703
rect 9493 36663 9551 36669
rect 10505 36703 10563 36709
rect 10505 36669 10517 36703
rect 10551 36700 10563 36703
rect 11054 36700 11060 36712
rect 10551 36672 11060 36700
rect 10551 36669 10563 36672
rect 10505 36663 10563 36669
rect 11054 36660 11060 36672
rect 11112 36660 11118 36712
rect 12452 36709 12480 36740
rect 12526 36728 12532 36740
rect 12584 36728 12590 36780
rect 12802 36768 12808 36780
rect 12763 36740 12808 36768
rect 12802 36728 12808 36740
rect 12860 36728 12866 36780
rect 14090 36768 14096 36780
rect 13004 36740 14096 36768
rect 12437 36703 12495 36709
rect 12437 36669 12449 36703
rect 12483 36669 12495 36703
rect 12618 36700 12624 36712
rect 12579 36672 12624 36700
rect 12437 36663 12495 36669
rect 12618 36660 12624 36672
rect 12676 36660 12682 36712
rect 12710 36660 12716 36712
rect 12768 36700 12774 36712
rect 13004 36709 13032 36740
rect 14090 36728 14096 36740
rect 14148 36728 14154 36780
rect 12989 36703 13047 36709
rect 12768 36672 12813 36700
rect 12768 36660 12774 36672
rect 12989 36669 13001 36703
rect 13035 36669 13047 36703
rect 12989 36663 13047 36669
rect 13078 36660 13084 36712
rect 13136 36700 13142 36712
rect 16301 36703 16359 36709
rect 16301 36700 16313 36703
rect 13136 36672 16313 36700
rect 13136 36660 13142 36672
rect 16301 36669 16313 36672
rect 16347 36669 16359 36703
rect 16301 36663 16359 36669
rect 16568 36703 16626 36709
rect 16568 36669 16580 36703
rect 16614 36700 16626 36703
rect 16942 36700 16948 36712
rect 16614 36672 16948 36700
rect 16614 36669 16626 36672
rect 16568 36663 16626 36669
rect 16942 36660 16948 36672
rect 17000 36660 17006 36712
rect 17494 36660 17500 36712
rect 17552 36700 17558 36712
rect 19536 36709 19564 36808
rect 19628 36808 19708 36836
rect 19628 36709 19656 36808
rect 19702 36796 19708 36808
rect 19760 36796 19766 36848
rect 21082 36796 21088 36848
rect 21140 36836 21146 36848
rect 21358 36836 21364 36848
rect 21140 36808 21364 36836
rect 21140 36796 21146 36808
rect 21358 36796 21364 36808
rect 21416 36796 21422 36848
rect 24854 36836 24860 36848
rect 22066 36808 24860 36836
rect 22066 36768 22094 36808
rect 24854 36796 24860 36808
rect 24912 36796 24918 36848
rect 26881 36839 26939 36845
rect 26881 36805 26893 36839
rect 26927 36836 26939 36839
rect 28442 36836 28448 36848
rect 26927 36808 28448 36836
rect 26927 36805 26939 36808
rect 26881 36799 26939 36805
rect 28442 36796 28448 36808
rect 28500 36796 28506 36848
rect 20732 36740 22094 36768
rect 19245 36703 19303 36709
rect 19245 36700 19257 36703
rect 17552 36672 19257 36700
rect 17552 36660 17558 36672
rect 19245 36669 19257 36672
rect 19291 36669 19303 36703
rect 19245 36663 19303 36669
rect 19429 36703 19487 36709
rect 19429 36669 19441 36703
rect 19475 36669 19487 36703
rect 19429 36663 19487 36669
rect 19521 36703 19579 36709
rect 19521 36669 19533 36703
rect 19567 36669 19579 36703
rect 19521 36663 19579 36669
rect 19613 36703 19671 36709
rect 19613 36669 19625 36703
rect 19659 36669 19671 36703
rect 19794 36700 19800 36712
rect 19755 36672 19800 36700
rect 19613 36663 19671 36669
rect 10410 36632 10416 36644
rect 8260 36604 9076 36632
rect 9140 36604 10416 36632
rect 8260 36592 8266 36604
rect 1670 36564 1676 36576
rect 1631 36536 1676 36564
rect 1670 36524 1676 36536
rect 1728 36524 1734 36576
rect 3053 36567 3111 36573
rect 3053 36533 3065 36567
rect 3099 36564 3111 36567
rect 3142 36564 3148 36576
rect 3099 36536 3148 36564
rect 3099 36533 3111 36536
rect 3053 36527 3111 36533
rect 3142 36524 3148 36536
rect 3200 36524 3206 36576
rect 6641 36567 6699 36573
rect 6641 36533 6653 36567
rect 6687 36564 6699 36567
rect 7006 36564 7012 36576
rect 6687 36536 7012 36564
rect 6687 36533 6699 36536
rect 6641 36527 6699 36533
rect 7006 36524 7012 36536
rect 7064 36524 7070 36576
rect 8386 36564 8392 36576
rect 8347 36536 8392 36564
rect 8386 36524 8392 36536
rect 8444 36524 8450 36576
rect 9048 36564 9076 36604
rect 10410 36592 10416 36604
rect 10468 36592 10474 36644
rect 10778 36641 10784 36644
rect 10772 36632 10784 36641
rect 10739 36604 10784 36632
rect 10772 36595 10784 36604
rect 10778 36592 10784 36595
rect 10836 36592 10842 36644
rect 14734 36632 14740 36644
rect 13096 36604 14740 36632
rect 13096 36564 13124 36604
rect 14734 36592 14740 36604
rect 14792 36592 14798 36644
rect 9048 36536 13124 36564
rect 13173 36567 13231 36573
rect 13173 36533 13185 36567
rect 13219 36564 13231 36567
rect 13262 36564 13268 36576
rect 13219 36536 13268 36564
rect 13219 36533 13231 36536
rect 13173 36527 13231 36533
rect 13262 36524 13268 36536
rect 13320 36524 13326 36576
rect 14090 36564 14096 36576
rect 14051 36536 14096 36564
rect 14090 36524 14096 36536
rect 14148 36524 14154 36576
rect 15562 36564 15568 36576
rect 15523 36536 15568 36564
rect 15562 36524 15568 36536
rect 15620 36524 15626 36576
rect 17310 36524 17316 36576
rect 17368 36564 17374 36576
rect 17681 36567 17739 36573
rect 17681 36564 17693 36567
rect 17368 36536 17693 36564
rect 17368 36524 17374 36536
rect 17681 36533 17693 36536
rect 17727 36564 17739 36567
rect 17862 36564 17868 36576
rect 17727 36536 17868 36564
rect 17727 36533 17739 36536
rect 17681 36527 17739 36533
rect 17862 36524 17868 36536
rect 17920 36524 17926 36576
rect 18138 36564 18144 36576
rect 18099 36536 18144 36564
rect 18138 36524 18144 36536
rect 18196 36524 18202 36576
rect 19444 36564 19472 36663
rect 19794 36660 19800 36672
rect 19852 36660 19858 36712
rect 20732 36564 20760 36740
rect 22186 36728 22192 36780
rect 22244 36768 22250 36780
rect 22554 36768 22560 36780
rect 22244 36740 22560 36768
rect 22244 36728 22250 36740
rect 22554 36728 22560 36740
rect 22612 36768 22618 36780
rect 23106 36768 23112 36780
rect 22612 36740 23112 36768
rect 22612 36728 22618 36740
rect 23106 36728 23112 36740
rect 23164 36728 23170 36780
rect 23750 36728 23756 36780
rect 23808 36768 23814 36780
rect 24765 36771 24823 36777
rect 24765 36768 24777 36771
rect 23808 36740 24777 36768
rect 23808 36728 23814 36740
rect 24765 36737 24777 36740
rect 24811 36737 24823 36771
rect 24765 36731 24823 36737
rect 27982 36728 27988 36780
rect 28040 36768 28046 36780
rect 28169 36771 28227 36777
rect 28169 36768 28181 36771
rect 28040 36740 28181 36768
rect 28040 36728 28046 36740
rect 28169 36737 28181 36740
rect 28215 36737 28227 36771
rect 28169 36731 28227 36737
rect 21085 36703 21143 36709
rect 21085 36669 21097 36703
rect 21131 36700 21143 36703
rect 21358 36700 21364 36712
rect 21131 36672 21364 36700
rect 21131 36669 21143 36672
rect 21085 36663 21143 36669
rect 21358 36660 21364 36672
rect 21416 36660 21422 36712
rect 22646 36700 22652 36712
rect 21744 36672 22652 36700
rect 21266 36632 21272 36644
rect 21227 36604 21272 36632
rect 21266 36592 21272 36604
rect 21324 36592 21330 36644
rect 21450 36592 21456 36644
rect 21508 36632 21514 36644
rect 21744 36641 21772 36672
rect 22646 36660 22652 36672
rect 22704 36660 22710 36712
rect 22925 36703 22983 36709
rect 22925 36669 22937 36703
rect 22971 36700 22983 36703
rect 23014 36700 23020 36712
rect 22971 36672 23020 36700
rect 22971 36669 22983 36672
rect 22925 36663 22983 36669
rect 23014 36660 23020 36672
rect 23072 36660 23078 36712
rect 23569 36703 23627 36709
rect 23569 36669 23581 36703
rect 23615 36700 23627 36703
rect 23842 36700 23848 36712
rect 23615 36672 23848 36700
rect 23615 36669 23627 36672
rect 23569 36663 23627 36669
rect 23842 36660 23848 36672
rect 23900 36660 23906 36712
rect 24581 36703 24639 36709
rect 24581 36669 24593 36703
rect 24627 36669 24639 36703
rect 24581 36663 24639 36669
rect 26053 36703 26111 36709
rect 26053 36669 26065 36703
rect 26099 36700 26111 36703
rect 26513 36703 26571 36709
rect 26513 36700 26525 36703
rect 26099 36672 26525 36700
rect 26099 36669 26111 36672
rect 26053 36663 26111 36669
rect 26513 36669 26525 36672
rect 26559 36669 26571 36703
rect 26513 36663 26571 36669
rect 21729 36635 21787 36641
rect 21729 36632 21741 36635
rect 21508 36604 21741 36632
rect 21508 36592 21514 36604
rect 21729 36601 21741 36604
rect 21775 36601 21787 36635
rect 21729 36595 21787 36601
rect 21818 36592 21824 36644
rect 21876 36632 21882 36644
rect 21913 36635 21971 36641
rect 21913 36632 21925 36635
rect 21876 36604 21925 36632
rect 21876 36592 21882 36604
rect 21913 36601 21925 36604
rect 21959 36632 21971 36635
rect 22554 36632 22560 36644
rect 21959 36604 22560 36632
rect 21959 36601 21971 36604
rect 21913 36595 21971 36601
rect 22554 36592 22560 36604
rect 22612 36592 22618 36644
rect 23198 36592 23204 36644
rect 23256 36632 23262 36644
rect 23302 36635 23360 36641
rect 23302 36632 23314 36635
rect 23256 36604 23314 36632
rect 23256 36592 23262 36604
rect 23302 36601 23314 36604
rect 23348 36632 23360 36635
rect 24596 36632 24624 36663
rect 26602 36660 26608 36712
rect 26660 36700 26666 36712
rect 26697 36703 26755 36709
rect 26697 36700 26709 36703
rect 26660 36672 26709 36700
rect 26660 36660 26666 36672
rect 26697 36669 26709 36672
rect 26743 36669 26755 36703
rect 26697 36663 26755 36669
rect 26786 36660 26792 36712
rect 26844 36700 26850 36712
rect 26973 36703 27031 36709
rect 26844 36672 26889 36700
rect 26844 36660 26850 36672
rect 26973 36669 26985 36703
rect 27019 36700 27031 36703
rect 27062 36700 27068 36712
rect 27019 36672 27068 36700
rect 27019 36669 27031 36672
rect 26973 36663 27031 36669
rect 27062 36660 27068 36672
rect 27120 36660 27126 36712
rect 27154 36660 27160 36712
rect 27212 36700 27218 36712
rect 27890 36700 27896 36712
rect 27212 36672 27257 36700
rect 27851 36672 27896 36700
rect 27212 36660 27218 36672
rect 27890 36660 27896 36672
rect 27948 36660 27954 36712
rect 28074 36700 28080 36712
rect 28035 36672 28080 36700
rect 28074 36660 28080 36672
rect 28132 36660 28138 36712
rect 28261 36703 28319 36709
rect 28261 36669 28273 36703
rect 28307 36669 28319 36703
rect 28261 36663 28319 36669
rect 28445 36703 28503 36709
rect 28445 36669 28457 36703
rect 28491 36700 28503 36703
rect 29641 36703 29699 36709
rect 29641 36700 29653 36703
rect 28491 36672 29653 36700
rect 28491 36669 28503 36672
rect 28445 36663 28503 36669
rect 29641 36669 29653 36672
rect 29687 36669 29699 36703
rect 29641 36663 29699 36669
rect 29733 36703 29791 36709
rect 29733 36669 29745 36703
rect 29779 36669 29791 36703
rect 29733 36663 29791 36669
rect 23348 36604 24624 36632
rect 23348 36601 23360 36604
rect 23302 36595 23360 36601
rect 27798 36592 27804 36644
rect 27856 36632 27862 36644
rect 28276 36632 28304 36663
rect 27856 36604 28304 36632
rect 27856 36592 27862 36604
rect 29178 36592 29184 36644
rect 29236 36632 29242 36644
rect 29748 36632 29776 36663
rect 29236 36604 29776 36632
rect 29236 36592 29242 36604
rect 19444 36536 20760 36564
rect 22186 36524 22192 36576
rect 22244 36564 22250 36576
rect 24397 36567 24455 36573
rect 24397 36564 24409 36567
rect 22244 36536 24409 36564
rect 22244 36524 22250 36536
rect 24397 36533 24409 36536
rect 24443 36533 24455 36567
rect 24397 36527 24455 36533
rect 24946 36524 24952 36576
rect 25004 36564 25010 36576
rect 25225 36567 25283 36573
rect 25225 36564 25237 36567
rect 25004 36536 25237 36564
rect 25004 36524 25010 36536
rect 25225 36533 25237 36536
rect 25271 36533 25283 36567
rect 25225 36527 25283 36533
rect 25869 36567 25927 36573
rect 25869 36533 25881 36567
rect 25915 36564 25927 36567
rect 26050 36564 26056 36576
rect 25915 36536 26056 36564
rect 25915 36533 25927 36536
rect 25869 36527 25927 36533
rect 26050 36524 26056 36536
rect 26108 36524 26114 36576
rect 27522 36524 27528 36576
rect 27580 36564 27586 36576
rect 28629 36567 28687 36573
rect 28629 36564 28641 36567
rect 27580 36536 28641 36564
rect 27580 36524 27586 36536
rect 28629 36533 28641 36536
rect 28675 36533 28687 36567
rect 30834 36564 30840 36576
rect 30795 36536 30840 36564
rect 28629 36527 28687 36533
rect 30834 36524 30840 36536
rect 30892 36524 30898 36576
rect 1104 36474 32016 36496
rect 1104 36422 11253 36474
rect 11305 36422 11317 36474
rect 11369 36422 11381 36474
rect 11433 36422 11445 36474
rect 11497 36422 11509 36474
rect 11561 36422 21557 36474
rect 21609 36422 21621 36474
rect 21673 36422 21685 36474
rect 21737 36422 21749 36474
rect 21801 36422 21813 36474
rect 21865 36422 32016 36474
rect 1104 36400 32016 36422
rect 5074 36360 5080 36372
rect 5035 36332 5080 36360
rect 5074 36320 5080 36332
rect 5132 36320 5138 36372
rect 6914 36320 6920 36372
rect 6972 36360 6978 36372
rect 7101 36363 7159 36369
rect 7101 36360 7113 36363
rect 6972 36332 7113 36360
rect 6972 36320 6978 36332
rect 7101 36329 7113 36332
rect 7147 36329 7159 36363
rect 7101 36323 7159 36329
rect 8386 36320 8392 36372
rect 8444 36360 8450 36372
rect 10318 36360 10324 36372
rect 8444 36332 10324 36360
rect 8444 36320 8450 36332
rect 10318 36320 10324 36332
rect 10376 36320 10382 36372
rect 10594 36360 10600 36372
rect 10555 36332 10600 36360
rect 10594 36320 10600 36332
rect 10652 36320 10658 36372
rect 10965 36363 11023 36369
rect 10965 36329 10977 36363
rect 11011 36360 11023 36363
rect 11901 36363 11959 36369
rect 11901 36360 11913 36363
rect 11011 36332 11913 36360
rect 11011 36329 11023 36332
rect 10965 36323 11023 36329
rect 11901 36329 11913 36332
rect 11947 36329 11959 36363
rect 17678 36360 17684 36372
rect 11901 36323 11959 36329
rect 15856 36332 17684 36360
rect 3326 36292 3332 36304
rect 1412 36264 3332 36292
rect 1412 36233 1440 36264
rect 3326 36252 3332 36264
rect 3384 36292 3390 36304
rect 3878 36292 3884 36304
rect 3384 36264 3884 36292
rect 3384 36252 3390 36264
rect 3878 36252 3884 36264
rect 3936 36252 3942 36304
rect 4706 36252 4712 36304
rect 4764 36252 4770 36304
rect 7466 36252 7472 36304
rect 7524 36292 7530 36304
rect 7524 36264 7880 36292
rect 7524 36252 7530 36264
rect 1670 36233 1676 36236
rect 1397 36227 1455 36233
rect 1397 36193 1409 36227
rect 1443 36193 1455 36227
rect 1664 36224 1676 36233
rect 1631 36196 1676 36224
rect 1397 36187 1455 36193
rect 1664 36187 1676 36196
rect 1670 36184 1676 36187
rect 1728 36184 1734 36236
rect 3789 36227 3847 36233
rect 3789 36193 3801 36227
rect 3835 36224 3847 36227
rect 3970 36224 3976 36236
rect 3835 36196 3976 36224
rect 3835 36193 3847 36196
rect 3789 36187 3847 36193
rect 3970 36184 3976 36196
rect 4028 36184 4034 36236
rect 4341 36227 4399 36233
rect 4341 36193 4353 36227
rect 4387 36224 4399 36227
rect 4430 36224 4436 36236
rect 4387 36196 4436 36224
rect 4387 36193 4399 36196
rect 4341 36187 4399 36193
rect 4430 36184 4436 36196
rect 4488 36184 4494 36236
rect 4525 36227 4583 36233
rect 4525 36193 4537 36227
rect 4571 36224 4583 36227
rect 4724 36224 4752 36252
rect 4571 36196 4752 36224
rect 4893 36227 4951 36233
rect 4571 36193 4583 36196
rect 4525 36187 4583 36193
rect 4893 36193 4905 36227
rect 4939 36224 4951 36227
rect 6549 36227 6607 36233
rect 4939 36196 5580 36224
rect 4939 36193 4951 36196
rect 4893 36187 4951 36193
rect 5552 36168 5580 36196
rect 6549 36193 6561 36227
rect 6595 36224 6607 36227
rect 6914 36224 6920 36236
rect 6595 36196 6920 36224
rect 6595 36193 6607 36196
rect 6549 36187 6607 36193
rect 6914 36184 6920 36196
rect 6972 36184 6978 36236
rect 7282 36224 7288 36236
rect 7243 36196 7288 36224
rect 7282 36184 7288 36196
rect 7340 36184 7346 36236
rect 7650 36224 7656 36236
rect 7611 36196 7656 36224
rect 7650 36184 7656 36196
rect 7708 36184 7714 36236
rect 7852 36233 7880 36264
rect 10410 36252 10416 36304
rect 10468 36292 10474 36304
rect 10505 36295 10563 36301
rect 10505 36292 10517 36295
rect 10468 36264 10517 36292
rect 10468 36252 10474 36264
rect 10505 36261 10517 36264
rect 10551 36261 10563 36295
rect 10505 36255 10563 36261
rect 11701 36295 11759 36301
rect 11701 36261 11713 36295
rect 11747 36292 11759 36295
rect 11790 36292 11796 36304
rect 11747 36264 11796 36292
rect 11747 36261 11759 36264
rect 11701 36255 11759 36261
rect 11790 36252 11796 36264
rect 11848 36252 11854 36304
rect 15856 36301 15884 36332
rect 17678 36320 17684 36332
rect 17736 36320 17742 36372
rect 18230 36360 18236 36372
rect 18191 36332 18236 36360
rect 18230 36320 18236 36332
rect 18288 36320 18294 36372
rect 21177 36363 21235 36369
rect 21177 36329 21189 36363
rect 21223 36360 21235 36363
rect 21450 36360 21456 36372
rect 21223 36332 21456 36360
rect 21223 36329 21235 36332
rect 21177 36323 21235 36329
rect 21450 36320 21456 36332
rect 21508 36320 21514 36372
rect 26050 36360 26056 36372
rect 26011 36332 26056 36360
rect 26050 36320 26056 36332
rect 26108 36320 26114 36372
rect 26145 36363 26203 36369
rect 26145 36329 26157 36363
rect 26191 36360 26203 36363
rect 26326 36360 26332 36372
rect 26191 36332 26332 36360
rect 26191 36329 26203 36332
rect 26145 36323 26203 36329
rect 26326 36320 26332 36332
rect 26384 36320 26390 36372
rect 26973 36363 27031 36369
rect 26973 36329 26985 36363
rect 27019 36360 27031 36363
rect 27154 36360 27160 36372
rect 27019 36332 27160 36360
rect 27019 36329 27031 36332
rect 26973 36323 27031 36329
rect 27154 36320 27160 36332
rect 27212 36320 27218 36372
rect 15841 36295 15899 36301
rect 15841 36261 15853 36295
rect 15887 36261 15899 36295
rect 15841 36255 15899 36261
rect 17402 36252 17408 36304
rect 17460 36292 17466 36304
rect 17862 36292 17868 36304
rect 17460 36264 17868 36292
rect 17460 36252 17466 36264
rect 17862 36252 17868 36264
rect 17920 36252 17926 36304
rect 21821 36295 21879 36301
rect 21821 36261 21833 36295
rect 21867 36292 21879 36295
rect 22094 36292 22100 36304
rect 21867 36264 22100 36292
rect 21867 36261 21879 36264
rect 21821 36255 21879 36261
rect 22094 36252 22100 36264
rect 22152 36252 22158 36304
rect 22189 36295 22247 36301
rect 22189 36261 22201 36295
rect 22235 36292 22247 36295
rect 22278 36292 22284 36304
rect 22235 36264 22284 36292
rect 22235 36261 22247 36264
rect 22189 36255 22247 36261
rect 22278 36252 22284 36264
rect 22336 36252 22342 36304
rect 23566 36292 23572 36304
rect 23527 36264 23572 36292
rect 23566 36252 23572 36264
rect 23624 36252 23630 36304
rect 24489 36295 24547 36301
rect 24489 36261 24501 36295
rect 24535 36292 24547 36295
rect 26510 36292 26516 36304
rect 24535 36264 26516 36292
rect 24535 36261 24547 36264
rect 24489 36255 24547 36261
rect 26510 36252 26516 36264
rect 26568 36252 26574 36304
rect 27338 36252 27344 36304
rect 27396 36292 27402 36304
rect 29086 36292 29092 36304
rect 27396 36264 27752 36292
rect 27396 36252 27402 36264
rect 7837 36227 7895 36233
rect 7837 36193 7849 36227
rect 7883 36224 7895 36227
rect 8297 36227 8355 36233
rect 8297 36224 8309 36227
rect 7883 36196 8309 36224
rect 7883 36193 7895 36196
rect 7837 36187 7895 36193
rect 8297 36193 8309 36196
rect 8343 36193 8355 36227
rect 9214 36224 9220 36236
rect 9175 36196 9220 36224
rect 8297 36187 8355 36193
rect 9214 36184 9220 36196
rect 9272 36184 9278 36236
rect 12989 36227 13047 36233
rect 12989 36193 13001 36227
rect 13035 36224 13047 36227
rect 13078 36224 13084 36236
rect 13035 36196 13084 36224
rect 13035 36193 13047 36196
rect 12989 36187 13047 36193
rect 13078 36184 13084 36196
rect 13136 36184 13142 36236
rect 13262 36233 13268 36236
rect 13256 36224 13268 36233
rect 13223 36196 13268 36224
rect 13256 36187 13268 36196
rect 13262 36184 13268 36187
rect 13320 36184 13326 36236
rect 15010 36184 15016 36236
rect 15068 36224 15074 36236
rect 15565 36227 15623 36233
rect 15565 36224 15577 36227
rect 15068 36196 15577 36224
rect 15068 36184 15074 36196
rect 15565 36193 15577 36196
rect 15611 36193 15623 36227
rect 15565 36187 15623 36193
rect 15933 36227 15991 36233
rect 15933 36193 15945 36227
rect 15979 36193 15991 36227
rect 15933 36187 15991 36193
rect 16853 36227 16911 36233
rect 16853 36193 16865 36227
rect 16899 36224 16911 36227
rect 17218 36224 17224 36236
rect 16899 36196 17224 36224
rect 16899 36193 16911 36196
rect 16853 36187 16911 36193
rect 4246 36116 4252 36168
rect 4304 36156 4310 36168
rect 4617 36159 4675 36165
rect 4617 36156 4629 36159
rect 4304 36128 4629 36156
rect 4304 36116 4310 36128
rect 4617 36125 4629 36128
rect 4663 36125 4675 36159
rect 4617 36119 4675 36125
rect 4709 36159 4767 36165
rect 4709 36125 4721 36159
rect 4755 36125 4767 36159
rect 4709 36119 4767 36125
rect 3418 36088 3424 36100
rect 2332 36060 3424 36088
rect 2130 35980 2136 36032
rect 2188 36020 2194 36032
rect 2332 36020 2360 36060
rect 3418 36048 3424 36060
rect 3476 36048 3482 36100
rect 4724 36088 4752 36119
rect 5534 36116 5540 36168
rect 5592 36156 5598 36168
rect 6365 36159 6423 36165
rect 6365 36156 6377 36159
rect 5592 36128 6377 36156
rect 5592 36116 5598 36128
rect 6365 36125 6377 36128
rect 6411 36125 6423 36159
rect 6365 36119 6423 36125
rect 7374 36116 7380 36168
rect 7432 36156 7438 36168
rect 7469 36159 7527 36165
rect 7469 36156 7481 36159
rect 7432 36128 7481 36156
rect 7432 36116 7438 36128
rect 7469 36125 7481 36128
rect 7515 36125 7527 36159
rect 7469 36119 7527 36125
rect 7561 36159 7619 36165
rect 7561 36125 7573 36159
rect 7607 36125 7619 36159
rect 7561 36119 7619 36125
rect 8941 36159 8999 36165
rect 8941 36125 8953 36159
rect 8987 36156 8999 36159
rect 8987 36128 9260 36156
rect 8987 36125 8999 36128
rect 8941 36119 8999 36125
rect 4172 36060 4752 36088
rect 4172 36032 4200 36060
rect 7282 36048 7288 36100
rect 7340 36088 7346 36100
rect 7576 36088 7604 36119
rect 9232 36100 9260 36128
rect 10226 36116 10232 36168
rect 10284 36156 10290 36168
rect 10321 36159 10379 36165
rect 10321 36156 10333 36159
rect 10284 36128 10333 36156
rect 10284 36116 10290 36128
rect 10321 36125 10333 36128
rect 10367 36125 10379 36159
rect 15470 36156 15476 36168
rect 15431 36128 15476 36156
rect 10321 36119 10379 36125
rect 15470 36116 15476 36128
rect 15528 36116 15534 36168
rect 15948 36156 15976 36187
rect 17218 36184 17224 36196
rect 17276 36184 17282 36236
rect 17494 36224 17500 36236
rect 17455 36196 17500 36224
rect 17494 36184 17500 36196
rect 17552 36184 17558 36236
rect 17681 36227 17739 36233
rect 17681 36193 17693 36227
rect 17727 36193 17739 36227
rect 17681 36187 17739 36193
rect 17037 36159 17095 36165
rect 15948 36128 16988 36156
rect 7340 36060 7604 36088
rect 7340 36048 7346 36060
rect 9214 36048 9220 36100
rect 9272 36048 9278 36100
rect 12894 36088 12900 36100
rect 11900 36060 12900 36088
rect 2188 35992 2360 36020
rect 2188 35980 2194 35992
rect 2774 35980 2780 36032
rect 2832 36020 2838 36032
rect 3697 36023 3755 36029
rect 2832 35992 2877 36020
rect 2832 35980 2838 35992
rect 3697 35989 3709 36023
rect 3743 36020 3755 36023
rect 3786 36020 3792 36032
rect 3743 35992 3792 36020
rect 3743 35989 3755 35992
rect 3697 35983 3755 35989
rect 3786 35980 3792 35992
rect 3844 36020 3850 36032
rect 4154 36020 4160 36032
rect 3844 35992 4160 36020
rect 3844 35980 3850 35992
rect 4154 35980 4160 35992
rect 4212 35980 4218 36032
rect 5166 35980 5172 36032
rect 5224 36020 5230 36032
rect 11900 36029 11928 36060
rect 12894 36048 12900 36060
rect 12952 36048 12958 36100
rect 5537 36023 5595 36029
rect 5537 36020 5549 36023
rect 5224 35992 5549 36020
rect 5224 35980 5230 35992
rect 5537 35989 5549 35992
rect 5583 35989 5595 36023
rect 5537 35983 5595 35989
rect 11885 36023 11943 36029
rect 11885 35989 11897 36023
rect 11931 35989 11943 36023
rect 11885 35983 11943 35989
rect 11974 35980 11980 36032
rect 12032 36020 12038 36032
rect 12069 36023 12127 36029
rect 12069 36020 12081 36023
rect 12032 35992 12081 36020
rect 12032 35980 12038 35992
rect 12069 35989 12081 35992
rect 12115 35989 12127 36023
rect 12069 35983 12127 35989
rect 13722 35980 13728 36032
rect 13780 36020 13786 36032
rect 14090 36020 14096 36032
rect 13780 35992 14096 36020
rect 13780 35980 13786 35992
rect 14090 35980 14096 35992
rect 14148 36020 14154 36032
rect 14369 36023 14427 36029
rect 14369 36020 14381 36023
rect 14148 35992 14381 36020
rect 14148 35980 14154 35992
rect 14369 35989 14381 35992
rect 14415 35989 14427 36023
rect 14369 35983 14427 35989
rect 16669 36023 16727 36029
rect 16669 35989 16681 36023
rect 16715 36020 16727 36023
rect 16850 36020 16856 36032
rect 16715 35992 16856 36020
rect 16715 35989 16727 35992
rect 16669 35983 16727 35989
rect 16850 35980 16856 35992
rect 16908 35980 16914 36032
rect 16960 36020 16988 36128
rect 17037 36125 17049 36159
rect 17083 36156 17095 36159
rect 17696 36156 17724 36187
rect 17770 36184 17776 36236
rect 17828 36224 17834 36236
rect 17828 36196 17873 36224
rect 17828 36184 17834 36196
rect 17954 36184 17960 36236
rect 18012 36224 18018 36236
rect 18049 36227 18107 36233
rect 18049 36224 18061 36227
rect 18012 36196 18061 36224
rect 18012 36184 18018 36196
rect 18049 36193 18061 36196
rect 18095 36193 18107 36227
rect 18049 36187 18107 36193
rect 21269 36227 21327 36233
rect 21269 36193 21281 36227
rect 21315 36224 21327 36227
rect 21358 36224 21364 36236
rect 21315 36196 21364 36224
rect 21315 36193 21327 36196
rect 21269 36187 21327 36193
rect 21358 36184 21364 36196
rect 21416 36184 21422 36236
rect 21450 36184 21456 36236
rect 21508 36224 21514 36236
rect 21965 36227 22023 36233
rect 21965 36224 21977 36227
rect 21508 36196 21977 36224
rect 21508 36184 21514 36196
rect 21965 36193 21977 36196
rect 22011 36193 22023 36227
rect 21965 36187 22023 36193
rect 23201 36227 23259 36233
rect 23201 36193 23213 36227
rect 23247 36224 23259 36227
rect 23290 36224 23296 36236
rect 23247 36196 23296 36224
rect 23247 36193 23259 36196
rect 23201 36187 23259 36193
rect 23290 36184 23296 36196
rect 23348 36184 23354 36236
rect 23934 36184 23940 36236
rect 23992 36224 23998 36236
rect 24305 36227 24363 36233
rect 24305 36224 24317 36227
rect 23992 36196 24317 36224
rect 23992 36184 23998 36196
rect 24305 36193 24317 36196
rect 24351 36193 24363 36227
rect 24305 36187 24363 36193
rect 26050 36184 26056 36236
rect 26108 36224 26114 36236
rect 27157 36227 27215 36233
rect 27157 36224 27169 36227
rect 26108 36196 27169 36224
rect 26108 36184 26114 36196
rect 27157 36193 27169 36196
rect 27203 36193 27215 36227
rect 27430 36224 27436 36236
rect 27391 36196 27436 36224
rect 27157 36187 27215 36193
rect 27430 36184 27436 36196
rect 27488 36184 27494 36236
rect 27614 36224 27620 36236
rect 27575 36196 27620 36224
rect 27614 36184 27620 36196
rect 27672 36184 27678 36236
rect 17862 36156 17868 36168
rect 17083 36128 17724 36156
rect 17823 36128 17868 36156
rect 17083 36125 17095 36128
rect 17037 36119 17095 36125
rect 17696 36088 17724 36128
rect 17862 36116 17868 36128
rect 17920 36116 17926 36168
rect 18785 36159 18843 36165
rect 18785 36125 18797 36159
rect 18831 36156 18843 36159
rect 20162 36156 20168 36168
rect 18831 36128 20168 36156
rect 18831 36125 18843 36128
rect 18785 36119 18843 36125
rect 18046 36088 18052 36100
rect 17696 36060 18052 36088
rect 18046 36048 18052 36060
rect 18104 36048 18110 36100
rect 18800 36020 18828 36119
rect 20162 36116 20168 36128
rect 20220 36156 20226 36168
rect 21174 36156 21180 36168
rect 20220 36128 21180 36156
rect 20220 36116 20226 36128
rect 21174 36116 21180 36128
rect 21232 36116 21238 36168
rect 26329 36159 26387 36165
rect 26329 36125 26341 36159
rect 26375 36156 26387 36159
rect 26418 36156 26424 36168
rect 26375 36128 26424 36156
rect 26375 36125 26387 36128
rect 26329 36119 26387 36125
rect 26418 36116 26424 36128
rect 26476 36116 26482 36168
rect 27338 36156 27344 36168
rect 27299 36128 27344 36156
rect 27338 36116 27344 36128
rect 27396 36116 27402 36168
rect 18874 36048 18880 36100
rect 18932 36088 18938 36100
rect 22002 36088 22008 36100
rect 18932 36060 22008 36088
rect 18932 36048 18938 36060
rect 22002 36048 22008 36060
rect 22060 36048 22066 36100
rect 24486 36048 24492 36100
rect 24544 36088 24550 36100
rect 26786 36088 26792 36100
rect 24544 36060 26792 36088
rect 24544 36048 24550 36060
rect 26786 36048 26792 36060
rect 26844 36088 26850 36100
rect 27249 36091 27307 36097
rect 27249 36088 27261 36091
rect 26844 36060 27261 36088
rect 26844 36048 26850 36060
rect 27249 36057 27261 36060
rect 27295 36057 27307 36091
rect 27724 36088 27752 36264
rect 28368 36264 29092 36292
rect 28368 36233 28396 36264
rect 29086 36252 29092 36264
rect 29144 36252 29150 36304
rect 28261 36227 28319 36233
rect 28261 36193 28273 36227
rect 28307 36193 28319 36227
rect 28261 36187 28319 36193
rect 28353 36227 28411 36233
rect 28353 36193 28365 36227
rect 28399 36193 28411 36227
rect 28353 36187 28411 36193
rect 28629 36227 28687 36233
rect 28629 36193 28641 36227
rect 28675 36224 28687 36227
rect 29181 36227 29239 36233
rect 29181 36224 29193 36227
rect 28675 36196 29193 36224
rect 28675 36193 28687 36196
rect 28629 36187 28687 36193
rect 29181 36193 29193 36196
rect 29227 36193 29239 36227
rect 29181 36187 29239 36193
rect 29273 36227 29331 36233
rect 29273 36193 29285 36227
rect 29319 36224 29331 36227
rect 30098 36224 30104 36236
rect 29319 36196 30104 36224
rect 29319 36193 29331 36196
rect 29273 36187 29331 36193
rect 28276 36156 28304 36187
rect 30098 36184 30104 36196
rect 30156 36184 30162 36236
rect 30742 36184 30748 36236
rect 30800 36224 30806 36236
rect 31113 36227 31171 36233
rect 31113 36224 31125 36227
rect 30800 36196 31125 36224
rect 30800 36184 30806 36196
rect 31113 36193 31125 36196
rect 31159 36193 31171 36227
rect 31113 36187 31171 36193
rect 29914 36156 29920 36168
rect 28276 36128 29920 36156
rect 29914 36116 29920 36128
rect 29972 36116 29978 36168
rect 28537 36091 28595 36097
rect 28537 36088 28549 36091
rect 27724 36060 28549 36088
rect 27249 36051 27307 36057
rect 28537 36057 28549 36060
rect 28583 36057 28595 36091
rect 28537 36051 28595 36057
rect 16960 35992 18828 36020
rect 19150 35980 19156 36032
rect 19208 36020 19214 36032
rect 19245 36023 19303 36029
rect 19245 36020 19257 36023
rect 19208 35992 19257 36020
rect 19208 35980 19214 35992
rect 19245 35989 19257 35992
rect 19291 35989 19303 36023
rect 19245 35983 19303 35989
rect 20349 36023 20407 36029
rect 20349 35989 20361 36023
rect 20395 36020 20407 36023
rect 20806 36020 20812 36032
rect 20395 35992 20812 36020
rect 20395 35989 20407 35992
rect 20349 35983 20407 35989
rect 20806 35980 20812 35992
rect 20864 35980 20870 36032
rect 22738 36020 22744 36032
rect 22699 35992 22744 36020
rect 22738 35980 22744 35992
rect 22796 35980 22802 36032
rect 23014 35980 23020 36032
rect 23072 36020 23078 36032
rect 23569 36023 23627 36029
rect 23569 36020 23581 36023
rect 23072 35992 23581 36020
rect 23072 35980 23078 35992
rect 23569 35989 23581 35992
rect 23615 35989 23627 36023
rect 23569 35983 23627 35989
rect 23658 35980 23664 36032
rect 23716 36020 23722 36032
rect 23753 36023 23811 36029
rect 23753 36020 23765 36023
rect 23716 35992 23765 36020
rect 23716 35980 23722 35992
rect 23753 35989 23765 35992
rect 23799 35989 23811 36023
rect 25130 36020 25136 36032
rect 25091 35992 25136 36020
rect 23753 35983 23811 35989
rect 25130 35980 25136 35992
rect 25188 35980 25194 36032
rect 25498 35980 25504 36032
rect 25556 36020 25562 36032
rect 25685 36023 25743 36029
rect 25685 36020 25697 36023
rect 25556 35992 25697 36020
rect 25556 35980 25562 35992
rect 25685 35989 25697 35992
rect 25731 35989 25743 36023
rect 25685 35983 25743 35989
rect 28077 36023 28135 36029
rect 28077 35989 28089 36023
rect 28123 36020 28135 36023
rect 28258 36020 28264 36032
rect 28123 35992 28264 36020
rect 28123 35989 28135 35992
rect 28077 35983 28135 35989
rect 28258 35980 28264 35992
rect 28316 35980 28322 36032
rect 29730 36020 29736 36032
rect 29691 35992 29736 36020
rect 29730 35980 29736 35992
rect 29788 35980 29794 36032
rect 30374 36020 30380 36032
rect 30335 35992 30380 36020
rect 30374 35980 30380 35992
rect 30432 36020 30438 36032
rect 30650 36020 30656 36032
rect 30432 35992 30656 36020
rect 30432 35980 30438 35992
rect 30650 35980 30656 35992
rect 30708 35980 30714 36032
rect 31297 36023 31355 36029
rect 31297 35989 31309 36023
rect 31343 36020 31355 36023
rect 31343 35992 32076 36020
rect 31343 35989 31355 35992
rect 31297 35983 31355 35989
rect 1104 35930 32016 35952
rect 1104 35878 6102 35930
rect 6154 35878 6166 35930
rect 6218 35878 6230 35930
rect 6282 35878 6294 35930
rect 6346 35878 6358 35930
rect 6410 35878 16405 35930
rect 16457 35878 16469 35930
rect 16521 35878 16533 35930
rect 16585 35878 16597 35930
rect 16649 35878 16661 35930
rect 16713 35878 26709 35930
rect 26761 35878 26773 35930
rect 26825 35878 26837 35930
rect 26889 35878 26901 35930
rect 26953 35878 26965 35930
rect 27017 35878 32016 35930
rect 1104 35856 32016 35878
rect 1581 35819 1639 35825
rect 1581 35785 1593 35819
rect 1627 35816 1639 35819
rect 5442 35816 5448 35828
rect 1627 35788 5448 35816
rect 1627 35785 1639 35788
rect 1581 35779 1639 35785
rect 5442 35776 5448 35788
rect 5500 35776 5506 35828
rect 17773 35819 17831 35825
rect 9876 35788 16988 35816
rect 0 35748 800 35762
rect 3050 35748 3056 35760
rect 0 35720 3056 35748
rect 0 35706 800 35720
rect 3050 35708 3056 35720
rect 3108 35708 3114 35760
rect 3970 35708 3976 35760
rect 4028 35748 4034 35760
rect 4028 35720 5948 35748
rect 4028 35708 4034 35720
rect 5920 35692 5948 35720
rect 6730 35708 6736 35760
rect 6788 35748 6794 35760
rect 9490 35748 9496 35760
rect 6788 35720 9496 35748
rect 6788 35708 6794 35720
rect 9490 35708 9496 35720
rect 9548 35708 9554 35760
rect 2406 35640 2412 35692
rect 2464 35680 2470 35692
rect 2593 35683 2651 35689
rect 2593 35680 2605 35683
rect 2464 35652 2605 35680
rect 2464 35640 2470 35652
rect 2593 35649 2605 35652
rect 2639 35649 2651 35683
rect 4246 35680 4252 35692
rect 4207 35652 4252 35680
rect 2593 35643 2651 35649
rect 4246 35640 4252 35652
rect 4304 35640 4310 35692
rect 5718 35680 5724 35692
rect 4356 35652 5724 35680
rect 2869 35615 2927 35621
rect 2869 35581 2881 35615
rect 2915 35612 2927 35615
rect 3142 35612 3148 35624
rect 2915 35584 3148 35612
rect 2915 35581 2927 35584
rect 2869 35575 2927 35581
rect 3142 35572 3148 35584
rect 3200 35612 3206 35624
rect 3973 35615 4031 35621
rect 3200 35584 3924 35612
rect 3200 35572 3206 35584
rect 3602 35436 3608 35488
rect 3660 35476 3666 35488
rect 3789 35479 3847 35485
rect 3789 35476 3801 35479
rect 3660 35448 3801 35476
rect 3660 35436 3666 35448
rect 3789 35445 3801 35448
rect 3835 35445 3847 35479
rect 3896 35476 3924 35584
rect 3973 35581 3985 35615
rect 4019 35581 4031 35615
rect 4154 35612 4160 35624
rect 4115 35584 4160 35612
rect 3973 35575 4031 35581
rect 3988 35544 4016 35575
rect 4154 35572 4160 35584
rect 4212 35572 4218 35624
rect 4356 35621 4384 35652
rect 5718 35640 5724 35652
rect 5776 35640 5782 35692
rect 5902 35640 5908 35692
rect 5960 35680 5966 35692
rect 6825 35683 6883 35689
rect 6825 35680 6837 35683
rect 5960 35652 6837 35680
rect 5960 35640 5966 35652
rect 6825 35649 6837 35652
rect 6871 35649 6883 35683
rect 6825 35643 6883 35649
rect 7374 35640 7380 35692
rect 7432 35640 7438 35692
rect 4341 35615 4399 35621
rect 4341 35581 4353 35615
rect 4387 35581 4399 35615
rect 4341 35575 4399 35581
rect 4430 35572 4436 35624
rect 4488 35612 4494 35624
rect 4525 35615 4583 35621
rect 4525 35612 4537 35615
rect 4488 35584 4537 35612
rect 4488 35572 4494 35584
rect 4525 35581 4537 35584
rect 4571 35612 4583 35615
rect 5074 35612 5080 35624
rect 4571 35584 5080 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 5074 35572 5080 35584
rect 5132 35572 5138 35624
rect 6365 35615 6423 35621
rect 6365 35581 6377 35615
rect 6411 35612 6423 35615
rect 6454 35612 6460 35624
rect 6411 35584 6460 35612
rect 6411 35581 6423 35584
rect 6365 35575 6423 35581
rect 6454 35572 6460 35584
rect 6512 35572 6518 35624
rect 7101 35615 7159 35621
rect 7101 35581 7113 35615
rect 7147 35612 7159 35615
rect 7392 35612 7420 35640
rect 7926 35612 7932 35624
rect 7147 35584 7932 35612
rect 7147 35581 7159 35584
rect 7101 35575 7159 35581
rect 7926 35572 7932 35584
rect 7984 35572 7990 35624
rect 9876 35621 9904 35788
rect 9953 35683 10011 35689
rect 9953 35649 9965 35683
rect 9999 35680 10011 35683
rect 10318 35680 10324 35692
rect 9999 35652 10324 35680
rect 9999 35649 10011 35652
rect 9953 35643 10011 35649
rect 10318 35640 10324 35652
rect 10376 35640 10382 35692
rect 11793 35683 11851 35689
rect 11793 35649 11805 35683
rect 11839 35680 11851 35683
rect 11882 35680 11888 35692
rect 11839 35652 11888 35680
rect 11839 35649 11851 35652
rect 11793 35643 11851 35649
rect 11882 35640 11888 35652
rect 11940 35640 11946 35692
rect 12989 35683 13047 35689
rect 12989 35649 13001 35683
rect 13035 35680 13047 35683
rect 13446 35680 13452 35692
rect 13035 35652 13452 35680
rect 13035 35649 13047 35652
rect 12989 35643 13047 35649
rect 13446 35640 13452 35652
rect 13504 35680 13510 35692
rect 13504 35652 15056 35680
rect 13504 35640 13510 35652
rect 8113 35615 8171 35621
rect 8113 35581 8125 35615
rect 8159 35581 8171 35615
rect 8113 35575 8171 35581
rect 9677 35615 9735 35621
rect 9677 35581 9689 35615
rect 9723 35581 9735 35615
rect 9677 35575 9735 35581
rect 9861 35615 9919 35621
rect 9861 35581 9873 35615
rect 9907 35581 9919 35615
rect 9861 35575 9919 35581
rect 10045 35615 10103 35621
rect 10045 35581 10057 35615
rect 10091 35612 10103 35615
rect 10134 35612 10140 35624
rect 10091 35584 10140 35612
rect 10091 35581 10103 35584
rect 10045 35575 10103 35581
rect 4706 35544 4712 35556
rect 3988 35516 4712 35544
rect 4706 35504 4712 35516
rect 4764 35504 4770 35556
rect 5166 35544 5172 35556
rect 4816 35516 5172 35544
rect 4154 35476 4160 35488
rect 3896 35448 4160 35476
rect 3789 35439 3847 35445
rect 4154 35436 4160 35448
rect 4212 35476 4218 35488
rect 4816 35476 4844 35516
rect 5166 35504 5172 35516
rect 5224 35504 5230 35556
rect 6914 35504 6920 35556
rect 6972 35544 6978 35556
rect 8128 35544 8156 35575
rect 6972 35516 8156 35544
rect 9692 35544 9720 35575
rect 10134 35572 10140 35584
rect 10192 35572 10198 35624
rect 10226 35572 10232 35624
rect 10284 35612 10290 35624
rect 10410 35612 10416 35624
rect 10284 35584 10416 35612
rect 10284 35572 10290 35584
rect 10410 35572 10416 35584
rect 10468 35572 10474 35624
rect 11974 35612 11980 35624
rect 11935 35584 11980 35612
rect 11974 35572 11980 35584
rect 12032 35612 12038 35624
rect 13173 35615 13231 35621
rect 13173 35612 13185 35615
rect 12032 35584 13185 35612
rect 12032 35572 12038 35584
rect 13173 35581 13185 35584
rect 13219 35581 13231 35615
rect 14366 35612 14372 35624
rect 14327 35584 14372 35612
rect 13173 35575 13231 35581
rect 14366 35572 14372 35584
rect 14424 35572 14430 35624
rect 10594 35544 10600 35556
rect 9692 35516 10600 35544
rect 6972 35504 6978 35516
rect 10594 35504 10600 35516
rect 10652 35544 10658 35556
rect 11146 35544 11152 35556
rect 10652 35516 11152 35544
rect 10652 35504 10658 35516
rect 11146 35504 11152 35516
rect 11204 35504 11210 35556
rect 12618 35504 12624 35556
rect 12676 35544 12682 35556
rect 13538 35544 13544 35556
rect 12676 35516 13308 35544
rect 13499 35516 13544 35544
rect 12676 35504 12682 35516
rect 5074 35476 5080 35488
rect 4212 35448 4844 35476
rect 5035 35448 5080 35476
rect 4212 35436 4218 35448
rect 5074 35436 5080 35448
rect 5132 35436 5138 35488
rect 6273 35479 6331 35485
rect 6273 35445 6285 35479
rect 6319 35476 6331 35479
rect 7190 35476 7196 35488
rect 6319 35448 7196 35476
rect 6319 35445 6331 35448
rect 6273 35439 6331 35445
rect 7190 35436 7196 35448
rect 7248 35436 7254 35488
rect 7282 35436 7288 35488
rect 7340 35476 7346 35488
rect 8205 35479 8263 35485
rect 8205 35476 8217 35479
rect 7340 35448 8217 35476
rect 7340 35436 7346 35448
rect 8205 35445 8217 35448
rect 8251 35445 8263 35479
rect 9214 35476 9220 35488
rect 9175 35448 9220 35476
rect 8205 35439 8263 35445
rect 9214 35436 9220 35448
rect 9272 35436 9278 35488
rect 9398 35436 9404 35488
rect 9456 35476 9462 35488
rect 10134 35476 10140 35488
rect 9456 35448 10140 35476
rect 9456 35436 9462 35448
rect 10134 35436 10140 35448
rect 10192 35436 10198 35488
rect 10410 35476 10416 35488
rect 10371 35448 10416 35476
rect 10410 35436 10416 35448
rect 10468 35436 10474 35488
rect 10870 35476 10876 35488
rect 10831 35448 10876 35476
rect 10870 35436 10876 35448
rect 10928 35436 10934 35488
rect 12158 35476 12164 35488
rect 12119 35448 12164 35476
rect 12158 35436 12164 35448
rect 12216 35436 12222 35488
rect 13280 35485 13308 35516
rect 13538 35504 13544 35516
rect 13596 35504 13602 35556
rect 14277 35547 14335 35553
rect 14277 35513 14289 35547
rect 14323 35544 14335 35547
rect 14918 35544 14924 35556
rect 14323 35516 14924 35544
rect 14323 35513 14335 35516
rect 14277 35507 14335 35513
rect 14918 35504 14924 35516
rect 14976 35504 14982 35556
rect 13265 35479 13323 35485
rect 13265 35445 13277 35479
rect 13311 35445 13323 35479
rect 13265 35439 13323 35445
rect 13357 35479 13415 35485
rect 13357 35445 13369 35479
rect 13403 35476 13415 35479
rect 14090 35476 14096 35488
rect 13403 35448 14096 35476
rect 13403 35445 13415 35448
rect 13357 35439 13415 35445
rect 14090 35436 14096 35448
rect 14148 35436 14154 35488
rect 14366 35436 14372 35488
rect 14424 35476 14430 35488
rect 14829 35479 14887 35485
rect 14829 35476 14841 35479
rect 14424 35448 14841 35476
rect 14424 35436 14430 35448
rect 14829 35445 14841 35448
rect 14875 35445 14887 35479
rect 15028 35476 15056 35652
rect 15102 35572 15108 35624
rect 15160 35612 15166 35624
rect 16209 35615 16267 35621
rect 16209 35612 16221 35615
rect 15160 35584 16221 35612
rect 15160 35572 15166 35584
rect 16209 35581 16221 35584
rect 16255 35581 16267 35615
rect 16209 35575 16267 35581
rect 16761 35615 16819 35621
rect 16761 35581 16773 35615
rect 16807 35612 16819 35615
rect 16850 35612 16856 35624
rect 16807 35584 16856 35612
rect 16807 35581 16819 35584
rect 16761 35575 16819 35581
rect 16850 35572 16856 35584
rect 16908 35572 16914 35624
rect 16960 35612 16988 35788
rect 17773 35785 17785 35819
rect 17819 35816 17831 35819
rect 17954 35816 17960 35828
rect 17819 35788 17960 35816
rect 17819 35785 17831 35788
rect 17773 35779 17831 35785
rect 17954 35776 17960 35788
rect 18012 35776 18018 35828
rect 19242 35816 19248 35828
rect 18064 35788 19248 35816
rect 17862 35708 17868 35760
rect 17920 35748 17926 35760
rect 18064 35748 18092 35788
rect 19242 35776 19248 35788
rect 19300 35776 19306 35828
rect 19518 35776 19524 35828
rect 19576 35816 19582 35828
rect 19576 35788 20208 35816
rect 19576 35776 19582 35788
rect 17920 35720 18092 35748
rect 17920 35708 17926 35720
rect 18322 35708 18328 35760
rect 18380 35748 18386 35760
rect 20180 35748 20208 35788
rect 21266 35776 21272 35828
rect 21324 35816 21330 35828
rect 21361 35819 21419 35825
rect 21361 35816 21373 35819
rect 21324 35788 21373 35816
rect 21324 35776 21330 35788
rect 21361 35785 21373 35788
rect 21407 35785 21419 35819
rect 21361 35779 21419 35785
rect 21542 35776 21548 35828
rect 21600 35816 21606 35828
rect 27154 35816 27160 35828
rect 21600 35788 27160 35816
rect 21600 35776 21606 35788
rect 27154 35776 27160 35788
rect 27212 35776 27218 35828
rect 27338 35776 27344 35828
rect 27396 35816 27402 35828
rect 27525 35819 27583 35825
rect 27525 35816 27537 35819
rect 27396 35788 27537 35816
rect 27396 35776 27402 35788
rect 27525 35785 27537 35788
rect 27571 35785 27583 35819
rect 27525 35779 27583 35785
rect 28074 35776 28080 35828
rect 28132 35816 28138 35828
rect 28813 35819 28871 35825
rect 28813 35816 28825 35819
rect 28132 35788 28825 35816
rect 28132 35776 28138 35788
rect 28813 35785 28825 35788
rect 28859 35785 28871 35819
rect 28813 35779 28871 35785
rect 23198 35748 23204 35760
rect 18380 35720 19288 35748
rect 20180 35720 23204 35748
rect 18380 35708 18386 35720
rect 17494 35640 17500 35692
rect 17552 35680 17558 35692
rect 18509 35683 18567 35689
rect 18509 35680 18521 35683
rect 17552 35652 18521 35680
rect 17552 35640 17558 35652
rect 18509 35649 18521 35652
rect 18555 35649 18567 35683
rect 19260 35680 19288 35720
rect 23198 35708 23204 35720
rect 23256 35748 23262 35760
rect 24946 35748 24952 35760
rect 23256 35720 24952 35748
rect 23256 35708 23262 35720
rect 23400 35689 23428 35720
rect 24946 35708 24952 35720
rect 25004 35708 25010 35760
rect 26697 35751 26755 35757
rect 26697 35717 26709 35751
rect 26743 35748 26755 35751
rect 27614 35748 27620 35760
rect 26743 35720 27620 35748
rect 26743 35717 26755 35720
rect 26697 35711 26755 35717
rect 27614 35708 27620 35720
rect 27672 35708 27678 35760
rect 27706 35708 27712 35760
rect 27764 35748 27770 35760
rect 27890 35748 27896 35760
rect 27764 35720 27896 35748
rect 27764 35708 27770 35720
rect 27890 35708 27896 35720
rect 27948 35708 27954 35760
rect 28994 35708 29000 35760
rect 29052 35748 29058 35760
rect 32048 35748 32076 35992
rect 32320 35748 33120 35762
rect 29052 35720 29960 35748
rect 32048 35720 33120 35748
rect 29052 35708 29058 35720
rect 23385 35683 23443 35689
rect 19260 35652 19380 35680
rect 18509 35643 18567 35649
rect 17310 35612 17316 35624
rect 16960 35584 17316 35612
rect 17310 35572 17316 35584
rect 17368 35612 17374 35624
rect 17405 35615 17463 35621
rect 17405 35612 17417 35615
rect 17368 35584 17417 35612
rect 17368 35572 17374 35584
rect 17405 35581 17417 35584
rect 17451 35581 17463 35615
rect 18046 35612 18052 35624
rect 18007 35584 18052 35612
rect 17405 35575 17463 35581
rect 18046 35572 18052 35584
rect 18104 35572 18110 35624
rect 19242 35612 19248 35624
rect 19203 35584 19248 35612
rect 19242 35572 19248 35584
rect 19300 35572 19306 35624
rect 19352 35612 19380 35652
rect 23385 35649 23397 35683
rect 23431 35649 23443 35683
rect 23842 35680 23848 35692
rect 23803 35652 23848 35680
rect 23385 35643 23443 35649
rect 23842 35640 23848 35652
rect 23900 35640 23906 35692
rect 25041 35683 25099 35689
rect 25041 35649 25053 35683
rect 25087 35680 25099 35683
rect 27724 35680 27752 35708
rect 27982 35680 27988 35692
rect 25087 35652 27752 35680
rect 27943 35652 27988 35680
rect 25087 35649 25099 35652
rect 25041 35643 25099 35649
rect 19352 35584 20760 35612
rect 15378 35504 15384 35556
rect 15436 35544 15442 35556
rect 15942 35547 16000 35553
rect 15942 35544 15954 35547
rect 15436 35516 15954 35544
rect 15436 35504 15442 35516
rect 15942 35513 15954 35516
rect 15988 35513 16000 35547
rect 18966 35544 18972 35556
rect 15942 35507 16000 35513
rect 16040 35516 18972 35544
rect 16040 35476 16068 35516
rect 18966 35504 18972 35516
rect 19024 35504 19030 35556
rect 19518 35553 19524 35556
rect 19512 35507 19524 35553
rect 19576 35544 19582 35556
rect 19576 35516 19612 35544
rect 19518 35504 19524 35507
rect 19576 35504 19582 35516
rect 16942 35476 16948 35488
rect 15028 35448 16068 35476
rect 16903 35448 16948 35476
rect 14829 35439 14887 35445
rect 16942 35436 16948 35448
rect 17000 35436 17006 35488
rect 17218 35436 17224 35488
rect 17276 35476 17282 35488
rect 17782 35479 17840 35485
rect 17782 35476 17794 35479
rect 17276 35448 17794 35476
rect 17276 35436 17282 35448
rect 17782 35445 17794 35448
rect 17828 35445 17840 35479
rect 17782 35439 17840 35445
rect 19794 35436 19800 35488
rect 19852 35476 19858 35488
rect 20625 35479 20683 35485
rect 20625 35476 20637 35479
rect 19852 35448 20637 35476
rect 19852 35436 19858 35448
rect 20625 35445 20637 35448
rect 20671 35445 20683 35479
rect 20732 35476 20760 35584
rect 21174 35572 21180 35624
rect 21232 35612 21238 35624
rect 21269 35615 21327 35621
rect 21269 35612 21281 35615
rect 21232 35584 21281 35612
rect 21232 35572 21238 35584
rect 21269 35581 21281 35584
rect 21315 35581 21327 35615
rect 21450 35612 21456 35624
rect 21411 35584 21456 35612
rect 21269 35575 21327 35581
rect 21450 35572 21456 35584
rect 21508 35572 21514 35624
rect 22186 35612 22192 35624
rect 22147 35584 22192 35612
rect 22186 35572 22192 35584
rect 22244 35572 22250 35624
rect 23658 35612 23664 35624
rect 23619 35584 23664 35612
rect 23658 35572 23664 35584
rect 23716 35572 23722 35624
rect 24857 35615 24915 35621
rect 24857 35581 24869 35615
rect 24903 35612 24915 35615
rect 25130 35612 25136 35624
rect 24903 35584 25136 35612
rect 24903 35581 24915 35584
rect 24857 35575 24915 35581
rect 25130 35572 25136 35584
rect 25188 35572 25194 35624
rect 25700 35621 25728 35652
rect 27982 35640 27988 35652
rect 28040 35640 28046 35692
rect 28810 35640 28816 35692
rect 28868 35680 28874 35692
rect 29932 35689 29960 35720
rect 32320 35706 33120 35720
rect 29917 35683 29975 35689
rect 28868 35652 29592 35680
rect 28868 35640 28874 35652
rect 25685 35615 25743 35621
rect 25685 35581 25697 35615
rect 25731 35581 25743 35615
rect 25685 35575 25743 35581
rect 27065 35615 27123 35621
rect 27065 35581 27077 35615
rect 27111 35612 27123 35615
rect 27246 35612 27252 35624
rect 27111 35584 27252 35612
rect 27111 35581 27123 35584
rect 27065 35575 27123 35581
rect 27246 35572 27252 35584
rect 27304 35572 27310 35624
rect 27706 35612 27712 35624
rect 27667 35584 27712 35612
rect 27706 35572 27712 35584
rect 27764 35572 27770 35624
rect 27798 35572 27804 35624
rect 27856 35612 27862 35624
rect 27893 35615 27951 35621
rect 27893 35612 27905 35615
rect 27856 35584 27905 35612
rect 27856 35572 27862 35584
rect 27893 35581 27905 35584
rect 27939 35581 27951 35615
rect 27893 35575 27951 35581
rect 28077 35615 28135 35621
rect 28077 35581 28089 35615
rect 28123 35581 28135 35615
rect 28258 35612 28264 35624
rect 28219 35584 28264 35612
rect 28077 35575 28135 35581
rect 20990 35504 20996 35556
rect 21048 35544 21054 35556
rect 21542 35544 21548 35556
rect 21048 35516 21548 35544
rect 21048 35504 21054 35516
rect 21542 35504 21548 35516
rect 21600 35504 21606 35556
rect 22830 35544 22836 35556
rect 22791 35516 22836 35544
rect 22830 35504 22836 35516
rect 22888 35504 22894 35556
rect 23842 35504 23848 35556
rect 23900 35544 23906 35556
rect 25314 35544 25320 35556
rect 23900 35516 25320 35544
rect 23900 35504 23906 35516
rect 25314 35504 25320 35516
rect 25372 35504 25378 35556
rect 26602 35504 26608 35556
rect 26660 35544 26666 35556
rect 26881 35547 26939 35553
rect 26881 35544 26893 35547
rect 26660 35516 26893 35544
rect 26660 35504 26666 35516
rect 26881 35513 26893 35516
rect 26927 35513 26939 35547
rect 26881 35507 26939 35513
rect 27522 35504 27528 35556
rect 27580 35544 27586 35556
rect 28092 35544 28120 35575
rect 28258 35572 28264 35584
rect 28316 35572 28322 35624
rect 29564 35621 29592 35652
rect 29917 35649 29929 35683
rect 29963 35649 29975 35683
rect 29917 35643 29975 35649
rect 28905 35615 28963 35621
rect 28905 35581 28917 35615
rect 28951 35581 28963 35615
rect 28905 35575 28963 35581
rect 29549 35615 29607 35621
rect 29549 35581 29561 35615
rect 29595 35581 29607 35615
rect 29549 35575 29607 35581
rect 27580 35516 28120 35544
rect 28920 35544 28948 35575
rect 29638 35572 29644 35624
rect 29696 35612 29702 35624
rect 29733 35615 29791 35621
rect 29733 35612 29745 35615
rect 29696 35584 29745 35612
rect 29696 35572 29702 35584
rect 29733 35581 29745 35584
rect 29779 35581 29791 35615
rect 29733 35575 29791 35581
rect 29822 35572 29828 35624
rect 29880 35612 29886 35624
rect 30098 35612 30104 35624
rect 29880 35584 29925 35612
rect 30059 35584 30104 35612
rect 29880 35572 29886 35584
rect 30098 35572 30104 35584
rect 30156 35572 30162 35624
rect 29656 35544 29684 35572
rect 30374 35544 30380 35556
rect 28920 35516 29684 35544
rect 30116 35516 30380 35544
rect 27580 35504 27586 35516
rect 22186 35476 22192 35488
rect 20732 35448 22192 35476
rect 20625 35439 20683 35445
rect 22186 35436 22192 35448
rect 22244 35436 22250 35488
rect 22370 35476 22376 35488
rect 22331 35448 22376 35476
rect 22370 35436 22376 35448
rect 22428 35436 22434 35488
rect 25222 35436 25228 35488
rect 25280 35476 25286 35488
rect 25593 35479 25651 35485
rect 25593 35476 25605 35479
rect 25280 35448 25605 35476
rect 25280 35436 25286 35448
rect 25593 35445 25605 35448
rect 25639 35445 25651 35479
rect 25593 35439 25651 35445
rect 27154 35436 27160 35488
rect 27212 35476 27218 35488
rect 30116 35476 30144 35516
rect 30374 35504 30380 35516
rect 30432 35504 30438 35556
rect 30282 35476 30288 35488
rect 27212 35448 30144 35476
rect 30243 35448 30288 35476
rect 27212 35436 27218 35448
rect 30282 35436 30288 35448
rect 30340 35436 30346 35488
rect 30558 35436 30564 35488
rect 30616 35476 30622 35488
rect 30745 35479 30803 35485
rect 30745 35476 30757 35479
rect 30616 35448 30757 35476
rect 30616 35436 30622 35448
rect 30745 35445 30757 35448
rect 30791 35445 30803 35479
rect 30745 35439 30803 35445
rect 1104 35386 32016 35408
rect 1104 35334 11253 35386
rect 11305 35334 11317 35386
rect 11369 35334 11381 35386
rect 11433 35334 11445 35386
rect 11497 35334 11509 35386
rect 11561 35334 21557 35386
rect 21609 35334 21621 35386
rect 21673 35334 21685 35386
rect 21737 35334 21749 35386
rect 21801 35334 21813 35386
rect 21865 35334 32016 35386
rect 1104 35312 32016 35334
rect 2041 35275 2099 35281
rect 2041 35241 2053 35275
rect 2087 35272 2099 35275
rect 2222 35272 2228 35284
rect 2087 35244 2228 35272
rect 2087 35241 2099 35244
rect 2041 35235 2099 35241
rect 2222 35232 2228 35244
rect 2280 35272 2286 35284
rect 5810 35272 5816 35284
rect 2280 35244 5816 35272
rect 2280 35232 2286 35244
rect 5810 35232 5816 35244
rect 5868 35272 5874 35284
rect 9493 35275 9551 35281
rect 5868 35244 8524 35272
rect 5868 35232 5874 35244
rect 8496 35216 8524 35244
rect 9493 35241 9505 35275
rect 9539 35272 9551 35275
rect 10226 35272 10232 35284
rect 9539 35244 10232 35272
rect 9539 35241 9551 35244
rect 9493 35235 9551 35241
rect 10226 35232 10232 35244
rect 10284 35232 10290 35284
rect 12986 35272 12992 35284
rect 10336 35244 12992 35272
rect 2133 35207 2191 35213
rect 2133 35173 2145 35207
rect 2179 35204 2191 35207
rect 3050 35204 3056 35216
rect 2179 35176 3056 35204
rect 2179 35173 2191 35176
rect 2133 35167 2191 35173
rect 3050 35164 3056 35176
rect 3108 35164 3114 35216
rect 3344 35176 7604 35204
rect 3344 35148 3372 35176
rect 2685 35139 2743 35145
rect 2685 35105 2697 35139
rect 2731 35136 2743 35139
rect 2774 35136 2780 35148
rect 2731 35108 2780 35136
rect 2731 35105 2743 35108
rect 2685 35099 2743 35105
rect 2774 35096 2780 35108
rect 2832 35096 2838 35148
rect 3326 35136 3332 35148
rect 3287 35108 3332 35136
rect 3326 35096 3332 35108
rect 3384 35096 3390 35148
rect 3602 35145 3608 35148
rect 3596 35136 3608 35145
rect 3563 35108 3608 35136
rect 3596 35099 3608 35108
rect 3602 35096 3608 35099
rect 3660 35096 3666 35148
rect 5258 35096 5264 35148
rect 5316 35136 5322 35148
rect 5353 35139 5411 35145
rect 5353 35136 5365 35139
rect 5316 35108 5365 35136
rect 5316 35096 5322 35108
rect 5353 35105 5365 35108
rect 5399 35105 5411 35139
rect 5353 35099 5411 35105
rect 5718 35096 5724 35148
rect 5776 35136 5782 35148
rect 6365 35139 6423 35145
rect 6365 35136 6377 35139
rect 5776 35108 6377 35136
rect 5776 35096 5782 35108
rect 6365 35105 6377 35108
rect 6411 35105 6423 35139
rect 6365 35099 6423 35105
rect 7006 35096 7012 35148
rect 7064 35136 7070 35148
rect 7101 35139 7159 35145
rect 7101 35136 7113 35139
rect 7064 35108 7113 35136
rect 7064 35096 7070 35108
rect 7101 35105 7113 35108
rect 7147 35136 7159 35139
rect 7466 35136 7472 35148
rect 7147 35108 7472 35136
rect 7147 35105 7159 35108
rect 7101 35099 7159 35105
rect 7466 35096 7472 35108
rect 7524 35096 7530 35148
rect 7576 35145 7604 35176
rect 8478 35164 8484 35216
rect 8536 35164 8542 35216
rect 9398 35164 9404 35216
rect 9456 35204 9462 35216
rect 10336 35204 10364 35244
rect 12986 35232 12992 35244
rect 13044 35232 13050 35284
rect 13817 35275 13875 35281
rect 13817 35272 13829 35275
rect 13280 35244 13829 35272
rect 9456 35176 10364 35204
rect 9456 35164 9462 35176
rect 10410 35164 10416 35216
rect 10468 35204 10474 35216
rect 10606 35207 10664 35213
rect 10606 35204 10618 35207
rect 10468 35176 10618 35204
rect 10468 35164 10474 35176
rect 10606 35173 10618 35176
rect 10652 35173 10664 35207
rect 10606 35167 10664 35173
rect 11698 35164 11704 35216
rect 11756 35204 11762 35216
rect 12066 35204 12072 35216
rect 11756 35176 12072 35204
rect 11756 35164 11762 35176
rect 12066 35164 12072 35176
rect 12124 35164 12130 35216
rect 13112 35207 13170 35213
rect 13112 35173 13124 35207
rect 13158 35204 13170 35207
rect 13280 35204 13308 35244
rect 13817 35241 13829 35244
rect 13863 35241 13875 35275
rect 13817 35235 13875 35241
rect 14734 35232 14740 35284
rect 14792 35272 14798 35284
rect 15286 35272 15292 35284
rect 14792 35244 15292 35272
rect 14792 35232 14798 35244
rect 13158 35176 13308 35204
rect 13372 35176 14412 35204
rect 13158 35173 13170 35176
rect 13112 35167 13170 35173
rect 7834 35145 7840 35148
rect 7561 35139 7619 35145
rect 7561 35105 7573 35139
rect 7607 35105 7619 35139
rect 7561 35099 7619 35105
rect 7828 35099 7840 35145
rect 7892 35136 7898 35148
rect 8496 35136 8524 35164
rect 10226 35136 10232 35148
rect 7892 35108 7928 35136
rect 8496 35108 10232 35136
rect 7834 35096 7840 35099
rect 7892 35096 7898 35108
rect 10226 35096 10232 35108
rect 10284 35096 10290 35148
rect 10873 35139 10931 35145
rect 10873 35105 10885 35139
rect 10919 35136 10931 35139
rect 11054 35136 11060 35148
rect 10919 35108 11060 35136
rect 10919 35105 10931 35108
rect 10873 35099 10931 35105
rect 11054 35096 11060 35108
rect 11112 35096 11118 35148
rect 12158 35096 12164 35148
rect 12216 35136 12222 35148
rect 13372 35145 13400 35176
rect 13357 35139 13415 35145
rect 12216 35108 13308 35136
rect 12216 35096 12222 35108
rect 2038 35028 2044 35080
rect 2096 35068 2102 35080
rect 2866 35068 2872 35080
rect 2096 35040 2872 35068
rect 2096 35028 2102 35040
rect 2866 35028 2872 35040
rect 2924 35028 2930 35080
rect 4706 35000 4712 35012
rect 4619 34972 4712 35000
rect 4706 34960 4712 34972
rect 4764 35000 4770 35012
rect 5276 35000 5304 35096
rect 13280 35068 13308 35108
rect 13357 35105 13369 35139
rect 13403 35105 13415 35139
rect 13357 35099 13415 35105
rect 14001 35139 14059 35145
rect 14001 35105 14013 35139
rect 14047 35105 14059 35139
rect 14001 35099 14059 35105
rect 14016 35068 14044 35099
rect 13280 35040 14044 35068
rect 14384 35068 14412 35176
rect 14458 35096 14464 35148
rect 14516 35136 14522 35148
rect 14737 35139 14795 35145
rect 14737 35136 14749 35139
rect 14516 35108 14749 35136
rect 14516 35096 14522 35108
rect 14737 35105 14749 35108
rect 14783 35105 14795 35139
rect 14918 35136 14924 35148
rect 14879 35108 14924 35136
rect 14737 35099 14795 35105
rect 14918 35096 14924 35108
rect 14976 35096 14982 35148
rect 15120 35145 15148 35244
rect 15286 35232 15292 35244
rect 15344 35232 15350 35284
rect 15470 35272 15476 35284
rect 15431 35244 15476 35272
rect 15470 35232 15476 35244
rect 15528 35232 15534 35284
rect 17126 35272 17132 35284
rect 16868 35244 17132 35272
rect 16868 35216 16896 35244
rect 17126 35232 17132 35244
rect 17184 35272 17190 35284
rect 22462 35272 22468 35284
rect 17184 35244 22468 35272
rect 17184 35232 17190 35244
rect 22462 35232 22468 35244
rect 22520 35232 22526 35284
rect 23566 35232 23572 35284
rect 23624 35272 23630 35284
rect 23845 35275 23903 35281
rect 23845 35272 23857 35275
rect 23624 35244 23857 35272
rect 23624 35232 23630 35244
rect 23845 35241 23857 35244
rect 23891 35241 23903 35275
rect 24854 35272 24860 35284
rect 24815 35244 24860 35272
rect 23845 35235 23903 35241
rect 24854 35232 24860 35244
rect 24912 35272 24918 35284
rect 25406 35272 25412 35284
rect 24912 35244 25412 35272
rect 24912 35232 24918 35244
rect 25406 35232 25412 35244
rect 25464 35232 25470 35284
rect 26973 35275 27031 35281
rect 26973 35241 26985 35275
rect 27019 35272 27031 35275
rect 27062 35272 27068 35284
rect 27019 35244 27068 35272
rect 27019 35241 27031 35244
rect 26973 35235 27031 35241
rect 27062 35232 27068 35244
rect 27120 35232 27126 35284
rect 28534 35232 28540 35284
rect 28592 35272 28598 35284
rect 29730 35272 29736 35284
rect 28592 35244 29736 35272
rect 28592 35232 28598 35244
rect 29730 35232 29736 35244
rect 29788 35232 29794 35284
rect 16850 35204 16856 35216
rect 15212 35176 16856 35204
rect 15105 35139 15163 35145
rect 15105 35105 15117 35139
rect 15151 35105 15163 35139
rect 15105 35099 15163 35105
rect 14384 35040 14596 35068
rect 4764 34972 5304 35000
rect 14568 35000 14596 35040
rect 14642 35028 14648 35080
rect 14700 35068 14706 35080
rect 15013 35071 15071 35077
rect 15013 35068 15025 35071
rect 14700 35040 15025 35068
rect 14700 35028 14706 35040
rect 15013 35037 15025 35040
rect 15059 35037 15071 35071
rect 15013 35031 15071 35037
rect 15212 35000 15240 35176
rect 16684 35145 16712 35176
rect 16850 35164 16856 35176
rect 16908 35164 16914 35216
rect 18693 35207 18751 35213
rect 18693 35204 18705 35207
rect 18064 35176 18705 35204
rect 16942 35145 16948 35148
rect 15289 35139 15347 35145
rect 15289 35105 15301 35139
rect 15335 35105 15347 35139
rect 15289 35099 15347 35105
rect 16669 35139 16727 35145
rect 16669 35105 16681 35139
rect 16715 35105 16727 35139
rect 16936 35136 16948 35145
rect 16903 35108 16948 35136
rect 16669 35099 16727 35105
rect 16936 35099 16948 35108
rect 15315 35068 15343 35099
rect 16942 35096 16948 35099
rect 17000 35096 17006 35148
rect 15470 35068 15476 35080
rect 15315 35040 15476 35068
rect 15470 35028 15476 35040
rect 15528 35028 15534 35080
rect 14568 34972 15240 35000
rect 4764 34960 4770 34972
rect 15286 34960 15292 35012
rect 15344 35000 15350 35012
rect 18064 35009 18092 35176
rect 18693 35173 18705 35176
rect 18739 35173 18751 35207
rect 18693 35167 18751 35173
rect 19334 35164 19340 35216
rect 19392 35204 19398 35216
rect 29546 35204 29552 35216
rect 19392 35176 19932 35204
rect 19392 35164 19398 35176
rect 19058 35136 19064 35148
rect 19019 35108 19064 35136
rect 19058 35096 19064 35108
rect 19116 35096 19122 35148
rect 19613 35139 19671 35145
rect 19613 35105 19625 35139
rect 19659 35105 19671 35139
rect 19794 35136 19800 35148
rect 19755 35108 19800 35136
rect 19613 35099 19671 35105
rect 18690 35028 18696 35080
rect 18748 35068 18754 35080
rect 19628 35068 19656 35099
rect 19794 35096 19800 35108
rect 19852 35096 19858 35148
rect 19904 35145 19932 35176
rect 22296 35176 29552 35204
rect 19889 35139 19947 35145
rect 19889 35105 19901 35139
rect 19935 35105 19947 35139
rect 19889 35099 19947 35105
rect 20165 35139 20223 35145
rect 20165 35105 20177 35139
rect 20211 35136 20223 35139
rect 20622 35136 20628 35148
rect 20211 35108 20628 35136
rect 20211 35105 20223 35108
rect 20165 35099 20223 35105
rect 20622 35096 20628 35108
rect 20680 35136 20686 35148
rect 21085 35139 21143 35145
rect 21085 35136 21097 35139
rect 20680 35108 21097 35136
rect 20680 35096 20686 35108
rect 21085 35105 21097 35108
rect 21131 35105 21143 35139
rect 21085 35099 21143 35105
rect 21818 35096 21824 35148
rect 21876 35136 21882 35148
rect 21913 35139 21971 35145
rect 21913 35136 21925 35139
rect 21876 35108 21925 35136
rect 21876 35096 21882 35108
rect 21913 35105 21925 35108
rect 21959 35105 21971 35139
rect 21913 35099 21971 35105
rect 22002 35096 22008 35148
rect 22060 35136 22066 35148
rect 22060 35108 22105 35136
rect 22060 35096 22066 35108
rect 19702 35068 19708 35080
rect 18748 35040 18828 35068
rect 19628 35040 19708 35068
rect 18748 35028 18754 35040
rect 15933 35003 15991 35009
rect 15933 35000 15945 35003
rect 15344 34972 15945 35000
rect 15344 34960 15350 34972
rect 15933 34969 15945 34972
rect 15979 34969 15991 35003
rect 15933 34963 15991 34969
rect 18049 35003 18107 35009
rect 18049 34969 18061 35003
rect 18095 34969 18107 35003
rect 18800 35000 18828 35040
rect 19702 35028 19708 35040
rect 19760 35028 19766 35080
rect 19978 35068 19984 35080
rect 19939 35040 19984 35068
rect 19978 35028 19984 35040
rect 20036 35028 20042 35080
rect 22296 35068 22324 35176
rect 29546 35164 29552 35176
rect 29604 35164 29610 35216
rect 22370 35096 22376 35148
rect 22428 35136 22434 35148
rect 22721 35139 22779 35145
rect 22721 35136 22733 35139
rect 22428 35108 22733 35136
rect 22428 35096 22434 35108
rect 22721 35105 22733 35108
rect 22767 35105 22779 35139
rect 22721 35099 22779 35105
rect 25590 35096 25596 35148
rect 25648 35136 25654 35148
rect 25970 35139 26028 35145
rect 25970 35136 25982 35139
rect 25648 35108 25982 35136
rect 25648 35096 25654 35108
rect 25970 35105 25982 35108
rect 26016 35105 26028 35139
rect 25970 35099 26028 35105
rect 27341 35139 27399 35145
rect 27341 35105 27353 35139
rect 27387 35136 27399 35139
rect 27430 35136 27436 35148
rect 27387 35108 27436 35136
rect 27387 35105 27399 35108
rect 27341 35099 27399 35105
rect 27430 35096 27436 35108
rect 27488 35096 27494 35148
rect 27890 35096 27896 35148
rect 27948 35136 27954 35148
rect 27985 35139 28043 35145
rect 27985 35136 27997 35139
rect 27948 35108 27997 35136
rect 27948 35096 27954 35108
rect 27985 35105 27997 35108
rect 28031 35105 28043 35139
rect 27985 35099 28043 35105
rect 29730 35096 29736 35148
rect 29788 35136 29794 35148
rect 30662 35139 30720 35145
rect 30662 35136 30674 35139
rect 29788 35108 30674 35136
rect 29788 35096 29794 35108
rect 30662 35105 30674 35108
rect 30708 35105 30720 35139
rect 30662 35099 30720 35105
rect 22462 35068 22468 35080
rect 20180 35040 22324 35068
rect 22423 35040 22468 35068
rect 20180 35000 20208 35040
rect 22462 35028 22468 35040
rect 22520 35028 22526 35080
rect 26234 35068 26240 35080
rect 26195 35040 26240 35068
rect 26234 35028 26240 35040
rect 26292 35028 26298 35080
rect 27249 35071 27307 35077
rect 27249 35068 27261 35071
rect 26344 35040 27261 35068
rect 21177 35003 21235 35009
rect 18049 34963 18107 34969
rect 18340 34972 18736 35000
rect 18800 34972 20208 35000
rect 20272 34972 20576 35000
rect 2777 34935 2835 34941
rect 2777 34901 2789 34935
rect 2823 34932 2835 34935
rect 2866 34932 2872 34944
rect 2823 34904 2872 34932
rect 2823 34901 2835 34904
rect 2777 34895 2835 34901
rect 2866 34892 2872 34904
rect 2924 34892 2930 34944
rect 3510 34892 3516 34944
rect 3568 34932 3574 34944
rect 3694 34932 3700 34944
rect 3568 34904 3700 34932
rect 3568 34892 3574 34904
rect 3694 34892 3700 34904
rect 3752 34892 3758 34944
rect 5261 34935 5319 34941
rect 5261 34901 5273 34935
rect 5307 34932 5319 34935
rect 5350 34932 5356 34944
rect 5307 34904 5356 34932
rect 5307 34901 5319 34904
rect 5261 34895 5319 34901
rect 5350 34892 5356 34904
rect 5408 34892 5414 34944
rect 5810 34892 5816 34944
rect 5868 34932 5874 34944
rect 6457 34935 6515 34941
rect 6457 34932 6469 34935
rect 5868 34904 6469 34932
rect 5868 34892 5874 34904
rect 6457 34901 6469 34904
rect 6503 34901 6515 34935
rect 8938 34932 8944 34944
rect 8899 34904 8944 34932
rect 6457 34895 6515 34901
rect 8938 34892 8944 34904
rect 8996 34892 9002 34944
rect 9214 34892 9220 34944
rect 9272 34932 9278 34944
rect 10686 34932 10692 34944
rect 9272 34904 10692 34932
rect 9272 34892 9278 34904
rect 10686 34892 10692 34904
rect 10744 34892 10750 34944
rect 11977 34935 12035 34941
rect 11977 34901 11989 34935
rect 12023 34932 12035 34935
rect 13354 34932 13360 34944
rect 12023 34904 13360 34932
rect 12023 34901 12035 34904
rect 11977 34895 12035 34901
rect 13354 34892 13360 34904
rect 13412 34892 13418 34944
rect 14642 34892 14648 34944
rect 14700 34932 14706 34944
rect 15562 34932 15568 34944
rect 14700 34904 15568 34932
rect 14700 34892 14706 34904
rect 15562 34892 15568 34904
rect 15620 34892 15626 34944
rect 15948 34932 15976 34963
rect 17034 34932 17040 34944
rect 15948 34904 17040 34932
rect 17034 34892 17040 34904
rect 17092 34892 17098 34944
rect 17310 34892 17316 34944
rect 17368 34932 17374 34944
rect 18340 34932 18368 34972
rect 18506 34932 18512 34944
rect 17368 34904 18368 34932
rect 18467 34904 18512 34932
rect 17368 34892 17374 34904
rect 18506 34892 18512 34904
rect 18564 34892 18570 34944
rect 18708 34941 18736 34972
rect 18693 34935 18751 34941
rect 18693 34901 18705 34935
rect 18739 34901 18751 34935
rect 18693 34895 18751 34901
rect 18782 34892 18788 34944
rect 18840 34932 18846 34944
rect 20272 34932 20300 34972
rect 18840 34904 20300 34932
rect 20349 34935 20407 34941
rect 18840 34892 18846 34904
rect 20349 34901 20361 34935
rect 20395 34932 20407 34935
rect 20438 34932 20444 34944
rect 20395 34904 20444 34932
rect 20395 34901 20407 34904
rect 20349 34895 20407 34901
rect 20438 34892 20444 34904
rect 20496 34892 20502 34944
rect 20548 34932 20576 34972
rect 21177 34969 21189 35003
rect 21223 35000 21235 35003
rect 22370 35000 22376 35012
rect 21223 34972 22376 35000
rect 21223 34969 21235 34972
rect 21177 34963 21235 34969
rect 22370 34960 22376 34972
rect 22428 34960 22434 35012
rect 23934 34932 23940 34944
rect 20548 34904 23940 34932
rect 23934 34892 23940 34904
rect 23992 34932 23998 34944
rect 24305 34935 24363 34941
rect 24305 34932 24317 34935
rect 23992 34904 24317 34932
rect 23992 34892 23998 34904
rect 24305 34901 24317 34904
rect 24351 34901 24363 34935
rect 24305 34895 24363 34901
rect 24946 34892 24952 34944
rect 25004 34932 25010 34944
rect 26050 34932 26056 34944
rect 25004 34904 26056 34932
rect 25004 34892 25010 34904
rect 26050 34892 26056 34904
rect 26108 34932 26114 34944
rect 26344 34932 26372 35040
rect 27249 35037 27261 35040
rect 27295 35037 27307 35071
rect 27249 35031 27307 35037
rect 28261 35071 28319 35077
rect 28261 35037 28273 35071
rect 28307 35068 28319 35071
rect 29270 35068 29276 35080
rect 28307 35040 29276 35068
rect 28307 35037 28319 35040
rect 28261 35031 28319 35037
rect 29270 35028 29276 35040
rect 29328 35068 29334 35080
rect 29822 35068 29828 35080
rect 29328 35040 29828 35068
rect 29328 35028 29334 35040
rect 29822 35028 29828 35040
rect 29880 35028 29886 35080
rect 30926 35068 30932 35080
rect 30887 35040 30932 35068
rect 30926 35028 30932 35040
rect 30984 35028 30990 35080
rect 27246 34932 27252 34944
rect 26108 34904 26372 34932
rect 27207 34904 27252 34932
rect 26108 34892 26114 34904
rect 27246 34892 27252 34904
rect 27304 34892 27310 34944
rect 29546 34932 29552 34944
rect 29507 34904 29552 34932
rect 29546 34892 29552 34904
rect 29604 34892 29610 34944
rect 1104 34842 32016 34864
rect 1104 34790 6102 34842
rect 6154 34790 6166 34842
rect 6218 34790 6230 34842
rect 6282 34790 6294 34842
rect 6346 34790 6358 34842
rect 6410 34790 16405 34842
rect 16457 34790 16469 34842
rect 16521 34790 16533 34842
rect 16585 34790 16597 34842
rect 16649 34790 16661 34842
rect 16713 34790 26709 34842
rect 26761 34790 26773 34842
rect 26825 34790 26837 34842
rect 26889 34790 26901 34842
rect 26953 34790 26965 34842
rect 27017 34790 32016 34842
rect 1104 34768 32016 34790
rect 6488 34700 7604 34728
rect 2406 34620 2412 34672
rect 2464 34660 2470 34672
rect 2961 34663 3019 34669
rect 2961 34660 2973 34663
rect 2464 34632 2973 34660
rect 2464 34620 2470 34632
rect 2961 34629 2973 34632
rect 3007 34660 3019 34663
rect 3234 34660 3240 34672
rect 3007 34632 3240 34660
rect 3007 34629 3019 34632
rect 2961 34623 3019 34629
rect 3234 34620 3240 34632
rect 3292 34620 3298 34672
rect 5445 34663 5503 34669
rect 5445 34629 5457 34663
rect 5491 34660 5503 34663
rect 5491 34632 6408 34660
rect 5491 34629 5503 34632
rect 5445 34623 5503 34629
rect 6380 34536 6408 34632
rect 1581 34527 1639 34533
rect 1581 34493 1593 34527
rect 1627 34524 1639 34527
rect 1670 34524 1676 34536
rect 1627 34496 1676 34524
rect 1627 34493 1639 34496
rect 1581 34487 1639 34493
rect 1670 34484 1676 34496
rect 1728 34484 1734 34536
rect 2038 34524 2044 34536
rect 1999 34496 2044 34524
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2222 34524 2228 34536
rect 2183 34496 2228 34524
rect 2222 34484 2228 34496
rect 2280 34484 2286 34536
rect 4246 34484 4252 34536
rect 4304 34524 4310 34536
rect 4525 34527 4583 34533
rect 4525 34524 4537 34527
rect 4304 34496 4537 34524
rect 4304 34484 4310 34496
rect 4525 34493 4537 34496
rect 4571 34493 4583 34527
rect 4525 34487 4583 34493
rect 4706 34484 4712 34536
rect 4764 34524 4770 34536
rect 4801 34527 4859 34533
rect 4801 34524 4813 34527
rect 4764 34496 4813 34524
rect 4764 34484 4770 34496
rect 4801 34493 4813 34496
rect 4847 34493 4859 34527
rect 5258 34524 5264 34536
rect 5219 34496 5264 34524
rect 4801 34487 4859 34493
rect 5258 34484 5264 34496
rect 5316 34484 5322 34536
rect 5445 34527 5503 34533
rect 5445 34493 5457 34527
rect 5491 34524 5503 34527
rect 5718 34524 5724 34536
rect 5491 34496 5724 34524
rect 5491 34493 5503 34496
rect 5445 34487 5503 34493
rect 2774 34416 2780 34468
rect 2832 34456 2838 34468
rect 2832 34428 2877 34456
rect 2832 34416 2838 34428
rect 5166 34416 5172 34468
rect 5224 34456 5230 34468
rect 5460 34456 5488 34487
rect 5718 34484 5724 34496
rect 5776 34484 5782 34536
rect 6362 34484 6368 34536
rect 6420 34484 6426 34536
rect 6488 34533 6516 34700
rect 7374 34620 7380 34672
rect 7432 34620 7438 34672
rect 7576 34660 7604 34700
rect 7834 34688 7840 34740
rect 7892 34728 7898 34740
rect 7929 34731 7987 34737
rect 7929 34728 7941 34731
rect 7892 34700 7941 34728
rect 7892 34688 7898 34700
rect 7929 34697 7941 34700
rect 7975 34697 7987 34731
rect 7929 34691 7987 34697
rect 10134 34688 10140 34740
rect 10192 34728 10198 34740
rect 10321 34731 10379 34737
rect 10321 34728 10333 34731
rect 10192 34700 10333 34728
rect 10192 34688 10198 34700
rect 10321 34697 10333 34700
rect 10367 34697 10379 34731
rect 10321 34691 10379 34697
rect 10686 34688 10692 34740
rect 10744 34728 10750 34740
rect 11701 34731 11759 34737
rect 11701 34728 11713 34731
rect 10744 34700 11713 34728
rect 10744 34688 10750 34700
rect 11701 34697 11713 34700
rect 11747 34697 11759 34731
rect 11701 34691 11759 34697
rect 13357 34731 13415 34737
rect 13357 34697 13369 34731
rect 13403 34697 13415 34731
rect 13538 34728 13544 34740
rect 13499 34700 13544 34728
rect 13357 34691 13415 34697
rect 7650 34660 7656 34672
rect 7576 34632 7656 34660
rect 7650 34620 7656 34632
rect 7708 34660 7714 34672
rect 7708 34632 8064 34660
rect 7708 34620 7714 34632
rect 6733 34595 6791 34601
rect 6733 34561 6745 34595
rect 6779 34561 6791 34595
rect 7392 34592 7420 34620
rect 7469 34595 7527 34601
rect 7469 34592 7481 34595
rect 7392 34564 7481 34592
rect 6733 34555 6791 34561
rect 7469 34561 7481 34564
rect 7515 34561 7527 34595
rect 7926 34592 7932 34604
rect 7469 34555 7527 34561
rect 7668 34564 7932 34592
rect 6457 34527 6516 34533
rect 6457 34493 6469 34527
rect 6503 34496 6516 34527
rect 6549 34527 6607 34533
rect 6503 34493 6515 34496
rect 6457 34487 6515 34493
rect 6549 34493 6561 34527
rect 6595 34493 6607 34527
rect 6549 34487 6607 34493
rect 5224 34428 5488 34456
rect 5224 34416 5230 34428
rect 6564 34400 6592 34487
rect 6748 34456 6776 34555
rect 7006 34484 7012 34536
rect 7064 34524 7070 34536
rect 7193 34527 7251 34533
rect 7193 34524 7205 34527
rect 7064 34496 7205 34524
rect 7064 34484 7070 34496
rect 7193 34493 7205 34496
rect 7239 34493 7251 34527
rect 7374 34524 7380 34536
rect 7335 34496 7380 34524
rect 7193 34487 7251 34493
rect 7374 34484 7380 34496
rect 7432 34484 7438 34536
rect 7561 34527 7619 34533
rect 7561 34493 7573 34527
rect 7607 34526 7619 34527
rect 7668 34526 7696 34564
rect 7926 34552 7932 34564
rect 7984 34552 7990 34604
rect 7607 34498 7696 34526
rect 7745 34527 7803 34533
rect 7607 34493 7619 34498
rect 7561 34487 7619 34493
rect 7745 34493 7757 34527
rect 7791 34524 7803 34527
rect 8036 34524 8064 34632
rect 9674 34620 9680 34672
rect 9732 34660 9738 34672
rect 11057 34663 11115 34669
rect 11057 34660 11069 34663
rect 9732 34632 11069 34660
rect 9732 34620 9738 34632
rect 11057 34629 11069 34632
rect 11103 34629 11115 34663
rect 11057 34623 11115 34629
rect 12618 34620 12624 34672
rect 12676 34660 12682 34672
rect 12989 34663 13047 34669
rect 12989 34660 13001 34663
rect 12676 34632 13001 34660
rect 12676 34620 12682 34632
rect 12989 34629 13001 34632
rect 13035 34629 13047 34663
rect 13372 34660 13400 34691
rect 13538 34688 13544 34700
rect 13596 34688 13602 34740
rect 14366 34688 14372 34740
rect 14424 34728 14430 34740
rect 14737 34731 14795 34737
rect 14737 34728 14749 34731
rect 14424 34700 14749 34728
rect 14424 34688 14430 34700
rect 14737 34697 14749 34700
rect 14783 34697 14795 34731
rect 14737 34691 14795 34697
rect 14921 34731 14979 34737
rect 14921 34697 14933 34731
rect 14967 34728 14979 34731
rect 15010 34728 15016 34740
rect 14967 34700 15016 34728
rect 14967 34697 14979 34700
rect 14921 34691 14979 34697
rect 13722 34660 13728 34672
rect 13372 34632 13728 34660
rect 12989 34623 13047 34629
rect 13722 34620 13728 34632
rect 13780 34620 13786 34672
rect 8938 34592 8944 34604
rect 8851 34564 8944 34592
rect 8938 34552 8944 34564
rect 8996 34592 9002 34604
rect 8996 34564 9674 34592
rect 8996 34552 9002 34564
rect 8110 34524 8116 34536
rect 7791 34496 8116 34524
rect 7791 34493 7803 34496
rect 7745 34487 7803 34493
rect 8110 34484 8116 34496
rect 8168 34524 8174 34536
rect 9217 34527 9275 34533
rect 9217 34524 9229 34527
rect 8168 34496 9229 34524
rect 8168 34484 8174 34496
rect 9217 34493 9229 34496
rect 9263 34524 9275 34527
rect 9306 34524 9312 34536
rect 9263 34496 9312 34524
rect 9263 34493 9275 34496
rect 9217 34487 9275 34493
rect 9306 34484 9312 34496
rect 9364 34484 9370 34536
rect 9646 34524 9674 34564
rect 12158 34552 12164 34604
rect 12216 34592 12222 34604
rect 14642 34592 14648 34604
rect 12216 34564 14648 34592
rect 12216 34552 12222 34564
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 10965 34527 11023 34533
rect 10965 34524 10977 34527
rect 9646 34496 10977 34524
rect 10965 34493 10977 34496
rect 11011 34493 11023 34527
rect 10965 34487 11023 34493
rect 14369 34527 14427 34533
rect 14369 34493 14381 34527
rect 14415 34524 14427 34527
rect 14458 34524 14464 34536
rect 14415 34496 14464 34524
rect 14415 34493 14427 34496
rect 14369 34487 14427 34493
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 14752 34524 14780 34691
rect 15010 34688 15016 34700
rect 15068 34688 15074 34740
rect 15378 34728 15384 34740
rect 15339 34700 15384 34728
rect 15378 34688 15384 34700
rect 15436 34688 15442 34740
rect 17034 34688 17040 34740
rect 17092 34728 17098 34740
rect 17494 34728 17500 34740
rect 17092 34700 17500 34728
rect 17092 34688 17098 34700
rect 17494 34688 17500 34700
rect 17552 34688 17558 34740
rect 26145 34731 26203 34737
rect 18708 34700 25544 34728
rect 15470 34620 15476 34672
rect 15528 34660 15534 34672
rect 15528 34632 15976 34660
rect 15528 34620 15534 34632
rect 15378 34552 15384 34604
rect 15436 34592 15442 34604
rect 15749 34595 15807 34601
rect 15749 34592 15761 34595
rect 15436 34564 15761 34592
rect 15436 34552 15442 34564
rect 15749 34561 15761 34564
rect 15795 34561 15807 34595
rect 15749 34555 15807 34561
rect 15562 34524 15568 34536
rect 14752 34496 15568 34524
rect 15562 34484 15568 34496
rect 15620 34484 15626 34536
rect 15654 34484 15660 34536
rect 15712 34524 15718 34536
rect 15948 34533 15976 34632
rect 16206 34620 16212 34672
rect 16264 34660 16270 34672
rect 16264 34632 18644 34660
rect 16264 34620 16270 34632
rect 16853 34595 16911 34601
rect 16853 34592 16865 34595
rect 16040 34564 16865 34592
rect 15841 34527 15899 34533
rect 15841 34524 15853 34527
rect 15712 34496 15853 34524
rect 15712 34484 15718 34496
rect 15841 34493 15853 34496
rect 15887 34493 15899 34527
rect 15841 34487 15899 34493
rect 15933 34527 15991 34533
rect 15933 34493 15945 34527
rect 15979 34493 15991 34527
rect 15933 34487 15991 34493
rect 7650 34456 7656 34468
rect 6748 34428 7656 34456
rect 7650 34416 7656 34428
rect 7708 34416 7714 34468
rect 10413 34459 10471 34465
rect 10413 34425 10425 34459
rect 10459 34456 10471 34459
rect 10870 34456 10876 34468
rect 10459 34428 10876 34456
rect 10459 34425 10471 34428
rect 10413 34419 10471 34425
rect 10870 34416 10876 34428
rect 10928 34456 10934 34468
rect 11977 34459 12035 34465
rect 10928 34428 11836 34456
rect 10928 34416 10934 34428
rect 2133 34391 2191 34397
rect 2133 34357 2145 34391
rect 2179 34388 2191 34391
rect 2498 34388 2504 34400
rect 2179 34360 2504 34388
rect 2179 34357 2191 34360
rect 2133 34351 2191 34357
rect 2498 34348 2504 34360
rect 2556 34348 2562 34400
rect 5718 34348 5724 34400
rect 5776 34388 5782 34400
rect 5905 34391 5963 34397
rect 5905 34388 5917 34391
rect 5776 34360 5917 34388
rect 5776 34348 5782 34360
rect 5905 34357 5917 34360
rect 5951 34357 5963 34391
rect 5905 34351 5963 34357
rect 6546 34348 6552 34400
rect 6604 34348 6610 34400
rect 6730 34388 6736 34400
rect 6691 34360 6736 34388
rect 6730 34348 6736 34360
rect 6788 34348 6794 34400
rect 6822 34348 6828 34400
rect 6880 34388 6886 34400
rect 9214 34388 9220 34400
rect 6880 34360 9220 34388
rect 6880 34348 6886 34360
rect 9214 34348 9220 34360
rect 9272 34348 9278 34400
rect 11808 34388 11836 34428
rect 11977 34425 11989 34459
rect 12023 34456 12035 34459
rect 12986 34456 12992 34468
rect 12023 34428 12992 34456
rect 12023 34425 12035 34428
rect 11977 34419 12035 34425
rect 12986 34416 12992 34428
rect 13044 34416 13050 34468
rect 13354 34456 13360 34468
rect 13315 34428 13360 34456
rect 13354 34416 13360 34428
rect 13412 34416 13418 34468
rect 13446 34416 13452 34468
rect 13504 34456 13510 34468
rect 14182 34456 14188 34468
rect 13504 34428 14188 34456
rect 13504 34416 13510 34428
rect 14182 34416 14188 34428
rect 14240 34456 14246 34468
rect 16040 34456 16068 34564
rect 16853 34561 16865 34564
rect 16899 34561 16911 34595
rect 16853 34555 16911 34561
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34592 17831 34595
rect 18506 34592 18512 34604
rect 17819 34564 18512 34592
rect 17819 34561 17831 34564
rect 17773 34555 17831 34561
rect 18506 34552 18512 34564
rect 18564 34552 18570 34604
rect 16117 34527 16175 34533
rect 16117 34493 16129 34527
rect 16163 34493 16175 34527
rect 18046 34524 18052 34536
rect 18007 34496 18052 34524
rect 16117 34487 16175 34493
rect 14240 34428 16068 34456
rect 14240 34416 14246 34428
rect 12066 34388 12072 34400
rect 11808 34360 12072 34388
rect 12066 34348 12072 34360
rect 12124 34348 12130 34400
rect 14734 34388 14740 34400
rect 14695 34360 14740 34388
rect 14734 34348 14740 34360
rect 14792 34348 14798 34400
rect 15010 34348 15016 34400
rect 15068 34388 15074 34400
rect 15838 34388 15844 34400
rect 15068 34360 15844 34388
rect 15068 34348 15074 34360
rect 15838 34348 15844 34360
rect 15896 34388 15902 34400
rect 16132 34388 16160 34487
rect 18046 34484 18052 34496
rect 18104 34484 18110 34536
rect 18322 34484 18328 34536
rect 18380 34524 18386 34536
rect 18417 34527 18475 34533
rect 18417 34524 18429 34527
rect 18380 34496 18429 34524
rect 18380 34484 18386 34496
rect 18417 34493 18429 34496
rect 18463 34493 18475 34527
rect 18616 34524 18644 34632
rect 18708 34601 18736 34700
rect 18966 34620 18972 34672
rect 19024 34660 19030 34672
rect 19978 34660 19984 34672
rect 19024 34632 19984 34660
rect 19024 34620 19030 34632
rect 19978 34620 19984 34632
rect 20036 34620 20042 34672
rect 23934 34620 23940 34672
rect 23992 34660 23998 34672
rect 24302 34660 24308 34672
rect 23992 34632 24308 34660
rect 23992 34620 23998 34632
rect 24302 34620 24308 34632
rect 24360 34620 24366 34672
rect 25222 34620 25228 34672
rect 25280 34620 25286 34672
rect 18693 34595 18751 34601
rect 18693 34561 18705 34595
rect 18739 34561 18751 34595
rect 19337 34595 19395 34601
rect 19337 34592 19349 34595
rect 18693 34555 18751 34561
rect 18800 34564 19349 34592
rect 18800 34524 18828 34564
rect 19337 34561 19349 34564
rect 19383 34561 19395 34595
rect 19337 34555 19395 34561
rect 19610 34552 19616 34604
rect 19668 34592 19674 34604
rect 25133 34595 25191 34601
rect 19668 34564 20300 34592
rect 19668 34552 19674 34564
rect 18616 34496 18828 34524
rect 18417 34487 18475 34493
rect 19242 34484 19248 34536
rect 19300 34524 19306 34536
rect 20165 34527 20223 34533
rect 20165 34524 20177 34527
rect 19300 34496 20177 34524
rect 19300 34484 19306 34496
rect 20165 34493 20177 34496
rect 20211 34493 20223 34527
rect 20272 34524 20300 34564
rect 25133 34561 25145 34595
rect 25179 34592 25191 34595
rect 25240 34592 25268 34620
rect 25179 34564 25268 34592
rect 25516 34592 25544 34700
rect 26145 34697 26157 34731
rect 26191 34728 26203 34731
rect 26602 34728 26608 34740
rect 26191 34700 26608 34728
rect 26191 34697 26203 34700
rect 26145 34691 26203 34697
rect 26602 34688 26608 34700
rect 26660 34688 26666 34740
rect 29549 34731 29607 34737
rect 29549 34697 29561 34731
rect 29595 34728 29607 34731
rect 29638 34728 29644 34740
rect 29595 34700 29644 34728
rect 29595 34697 29607 34700
rect 29549 34691 29607 34697
rect 29638 34688 29644 34700
rect 29696 34728 29702 34740
rect 30006 34728 30012 34740
rect 29696 34700 30012 34728
rect 29696 34688 29702 34700
rect 30006 34688 30012 34700
rect 30064 34688 30070 34740
rect 25590 34620 25596 34672
rect 25648 34660 25654 34672
rect 28994 34660 29000 34672
rect 25648 34632 25693 34660
rect 25648 34620 25654 34632
rect 28966 34620 29000 34660
rect 29052 34620 29058 34672
rect 26602 34592 26608 34604
rect 25516 34564 26608 34592
rect 25179 34561 25191 34564
rect 25133 34555 25191 34561
rect 26602 34552 26608 34564
rect 26660 34552 26666 34604
rect 28721 34595 28779 34601
rect 28721 34561 28733 34595
rect 28767 34592 28779 34595
rect 28966 34592 28994 34620
rect 30926 34592 30932 34604
rect 28767 34564 28994 34592
rect 30887 34564 30932 34592
rect 28767 34561 28779 34564
rect 28721 34555 28779 34561
rect 30926 34552 30932 34564
rect 30984 34552 30990 34604
rect 22005 34527 22063 34533
rect 22005 34524 22017 34527
rect 20272 34496 22017 34524
rect 20165 34487 20223 34493
rect 22005 34493 22017 34496
rect 22051 34493 22063 34527
rect 22261 34527 22319 34533
rect 22261 34524 22273 34527
rect 22005 34487 22063 34493
rect 22112 34496 22273 34524
rect 16669 34459 16727 34465
rect 16669 34425 16681 34459
rect 16715 34456 16727 34459
rect 16758 34456 16764 34468
rect 16715 34428 16764 34456
rect 16715 34425 16727 34428
rect 16669 34419 16727 34425
rect 16758 34416 16764 34428
rect 16816 34456 16822 34468
rect 17034 34456 17040 34468
rect 16816 34428 17040 34456
rect 16816 34416 16822 34428
rect 17034 34416 17040 34428
rect 17092 34416 17098 34468
rect 17954 34416 17960 34468
rect 18012 34456 18018 34468
rect 19260 34456 19288 34484
rect 20438 34465 20444 34468
rect 20432 34456 20444 34465
rect 18012 34428 19288 34456
rect 20399 34428 20444 34456
rect 18012 34416 18018 34428
rect 20432 34419 20444 34428
rect 20438 34416 20444 34419
rect 20496 34416 20502 34468
rect 20714 34416 20720 34468
rect 20772 34456 20778 34468
rect 22112 34456 22140 34496
rect 22261 34493 22273 34496
rect 22307 34493 22319 34527
rect 24854 34524 24860 34536
rect 24815 34496 24860 34524
rect 22261 34487 22319 34493
rect 24854 34484 24860 34496
rect 24912 34484 24918 34536
rect 25041 34527 25099 34533
rect 25041 34493 25053 34527
rect 25087 34493 25099 34527
rect 25041 34487 25099 34493
rect 25225 34527 25283 34533
rect 25225 34493 25237 34527
rect 25271 34524 25283 34527
rect 25314 34524 25320 34536
rect 25271 34496 25320 34524
rect 25271 34493 25283 34496
rect 25225 34487 25283 34493
rect 20772 34428 22140 34456
rect 25056 34456 25084 34487
rect 25314 34484 25320 34496
rect 25372 34484 25378 34536
rect 25406 34484 25412 34536
rect 25464 34524 25470 34536
rect 26050 34524 26056 34536
rect 25464 34496 25509 34524
rect 26011 34496 26056 34524
rect 25464 34484 25470 34496
rect 26050 34484 26056 34496
rect 26108 34484 26114 34536
rect 26510 34484 26516 34536
rect 26568 34524 26574 34536
rect 28997 34527 29055 34533
rect 28997 34524 29009 34527
rect 26568 34496 29009 34524
rect 26568 34484 26574 34496
rect 26142 34456 26148 34468
rect 25056 34428 26148 34456
rect 20772 34416 20778 34428
rect 26142 34416 26148 34428
rect 26200 34416 26206 34468
rect 27264 34465 27292 34496
rect 28997 34493 29009 34496
rect 29043 34493 29055 34527
rect 28997 34487 29055 34493
rect 30282 34484 30288 34536
rect 30340 34524 30346 34536
rect 30662 34527 30720 34533
rect 30662 34524 30674 34527
rect 30340 34496 30674 34524
rect 30340 34484 30346 34496
rect 30662 34493 30674 34496
rect 30708 34493 30720 34527
rect 30662 34487 30720 34493
rect 27249 34459 27307 34465
rect 27249 34425 27261 34459
rect 27295 34456 27307 34459
rect 27295 34428 27329 34456
rect 27295 34425 27307 34428
rect 27249 34419 27307 34425
rect 15896 34360 16160 34388
rect 15896 34348 15902 34360
rect 16298 34348 16304 34400
rect 16356 34388 16362 34400
rect 20530 34388 20536 34400
rect 16356 34360 20536 34388
rect 16356 34348 16362 34360
rect 20530 34348 20536 34360
rect 20588 34348 20594 34400
rect 20622 34348 20628 34400
rect 20680 34388 20686 34400
rect 21545 34391 21603 34397
rect 21545 34388 21557 34391
rect 20680 34360 21557 34388
rect 20680 34348 20686 34360
rect 21545 34357 21557 34360
rect 21591 34357 21603 34391
rect 21545 34351 21603 34357
rect 22002 34348 22008 34400
rect 22060 34388 22066 34400
rect 22646 34388 22652 34400
rect 22060 34360 22652 34388
rect 22060 34348 22066 34360
rect 22646 34348 22652 34360
rect 22704 34388 22710 34400
rect 23385 34391 23443 34397
rect 23385 34388 23397 34391
rect 22704 34360 23397 34388
rect 22704 34348 22710 34360
rect 23385 34357 23397 34360
rect 23431 34357 23443 34391
rect 23385 34351 23443 34357
rect 25314 34348 25320 34400
rect 25372 34388 25378 34400
rect 27157 34391 27215 34397
rect 27157 34388 27169 34391
rect 25372 34360 27169 34388
rect 25372 34348 25378 34360
rect 27157 34357 27169 34360
rect 27203 34388 27215 34391
rect 28074 34388 28080 34400
rect 27203 34360 28080 34388
rect 27203 34357 27215 34360
rect 27157 34351 27215 34357
rect 28074 34348 28080 34360
rect 28132 34348 28138 34400
rect 1104 34298 32016 34320
rect 1104 34246 11253 34298
rect 11305 34246 11317 34298
rect 11369 34246 11381 34298
rect 11433 34246 11445 34298
rect 11497 34246 11509 34298
rect 11561 34246 21557 34298
rect 21609 34246 21621 34298
rect 21673 34246 21685 34298
rect 21737 34246 21749 34298
rect 21801 34246 21813 34298
rect 21865 34246 32016 34298
rect 1104 34224 32016 34246
rect 5350 34184 5356 34196
rect 4540 34156 5356 34184
rect 2498 34076 2504 34128
rect 2556 34116 2562 34128
rect 2593 34119 2651 34125
rect 2593 34116 2605 34119
rect 2556 34088 2605 34116
rect 2556 34076 2562 34088
rect 2593 34085 2605 34088
rect 2639 34085 2651 34119
rect 2593 34079 2651 34085
rect 1394 34048 1400 34060
rect 768 34020 1400 34048
rect 768 33844 796 34020
rect 1394 34008 1400 34020
rect 1452 34008 1458 34060
rect 2685 34051 2743 34057
rect 2685 34017 2697 34051
rect 2731 34048 2743 34051
rect 3326 34048 3332 34060
rect 2731 34020 3332 34048
rect 2731 34017 2743 34020
rect 2685 34011 2743 34017
rect 3326 34008 3332 34020
rect 3384 34008 3390 34060
rect 4540 34057 4568 34156
rect 5350 34144 5356 34156
rect 5408 34144 5414 34196
rect 6178 34144 6184 34196
rect 6236 34184 6242 34196
rect 6365 34187 6423 34193
rect 6365 34184 6377 34187
rect 6236 34156 6377 34184
rect 6236 34144 6242 34156
rect 6365 34153 6377 34156
rect 6411 34153 6423 34187
rect 6365 34147 6423 34153
rect 6454 34144 6460 34196
rect 6512 34184 6518 34196
rect 6822 34184 6828 34196
rect 6512 34156 6828 34184
rect 6512 34144 6518 34156
rect 6822 34144 6828 34156
rect 6880 34144 6886 34196
rect 9306 34144 9312 34196
rect 9364 34184 9370 34196
rect 9364 34156 10640 34184
rect 9364 34144 9370 34156
rect 4617 34119 4675 34125
rect 4617 34085 4629 34119
rect 4663 34116 4675 34119
rect 6733 34119 6791 34125
rect 6733 34116 6745 34119
rect 4663 34088 6745 34116
rect 4663 34085 4675 34088
rect 4617 34079 4675 34085
rect 6472 34060 6500 34088
rect 6733 34085 6745 34088
rect 6779 34085 6791 34119
rect 6733 34079 6791 34085
rect 8938 34076 8944 34128
rect 8996 34116 9002 34128
rect 9033 34119 9091 34125
rect 9033 34116 9045 34119
rect 8996 34088 9045 34116
rect 8996 34076 9002 34088
rect 9033 34085 9045 34088
rect 9079 34085 9091 34119
rect 9033 34079 9091 34085
rect 9122 34076 9128 34128
rect 9180 34076 9186 34128
rect 10612 34125 10640 34156
rect 14090 34144 14096 34196
rect 14148 34184 14154 34196
rect 15749 34187 15807 34193
rect 15749 34184 15761 34187
rect 14148 34156 15761 34184
rect 14148 34144 14154 34156
rect 15749 34153 15761 34156
rect 15795 34153 15807 34187
rect 15749 34147 15807 34153
rect 19429 34187 19487 34193
rect 19429 34153 19441 34187
rect 19475 34184 19487 34187
rect 19518 34184 19524 34196
rect 19475 34156 19524 34184
rect 19475 34153 19487 34156
rect 19429 34147 19487 34153
rect 19518 34144 19524 34156
rect 19576 34144 19582 34196
rect 20714 34184 20720 34196
rect 20675 34156 20720 34184
rect 20714 34144 20720 34156
rect 20772 34144 20778 34196
rect 23845 34187 23903 34193
rect 23845 34153 23857 34187
rect 23891 34153 23903 34187
rect 23845 34147 23903 34153
rect 10381 34119 10439 34125
rect 10381 34116 10393 34119
rect 9508 34088 10393 34116
rect 3973 34051 4031 34057
rect 3973 34017 3985 34051
rect 4019 34048 4031 34051
rect 4525 34051 4583 34057
rect 4019 34020 4476 34048
rect 4019 34017 4031 34020
rect 3973 34011 4031 34017
rect 2501 33983 2559 33989
rect 2501 33949 2513 33983
rect 2547 33949 2559 33983
rect 2501 33943 2559 33949
rect 2516 33912 2544 33943
rect 2774 33912 2780 33924
rect 2516 33884 2780 33912
rect 2774 33872 2780 33884
rect 2832 33872 2838 33924
rect 768 33816 888 33844
rect 0 33708 800 33722
rect 860 33708 888 33816
rect 1394 33804 1400 33856
rect 1452 33844 1458 33856
rect 1581 33847 1639 33853
rect 1581 33844 1593 33847
rect 1452 33816 1593 33844
rect 1452 33804 1458 33816
rect 1581 33813 1593 33816
rect 1627 33813 1639 33847
rect 3050 33844 3056 33856
rect 3011 33816 3056 33844
rect 1581 33807 1639 33813
rect 3050 33804 3056 33816
rect 3108 33804 3114 33856
rect 3418 33804 3424 33856
rect 3476 33844 3482 33856
rect 3881 33847 3939 33853
rect 3881 33844 3893 33847
rect 3476 33816 3893 33844
rect 3476 33804 3482 33816
rect 3881 33813 3893 33816
rect 3927 33844 3939 33847
rect 4062 33844 4068 33856
rect 3927 33816 4068 33844
rect 3927 33813 3939 33816
rect 3881 33807 3939 33813
rect 4062 33804 4068 33816
rect 4120 33804 4126 33856
rect 4448 33844 4476 34020
rect 4525 34017 4537 34051
rect 4571 34017 4583 34051
rect 4525 34011 4583 34017
rect 4709 34051 4767 34057
rect 4709 34017 4721 34051
rect 4755 34017 4767 34051
rect 5166 34048 5172 34060
rect 5127 34020 5172 34048
rect 4709 34011 4767 34017
rect 4724 33912 4752 34011
rect 5166 34008 5172 34020
rect 5224 34008 5230 34060
rect 5350 34048 5356 34060
rect 5311 34020 5356 34048
rect 5350 34008 5356 34020
rect 5408 34008 5414 34060
rect 5442 34008 5448 34060
rect 5500 34048 5506 34060
rect 5583 34051 5641 34057
rect 5500 34020 5545 34048
rect 5500 34008 5506 34020
rect 5583 34017 5595 34051
rect 5629 34048 5641 34051
rect 5629 34020 6316 34048
rect 5629 34017 5641 34020
rect 5583 34011 5641 34017
rect 5810 33940 5816 33992
rect 5868 33940 5874 33992
rect 5828 33912 5856 33940
rect 4724 33884 5856 33912
rect 6288 33912 6316 34020
rect 6454 34008 6460 34060
rect 6512 34008 6518 34060
rect 7929 34051 7987 34057
rect 7929 34017 7941 34051
rect 7975 34048 7987 34051
rect 8294 34048 8300 34060
rect 7975 34020 8300 34048
rect 7975 34017 7987 34020
rect 7929 34011 7987 34017
rect 8294 34008 8300 34020
rect 8352 34048 8358 34060
rect 9140 34048 9168 34076
rect 8352 34020 9168 34048
rect 8352 34008 8358 34020
rect 6914 33980 6920 33992
rect 6875 33952 6920 33980
rect 6914 33940 6920 33952
rect 6972 33940 6978 33992
rect 8846 33980 8852 33992
rect 8807 33952 8852 33980
rect 8846 33940 8852 33952
rect 8904 33940 8910 33992
rect 8941 33983 8999 33989
rect 8941 33949 8953 33983
rect 8987 33980 8999 33983
rect 9122 33980 9128 33992
rect 8987 33952 9128 33980
rect 8987 33949 8999 33952
rect 8941 33943 8999 33949
rect 9122 33940 9128 33952
rect 9180 33980 9186 33992
rect 9508 33980 9536 34088
rect 10381 34085 10393 34088
rect 10427 34085 10439 34119
rect 10381 34079 10439 34085
rect 10597 34119 10655 34125
rect 10597 34085 10609 34119
rect 10643 34085 10655 34119
rect 10597 34079 10655 34085
rect 12802 34076 12808 34128
rect 12860 34116 12866 34128
rect 13446 34116 13452 34128
rect 12860 34088 13452 34116
rect 12860 34076 12866 34088
rect 13446 34076 13452 34088
rect 13504 34076 13510 34128
rect 14826 34076 14832 34128
rect 14884 34116 14890 34128
rect 16298 34116 16304 34128
rect 14884 34088 16304 34116
rect 14884 34076 14890 34088
rect 16298 34076 16304 34088
rect 16356 34076 16362 34128
rect 18506 34076 18512 34128
rect 18564 34116 18570 34128
rect 19886 34116 19892 34128
rect 18564 34088 18920 34116
rect 18564 34076 18570 34088
rect 12345 34051 12403 34057
rect 12345 34017 12357 34051
rect 12391 34048 12403 34051
rect 13354 34048 13360 34060
rect 12391 34020 13360 34048
rect 12391 34017 12403 34020
rect 12345 34011 12403 34017
rect 13354 34008 13360 34020
rect 13412 34008 13418 34060
rect 13722 34008 13728 34060
rect 13780 34048 13786 34060
rect 15841 34051 15899 34057
rect 15841 34048 15853 34051
rect 13780 34020 15853 34048
rect 13780 34008 13786 34020
rect 15841 34017 15853 34020
rect 15887 34048 15899 34051
rect 16206 34048 16212 34060
rect 15887 34020 16212 34048
rect 15887 34017 15899 34020
rect 15841 34011 15899 34017
rect 16206 34008 16212 34020
rect 16264 34008 16270 34060
rect 18892 34057 18920 34088
rect 19076 34088 19892 34116
rect 19076 34057 19104 34088
rect 19886 34076 19892 34088
rect 19944 34076 19950 34128
rect 20622 34116 20628 34128
rect 20180 34088 20628 34116
rect 18693 34051 18751 34057
rect 18693 34017 18705 34051
rect 18739 34017 18751 34051
rect 18693 34011 18751 34017
rect 18877 34051 18935 34057
rect 18877 34017 18889 34051
rect 18923 34017 18935 34051
rect 18877 34011 18935 34017
rect 19061 34051 19119 34057
rect 19061 34017 19073 34051
rect 19107 34017 19119 34051
rect 19061 34011 19119 34017
rect 9180 33952 9536 33980
rect 9180 33940 9186 33952
rect 10226 33940 10232 33992
rect 10284 33980 10290 33992
rect 10284 33952 10456 33980
rect 10284 33940 10290 33952
rect 7282 33912 7288 33924
rect 6288 33884 7288 33912
rect 7282 33872 7288 33884
rect 7340 33872 7346 33924
rect 8113 33915 8171 33921
rect 8113 33881 8125 33915
rect 8159 33912 8171 33915
rect 10318 33912 10324 33924
rect 8159 33884 10324 33912
rect 8159 33881 8171 33884
rect 8113 33875 8171 33881
rect 10318 33872 10324 33884
rect 10376 33872 10382 33924
rect 4706 33844 4712 33856
rect 4448 33816 4712 33844
rect 4706 33804 4712 33816
rect 4764 33804 4770 33856
rect 5626 33804 5632 33856
rect 5684 33844 5690 33856
rect 5813 33847 5871 33853
rect 5813 33844 5825 33847
rect 5684 33816 5825 33844
rect 5684 33804 5690 33816
rect 5813 33813 5825 33816
rect 5859 33813 5871 33847
rect 5813 33807 5871 33813
rect 9401 33847 9459 33853
rect 9401 33813 9413 33847
rect 9447 33844 9459 33847
rect 9582 33844 9588 33856
rect 9447 33816 9588 33844
rect 9447 33813 9459 33816
rect 9401 33807 9459 33813
rect 9582 33804 9588 33816
rect 9640 33804 9646 33856
rect 9766 33804 9772 33856
rect 9824 33844 9830 33856
rect 10428 33853 10456 33952
rect 11974 33940 11980 33992
rect 12032 33980 12038 33992
rect 14826 33980 14832 33992
rect 12032 33952 14832 33980
rect 12032 33940 12038 33952
rect 14826 33940 14832 33952
rect 14884 33940 14890 33992
rect 15102 33980 15108 33992
rect 15063 33952 15108 33980
rect 15102 33940 15108 33952
rect 15160 33940 15166 33992
rect 15286 33940 15292 33992
rect 15344 33980 15350 33992
rect 17770 33980 17776 33992
rect 15344 33952 17776 33980
rect 15344 33940 15350 33952
rect 17770 33940 17776 33952
rect 17828 33940 17834 33992
rect 14734 33872 14740 33924
rect 14792 33912 14798 33924
rect 17313 33915 17371 33921
rect 17313 33912 17325 33915
rect 14792 33884 17325 33912
rect 14792 33872 14798 33884
rect 17313 33881 17325 33884
rect 17359 33912 17371 33915
rect 18598 33912 18604 33924
rect 17359 33884 18604 33912
rect 17359 33881 17371 33884
rect 17313 33875 17371 33881
rect 18598 33872 18604 33884
rect 18656 33872 18662 33924
rect 10229 33847 10287 33853
rect 10229 33844 10241 33847
rect 9824 33816 10241 33844
rect 9824 33804 9830 33816
rect 10229 33813 10241 33816
rect 10275 33813 10287 33847
rect 10229 33807 10287 33813
rect 10413 33847 10471 33853
rect 10413 33813 10425 33847
rect 10459 33844 10471 33847
rect 11514 33844 11520 33856
rect 10459 33816 11520 33844
rect 10459 33813 10471 33816
rect 10413 33807 10471 33813
rect 11514 33804 11520 33816
rect 11572 33804 11578 33856
rect 12066 33844 12072 33856
rect 12027 33816 12072 33844
rect 12066 33804 12072 33816
rect 12124 33804 12130 33856
rect 12986 33844 12992 33856
rect 12899 33816 12992 33844
rect 12986 33804 12992 33816
rect 13044 33844 13050 33856
rect 13630 33844 13636 33856
rect 13044 33816 13636 33844
rect 13044 33804 13050 33816
rect 13630 33804 13636 33816
rect 13688 33804 13694 33856
rect 14918 33804 14924 33856
rect 14976 33844 14982 33856
rect 16761 33847 16819 33853
rect 16761 33844 16773 33847
rect 14976 33816 16773 33844
rect 14976 33804 14982 33816
rect 16761 33813 16773 33816
rect 16807 33844 16819 33847
rect 17218 33844 17224 33856
rect 16807 33816 17224 33844
rect 16807 33813 16819 33816
rect 16761 33807 16819 33813
rect 17218 33804 17224 33816
rect 17276 33804 17282 33856
rect 18708 33844 18736 34011
rect 19150 34008 19156 34060
rect 19208 34048 19214 34060
rect 19245 34051 19303 34057
rect 19245 34048 19257 34051
rect 19208 34020 19257 34048
rect 19208 34008 19214 34020
rect 19245 34017 19257 34020
rect 19291 34048 19303 34051
rect 19794 34048 19800 34060
rect 19291 34020 19800 34048
rect 19291 34017 19303 34020
rect 19245 34011 19303 34017
rect 19794 34008 19800 34020
rect 19852 34008 19858 34060
rect 19981 34051 20039 34057
rect 19981 34017 19993 34051
rect 20027 34048 20039 34051
rect 20070 34048 20076 34060
rect 20027 34020 20076 34048
rect 20027 34017 20039 34020
rect 19981 34011 20039 34017
rect 20070 34008 20076 34020
rect 20128 34008 20134 34060
rect 20180 34057 20208 34088
rect 20622 34076 20628 34088
rect 20680 34116 20686 34128
rect 23658 34116 23664 34128
rect 20680 34088 22048 34116
rect 23619 34088 23664 34116
rect 20680 34076 20686 34088
rect 22020 34057 22048 34088
rect 23658 34076 23664 34088
rect 23716 34076 23722 34128
rect 20165 34051 20223 34057
rect 20165 34017 20177 34051
rect 20211 34017 20223 34051
rect 20165 34011 20223 34017
rect 20533 34051 20591 34057
rect 20533 34017 20545 34051
rect 20579 34017 20591 34051
rect 20533 34011 20591 34017
rect 22005 34051 22063 34057
rect 22005 34017 22017 34051
rect 22051 34017 22063 34051
rect 22370 34048 22376 34060
rect 22331 34020 22376 34048
rect 22005 34011 22063 34017
rect 18969 33983 19027 33989
rect 18969 33949 18981 33983
rect 19015 33949 19027 33983
rect 19334 33980 19340 33992
rect 18969 33943 19027 33949
rect 19260 33952 19340 33980
rect 18984 33912 19012 33943
rect 19058 33912 19064 33924
rect 18984 33884 19064 33912
rect 19058 33872 19064 33884
rect 19116 33912 19122 33924
rect 19260 33912 19288 33952
rect 19334 33940 19340 33952
rect 19392 33980 19398 33992
rect 20257 33983 20315 33989
rect 20257 33980 20269 33983
rect 19392 33952 20269 33980
rect 19392 33940 19398 33952
rect 20257 33949 20269 33952
rect 20303 33949 20315 33983
rect 20257 33943 20315 33949
rect 20349 33983 20407 33989
rect 20349 33949 20361 33983
rect 20395 33949 20407 33983
rect 20548 33980 20576 34011
rect 22370 34008 22376 34020
rect 22428 34008 22434 34060
rect 22557 34051 22615 34057
rect 22557 34017 22569 34051
rect 22603 34048 22615 34051
rect 22646 34048 22652 34060
rect 22603 34020 22652 34048
rect 22603 34017 22615 34020
rect 22557 34011 22615 34017
rect 22646 34008 22652 34020
rect 22704 34008 22710 34060
rect 23860 34048 23888 34147
rect 25590 34144 25596 34196
rect 25648 34184 25654 34196
rect 27522 34184 27528 34196
rect 25648 34156 27384 34184
rect 27483 34156 27528 34184
rect 25648 34144 25654 34156
rect 24305 34119 24363 34125
rect 24305 34085 24317 34119
rect 24351 34116 24363 34119
rect 24578 34116 24584 34128
rect 24351 34088 24584 34116
rect 24351 34085 24363 34088
rect 24305 34079 24363 34085
rect 24578 34076 24584 34088
rect 24636 34076 24642 34128
rect 25406 34076 25412 34128
rect 25464 34116 25470 34128
rect 25777 34119 25835 34125
rect 25777 34116 25789 34119
rect 25464 34088 25789 34116
rect 25464 34076 25470 34088
rect 25777 34085 25789 34088
rect 25823 34085 25835 34119
rect 25777 34079 25835 34085
rect 26050 34076 26056 34128
rect 26108 34116 26114 34128
rect 26154 34119 26212 34125
rect 26154 34116 26166 34119
rect 26108 34088 26166 34116
rect 26108 34076 26114 34088
rect 26154 34085 26166 34088
rect 26200 34085 26212 34119
rect 26154 34079 26212 34085
rect 25133 34051 25191 34057
rect 25133 34048 25145 34051
rect 23860 34020 25145 34048
rect 25133 34017 25145 34020
rect 25179 34017 25191 34051
rect 26510 34048 26516 34060
rect 25133 34011 25191 34017
rect 25240 34020 26516 34048
rect 21910 33980 21916 33992
rect 20548 33952 21916 33980
rect 20349 33943 20407 33949
rect 19116 33884 19288 33912
rect 19116 33872 19122 33884
rect 19886 33872 19892 33924
rect 19944 33912 19950 33924
rect 20364 33912 20392 33943
rect 21910 33940 21916 33952
rect 21968 33940 21974 33992
rect 22189 33983 22247 33989
rect 22189 33949 22201 33983
rect 22235 33949 22247 33983
rect 22189 33943 22247 33949
rect 19944 33884 20392 33912
rect 19944 33872 19950 33884
rect 20530 33872 20536 33924
rect 20588 33912 20594 33924
rect 21177 33915 21235 33921
rect 21177 33912 21189 33915
rect 20588 33884 21189 33912
rect 20588 33872 20594 33884
rect 21177 33881 21189 33884
rect 21223 33881 21235 33915
rect 22204 33912 22232 33943
rect 22278 33940 22284 33992
rect 22336 33980 22342 33992
rect 23382 33980 23388 33992
rect 22336 33952 23388 33980
rect 22336 33940 22342 33952
rect 23382 33940 23388 33952
rect 23440 33940 23446 33992
rect 24762 33940 24768 33992
rect 24820 33980 24826 33992
rect 24857 33983 24915 33989
rect 24857 33980 24869 33983
rect 24820 33952 24869 33980
rect 24820 33940 24826 33952
rect 24857 33949 24869 33952
rect 24903 33980 24915 33983
rect 25240 33980 25268 34020
rect 26510 34008 26516 34020
rect 26568 34008 26574 34060
rect 27356 34048 27384 34156
rect 27522 34144 27528 34156
rect 27580 34144 27586 34196
rect 27706 34144 27712 34196
rect 27764 34184 27770 34196
rect 28169 34187 28227 34193
rect 28169 34184 28181 34187
rect 27764 34156 28181 34184
rect 27764 34144 27770 34156
rect 28169 34153 28181 34156
rect 28215 34153 28227 34187
rect 29730 34184 29736 34196
rect 29691 34156 29736 34184
rect 28169 34147 28227 34153
rect 29730 34144 29736 34156
rect 29788 34144 29794 34196
rect 29914 34144 29920 34196
rect 29972 34184 29978 34196
rect 30285 34187 30343 34193
rect 30285 34184 30297 34187
rect 29972 34156 30297 34184
rect 29972 34144 29978 34156
rect 30285 34153 30297 34156
rect 30331 34153 30343 34187
rect 30285 34147 30343 34153
rect 27433 34051 27491 34057
rect 27433 34048 27445 34051
rect 27356 34020 27445 34048
rect 27433 34017 27445 34020
rect 27479 34048 27491 34051
rect 27982 34048 27988 34060
rect 27479 34020 27988 34048
rect 27479 34017 27491 34020
rect 27433 34011 27491 34017
rect 27982 34008 27988 34020
rect 28040 34008 28046 34060
rect 28261 34051 28319 34057
rect 28261 34017 28273 34051
rect 28307 34048 28319 34051
rect 28350 34048 28356 34060
rect 28307 34020 28356 34048
rect 28307 34017 28319 34020
rect 28261 34011 28319 34017
rect 28350 34008 28356 34020
rect 28408 34008 28414 34060
rect 28810 34008 28816 34060
rect 28868 34048 28874 34060
rect 28997 34051 29055 34057
rect 28997 34048 29009 34051
rect 28868 34020 29009 34048
rect 28868 34008 28874 34020
rect 28997 34017 29009 34020
rect 29043 34017 29055 34051
rect 29178 34048 29184 34060
rect 29139 34020 29184 34048
rect 28997 34011 29055 34017
rect 29178 34008 29184 34020
rect 29236 34008 29242 34060
rect 29270 34008 29276 34060
rect 29328 34048 29334 34060
rect 29546 34048 29552 34060
rect 29328 34020 29373 34048
rect 29507 34020 29552 34048
rect 29328 34008 29334 34020
rect 29546 34008 29552 34020
rect 29604 34008 29610 34060
rect 30006 34008 30012 34060
rect 30064 34048 30070 34060
rect 30377 34051 30435 34057
rect 30377 34048 30389 34051
rect 30064 34020 30389 34048
rect 30064 34008 30070 34020
rect 30377 34017 30389 34020
rect 30423 34017 30435 34051
rect 30377 34011 30435 34017
rect 31113 34051 31171 34057
rect 31113 34017 31125 34051
rect 31159 34048 31171 34051
rect 31662 34048 31668 34060
rect 31159 34020 31668 34048
rect 31159 34017 31171 34020
rect 31113 34011 31171 34017
rect 31662 34008 31668 34020
rect 31720 34008 31726 34060
rect 24903 33952 25268 33980
rect 25317 33983 25375 33989
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 25317 33949 25329 33983
rect 25363 33980 25375 33983
rect 25363 33952 26372 33980
rect 25363 33949 25375 33952
rect 25317 33943 25375 33949
rect 23014 33912 23020 33924
rect 22204 33884 23020 33912
rect 21177 33875 21235 33881
rect 23014 33872 23020 33884
rect 23072 33872 23078 33924
rect 23293 33915 23351 33921
rect 23293 33881 23305 33915
rect 23339 33881 23351 33915
rect 23293 33875 23351 33881
rect 19702 33844 19708 33856
rect 18708 33816 19708 33844
rect 19702 33804 19708 33816
rect 19760 33844 19766 33856
rect 20162 33844 20168 33856
rect 19760 33816 20168 33844
rect 19760 33804 19766 33816
rect 20162 33804 20168 33816
rect 20220 33804 20226 33856
rect 21821 33847 21879 33853
rect 21821 33813 21833 33847
rect 21867 33844 21879 33847
rect 21910 33844 21916 33856
rect 21867 33816 21916 33844
rect 21867 33813 21879 33816
rect 21821 33807 21879 33813
rect 21910 33804 21916 33816
rect 21968 33804 21974 33856
rect 22370 33804 22376 33856
rect 22428 33844 22434 33856
rect 22830 33844 22836 33856
rect 22428 33816 22836 33844
rect 22428 33804 22434 33816
rect 22830 33804 22836 33816
rect 22888 33804 22894 33856
rect 23308 33844 23336 33875
rect 25222 33872 25228 33924
rect 25280 33912 25286 33924
rect 25866 33912 25872 33924
rect 25280 33884 25872 33912
rect 25280 33872 25286 33884
rect 25866 33872 25872 33884
rect 25924 33872 25930 33924
rect 26344 33921 26372 33952
rect 29086 33940 29092 33992
rect 29144 33980 29150 33992
rect 29365 33983 29423 33989
rect 29365 33980 29377 33983
rect 29144 33952 29377 33980
rect 29144 33940 29150 33952
rect 29365 33949 29377 33952
rect 29411 33949 29423 33983
rect 29365 33943 29423 33949
rect 26329 33915 26387 33921
rect 26329 33881 26341 33915
rect 26375 33881 26387 33915
rect 26329 33875 26387 33881
rect 23382 33844 23388 33856
rect 23308 33816 23388 33844
rect 23382 33804 23388 33816
rect 23440 33804 23446 33856
rect 23661 33847 23719 33853
rect 23661 33813 23673 33847
rect 23707 33844 23719 33847
rect 25406 33844 25412 33856
rect 23707 33816 25412 33844
rect 23707 33813 23719 33816
rect 23661 33807 23719 33813
rect 25406 33804 25412 33816
rect 25464 33804 25470 33856
rect 26142 33844 26148 33856
rect 26103 33816 26148 33844
rect 26142 33804 26148 33816
rect 26200 33804 26206 33856
rect 31297 33847 31355 33853
rect 31297 33813 31309 33847
rect 31343 33844 31355 33847
rect 31343 33816 32076 33844
rect 31343 33813 31355 33816
rect 31297 33807 31355 33813
rect 0 33680 888 33708
rect 1104 33754 32016 33776
rect 1104 33702 6102 33754
rect 6154 33702 6166 33754
rect 6218 33702 6230 33754
rect 6282 33702 6294 33754
rect 6346 33702 6358 33754
rect 6410 33702 16405 33754
rect 16457 33702 16469 33754
rect 16521 33702 16533 33754
rect 16585 33702 16597 33754
rect 16649 33702 16661 33754
rect 16713 33702 26709 33754
rect 26761 33702 26773 33754
rect 26825 33702 26837 33754
rect 26889 33702 26901 33754
rect 26953 33702 26965 33754
rect 27017 33702 32016 33754
rect 1104 33680 32016 33702
rect 32048 33708 32076 33816
rect 32320 33708 33120 33722
rect 32048 33680 33120 33708
rect 0 33666 800 33680
rect 32320 33666 33120 33680
rect 3053 33643 3111 33649
rect 3053 33609 3065 33643
rect 3099 33640 3111 33643
rect 4522 33640 4528 33652
rect 3099 33612 4528 33640
rect 3099 33609 3111 33612
rect 3053 33603 3111 33609
rect 4522 33600 4528 33612
rect 4580 33640 4586 33652
rect 5442 33640 5448 33652
rect 4580 33612 5448 33640
rect 4580 33600 4586 33612
rect 5442 33600 5448 33612
rect 5500 33600 5506 33652
rect 5994 33600 6000 33652
rect 6052 33640 6058 33652
rect 6457 33643 6515 33649
rect 6457 33640 6469 33643
rect 6052 33612 6469 33640
rect 6052 33600 6058 33612
rect 6457 33609 6469 33612
rect 6503 33609 6515 33643
rect 6457 33603 6515 33609
rect 11790 33600 11796 33652
rect 11848 33640 11854 33652
rect 13170 33640 13176 33652
rect 11848 33612 13176 33640
rect 11848 33600 11854 33612
rect 13170 33600 13176 33612
rect 13228 33600 13234 33652
rect 13354 33600 13360 33652
rect 13412 33640 13418 33652
rect 13449 33643 13507 33649
rect 13449 33640 13461 33643
rect 13412 33612 13461 33640
rect 13412 33600 13418 33612
rect 13449 33609 13461 33612
rect 13495 33640 13507 33643
rect 18782 33640 18788 33652
rect 13495 33612 18788 33640
rect 13495 33609 13507 33612
rect 13449 33603 13507 33609
rect 18782 33600 18788 33612
rect 18840 33600 18846 33652
rect 19794 33600 19800 33652
rect 19852 33640 19858 33652
rect 19852 33612 20484 33640
rect 19852 33600 19858 33612
rect 2406 33572 2412 33584
rect 2056 33544 2412 33572
rect 2056 33448 2084 33544
rect 2406 33532 2412 33544
rect 2464 33532 2470 33584
rect 4246 33572 4252 33584
rect 2516 33544 4252 33572
rect 2516 33504 2544 33544
rect 4246 33532 4252 33544
rect 4304 33532 4310 33584
rect 5258 33532 5264 33584
rect 5316 33572 5322 33584
rect 5316 33544 5672 33572
rect 5316 33532 5322 33544
rect 3142 33504 3148 33516
rect 2148 33476 2544 33504
rect 2884 33476 3148 33504
rect 2038 33436 2044 33448
rect 1951 33408 2044 33436
rect 2038 33396 2044 33408
rect 2096 33396 2102 33448
rect 2148 33445 2176 33476
rect 2133 33439 2191 33445
rect 2133 33405 2145 33439
rect 2179 33405 2191 33439
rect 2133 33399 2191 33405
rect 2225 33439 2283 33445
rect 2225 33405 2237 33439
rect 2271 33405 2283 33439
rect 2225 33399 2283 33405
rect 2409 33439 2467 33445
rect 2409 33405 2421 33439
rect 2455 33436 2467 33439
rect 2884 33436 2912 33476
rect 3142 33464 3148 33476
rect 3200 33464 3206 33516
rect 2455 33408 2912 33436
rect 2455 33405 2467 33408
rect 2409 33399 2467 33405
rect 2240 33368 2268 33399
rect 3050 33396 3056 33448
rect 3108 33436 3114 33448
rect 5644 33445 5672 33544
rect 5718 33532 5724 33584
rect 5776 33572 5782 33584
rect 7285 33575 7343 33581
rect 7285 33572 7297 33575
rect 5776 33544 7297 33572
rect 5776 33532 5782 33544
rect 7285 33541 7297 33544
rect 7331 33572 7343 33575
rect 7331 33544 7788 33572
rect 7331 33541 7343 33544
rect 7285 33535 7343 33541
rect 7558 33504 7564 33516
rect 6196 33476 7564 33504
rect 3789 33439 3847 33445
rect 3789 33436 3801 33439
rect 3108 33408 3801 33436
rect 3108 33396 3114 33408
rect 3789 33405 3801 33408
rect 3835 33405 3847 33439
rect 3789 33399 3847 33405
rect 5425 33439 5483 33445
rect 5425 33405 5437 33439
rect 5471 33436 5483 33439
rect 5537 33439 5595 33445
rect 5471 33405 5488 33436
rect 5425 33399 5488 33405
rect 5537 33405 5549 33439
rect 5583 33405 5595 33439
rect 5537 33399 5595 33405
rect 5629 33439 5687 33445
rect 5629 33405 5641 33439
rect 5675 33405 5687 33439
rect 5810 33436 5816 33448
rect 5771 33408 5816 33436
rect 5629 33399 5687 33405
rect 2590 33368 2596 33380
rect 2148 33340 2596 33368
rect 2148 33312 2176 33340
rect 2590 33328 2596 33340
rect 2648 33328 2654 33380
rect 2866 33368 2872 33380
rect 2827 33340 2872 33368
rect 2866 33328 2872 33340
rect 2924 33328 2930 33380
rect 3326 33368 3332 33380
rect 3068 33340 3332 33368
rect 1765 33303 1823 33309
rect 1765 33269 1777 33303
rect 1811 33300 1823 33303
rect 1946 33300 1952 33312
rect 1811 33272 1952 33300
rect 1811 33269 1823 33272
rect 1765 33263 1823 33269
rect 1946 33260 1952 33272
rect 2004 33260 2010 33312
rect 2130 33260 2136 33312
rect 2188 33260 2194 33312
rect 3068 33309 3096 33340
rect 3326 33328 3332 33340
rect 3384 33328 3390 33380
rect 3068 33303 3127 33309
rect 3068 33272 3081 33303
rect 3069 33269 3081 33272
rect 3115 33269 3127 33303
rect 3234 33300 3240 33312
rect 3195 33272 3240 33300
rect 3069 33263 3127 33269
rect 3234 33260 3240 33272
rect 3292 33260 3298 33312
rect 3878 33300 3884 33312
rect 3839 33272 3884 33300
rect 3878 33260 3884 33272
rect 3936 33260 3942 33312
rect 4890 33260 4896 33312
rect 4948 33300 4954 33312
rect 5169 33303 5227 33309
rect 5169 33300 5181 33303
rect 4948 33272 5181 33300
rect 4948 33260 4954 33272
rect 5169 33269 5181 33272
rect 5215 33269 5227 33303
rect 5460 33300 5488 33399
rect 5552 33368 5580 33399
rect 5810 33396 5816 33408
rect 5868 33396 5874 33448
rect 5718 33368 5724 33380
rect 5552 33340 5724 33368
rect 5718 33328 5724 33340
rect 5776 33368 5782 33380
rect 6196 33368 6224 33476
rect 7558 33464 7564 33476
rect 7616 33464 7622 33516
rect 7282 33436 7288 33448
rect 6288 33408 7288 33436
rect 6288 33377 6316 33408
rect 7282 33396 7288 33408
rect 7340 33396 7346 33448
rect 7760 33445 7788 33544
rect 10042 33532 10048 33584
rect 10100 33572 10106 33584
rect 10689 33575 10747 33581
rect 10689 33572 10701 33575
rect 10100 33544 10701 33572
rect 10100 33532 10106 33544
rect 10689 33541 10701 33544
rect 10735 33541 10747 33575
rect 10689 33535 10747 33541
rect 11716 33544 12756 33572
rect 9309 33507 9367 33513
rect 9309 33504 9321 33507
rect 8772 33476 9321 33504
rect 7653 33439 7711 33445
rect 7653 33405 7665 33439
rect 7699 33405 7711 33439
rect 7653 33399 7711 33405
rect 7745 33439 7803 33445
rect 7745 33405 7757 33439
rect 7791 33405 7803 33439
rect 7745 33399 7803 33405
rect 5776 33340 6224 33368
rect 6273 33371 6331 33377
rect 5776 33328 5782 33340
rect 6273 33337 6285 33371
rect 6319 33337 6331 33371
rect 6273 33331 6331 33337
rect 6288 33300 6316 33331
rect 6454 33328 6460 33380
rect 6512 33377 6518 33380
rect 6512 33371 6531 33377
rect 6519 33337 6531 33371
rect 7668 33368 7696 33399
rect 7834 33396 7840 33448
rect 7892 33436 7898 33448
rect 8021 33439 8079 33445
rect 7892 33408 7937 33436
rect 7892 33396 7898 33408
rect 8021 33405 8033 33439
rect 8067 33436 8079 33439
rect 8662 33436 8668 33448
rect 8067 33408 8668 33436
rect 8067 33405 8079 33408
rect 8021 33399 8079 33405
rect 8662 33396 8668 33408
rect 8720 33396 8726 33448
rect 8772 33368 8800 33476
rect 9309 33473 9321 33476
rect 9355 33504 9367 33507
rect 9766 33504 9772 33516
rect 9355 33476 9674 33504
rect 9727 33476 9772 33504
rect 9355 33473 9367 33476
rect 9309 33467 9367 33473
rect 9646 33448 9674 33476
rect 9766 33464 9772 33476
rect 9824 33464 9830 33516
rect 11146 33464 11152 33516
rect 11204 33504 11210 33516
rect 11716 33504 11744 33544
rect 11974 33504 11980 33516
rect 11204 33476 11744 33504
rect 11935 33476 11980 33504
rect 11204 33464 11210 33476
rect 8938 33436 8944 33448
rect 8899 33408 8944 33436
rect 8938 33396 8944 33408
rect 8996 33396 9002 33448
rect 9214 33436 9220 33448
rect 9175 33408 9220 33436
rect 9214 33396 9220 33408
rect 9272 33396 9278 33448
rect 9646 33408 9680 33448
rect 9674 33396 9680 33408
rect 9732 33396 9738 33448
rect 10686 33436 10692 33448
rect 10647 33408 10692 33436
rect 10686 33396 10692 33408
rect 10744 33396 10750 33448
rect 11716 33445 11744 33476
rect 11974 33464 11980 33476
rect 12032 33464 12038 33516
rect 12084 33476 12664 33504
rect 10873 33439 10931 33445
rect 10873 33405 10885 33439
rect 10919 33436 10931 33439
rect 11517 33439 11575 33445
rect 11517 33436 11529 33439
rect 10919 33408 11529 33436
rect 10919 33405 10931 33408
rect 10873 33399 10931 33405
rect 11517 33405 11529 33408
rect 11563 33405 11575 33439
rect 11517 33399 11575 33405
rect 11701 33439 11759 33445
rect 11701 33405 11713 33439
rect 11747 33405 11759 33439
rect 11701 33399 11759 33405
rect 11790 33396 11796 33448
rect 11848 33436 11854 33448
rect 12084 33445 12112 33476
rect 11885 33439 11943 33445
rect 11885 33436 11897 33439
rect 11848 33408 11897 33436
rect 11848 33396 11854 33408
rect 11885 33405 11897 33408
rect 11931 33405 11943 33439
rect 11885 33399 11943 33405
rect 12069 33439 12127 33445
rect 12069 33405 12081 33439
rect 12115 33405 12127 33439
rect 12250 33436 12256 33448
rect 12211 33408 12256 33436
rect 12069 33399 12127 33405
rect 12250 33396 12256 33408
rect 12308 33396 12314 33448
rect 7668 33340 8800 33368
rect 6512 33331 6531 33337
rect 6512 33328 6518 33331
rect 8036 33312 8064 33340
rect 9306 33328 9312 33380
rect 9364 33368 9370 33380
rect 9585 33371 9643 33377
rect 9585 33368 9597 33371
rect 9364 33340 9597 33368
rect 9364 33328 9370 33340
rect 9585 33337 9597 33340
rect 9631 33337 9643 33371
rect 9585 33331 9643 33337
rect 11057 33371 11115 33377
rect 11057 33337 11069 33371
rect 11103 33337 11115 33371
rect 12636 33368 12664 33476
rect 12728 33445 12756 33544
rect 17218 33532 17224 33584
rect 17276 33572 17282 33584
rect 20456 33581 20484 33612
rect 20530 33600 20536 33652
rect 20588 33640 20594 33652
rect 20809 33643 20867 33649
rect 20809 33640 20821 33643
rect 20588 33612 20821 33640
rect 20588 33600 20594 33612
rect 20809 33609 20821 33612
rect 20855 33609 20867 33643
rect 21450 33640 21456 33652
rect 21411 33612 21456 33640
rect 20809 33603 20867 33609
rect 21450 33600 21456 33612
rect 21508 33600 21514 33652
rect 30745 33643 30803 33649
rect 30745 33640 30757 33643
rect 21560 33612 30757 33640
rect 20441 33575 20499 33581
rect 17276 33544 20116 33572
rect 17276 33532 17282 33544
rect 15102 33464 15108 33516
rect 15160 33504 15166 33516
rect 15933 33507 15991 33513
rect 15933 33504 15945 33507
rect 15160 33476 15945 33504
rect 15160 33464 15166 33476
rect 15933 33473 15945 33476
rect 15979 33473 15991 33507
rect 15933 33467 15991 33473
rect 19242 33464 19248 33516
rect 19300 33504 19306 33516
rect 19515 33507 19573 33513
rect 19515 33504 19527 33507
rect 19300 33476 19527 33504
rect 19300 33464 19306 33476
rect 19515 33473 19527 33476
rect 19561 33473 19573 33507
rect 19978 33504 19984 33516
rect 19515 33467 19573 33473
rect 19720 33476 19984 33504
rect 12713 33439 12771 33445
rect 12713 33405 12725 33439
rect 12759 33405 12771 33439
rect 14090 33436 14096 33448
rect 14003 33408 14096 33436
rect 12713 33399 12771 33405
rect 14090 33396 14096 33408
rect 14148 33436 14154 33448
rect 15120 33436 15148 33464
rect 17773 33439 17831 33445
rect 17773 33436 17785 33439
rect 14148 33408 15148 33436
rect 16408 33408 17785 33436
rect 14148 33396 14154 33408
rect 12805 33371 12863 33377
rect 12805 33368 12817 33371
rect 12636 33340 12817 33368
rect 11057 33331 11115 33337
rect 12805 33337 12817 33340
rect 12851 33337 12863 33371
rect 12805 33331 12863 33337
rect 5460 33272 6316 33300
rect 6641 33303 6699 33309
rect 5169 33263 5227 33269
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 7098 33300 7104 33312
rect 6687 33272 7104 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 7098 33260 7104 33272
rect 7156 33260 7162 33312
rect 7282 33300 7288 33312
rect 7243 33272 7288 33300
rect 7282 33260 7288 33272
rect 7340 33260 7346 33312
rect 7377 33303 7435 33309
rect 7377 33269 7389 33303
rect 7423 33300 7435 33303
rect 7558 33300 7564 33312
rect 7423 33272 7564 33300
rect 7423 33269 7435 33272
rect 7377 33263 7435 33269
rect 7558 33260 7564 33272
rect 7616 33260 7622 33312
rect 8018 33260 8024 33312
rect 8076 33260 8082 33312
rect 11072 33300 11100 33331
rect 13814 33328 13820 33380
rect 13872 33368 13878 33380
rect 14338 33371 14396 33377
rect 14338 33368 14350 33371
rect 13872 33340 14350 33368
rect 13872 33328 13878 33340
rect 14338 33337 14350 33340
rect 14384 33337 14396 33371
rect 14338 33331 14396 33337
rect 15746 33328 15752 33380
rect 15804 33368 15810 33380
rect 16178 33371 16236 33377
rect 16178 33368 16190 33371
rect 15804 33340 16190 33368
rect 15804 33328 15810 33340
rect 16178 33337 16190 33340
rect 16224 33337 16236 33371
rect 16178 33331 16236 33337
rect 16298 33328 16304 33380
rect 16356 33368 16362 33380
rect 16408 33368 16436 33408
rect 17773 33405 17785 33408
rect 17819 33405 17831 33439
rect 18506 33436 18512 33448
rect 18467 33408 18512 33436
rect 17773 33399 17831 33405
rect 18506 33396 18512 33408
rect 18564 33396 18570 33448
rect 19150 33396 19156 33448
rect 19208 33436 19214 33448
rect 19208 33435 19288 33436
rect 19208 33429 19307 33435
rect 19208 33408 19261 33429
rect 19208 33396 19214 33408
rect 19249 33395 19261 33408
rect 19295 33395 19307 33429
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 19720 33446 19748 33476
rect 19978 33464 19984 33476
rect 20036 33464 20042 33516
rect 20088 33504 20116 33544
rect 20441 33541 20453 33575
rect 20487 33541 20499 33575
rect 21560 33572 21588 33612
rect 30745 33609 30757 33612
rect 30791 33609 30803 33643
rect 30745 33603 30803 33609
rect 25590 33572 25596 33584
rect 20441 33535 20499 33541
rect 20548 33544 21588 33572
rect 24964 33544 25596 33572
rect 20548 33504 20576 33544
rect 20088 33476 20576 33504
rect 20622 33464 20628 33516
rect 20680 33504 20686 33516
rect 21729 33507 21787 33513
rect 21729 33504 21741 33507
rect 20680 33476 21741 33504
rect 20680 33464 20686 33476
rect 21729 33473 21741 33476
rect 21775 33473 21787 33507
rect 21910 33504 21916 33516
rect 21871 33476 21916 33504
rect 21729 33467 21787 33473
rect 21910 33464 21916 33476
rect 21968 33464 21974 33516
rect 23198 33504 23204 33516
rect 23159 33476 23204 33504
rect 23198 33464 23204 33476
rect 23256 33464 23262 33516
rect 19628 33445 19748 33446
rect 19613 33439 19748 33445
rect 19484 33408 19529 33436
rect 19484 33396 19490 33408
rect 19613 33405 19625 33439
rect 19659 33418 19748 33439
rect 19659 33405 19671 33418
rect 19613 33399 19671 33405
rect 19794 33396 19800 33448
rect 19852 33436 19858 33448
rect 19852 33408 19897 33436
rect 19852 33396 19858 33408
rect 20070 33396 20076 33448
rect 20128 33436 20134 33448
rect 20898 33436 20904 33448
rect 20128 33408 20904 33436
rect 20128 33396 20134 33408
rect 20898 33396 20904 33408
rect 20956 33436 20962 33448
rect 21637 33439 21695 33445
rect 21637 33436 21649 33439
rect 20956 33408 21649 33436
rect 20956 33396 20962 33408
rect 21637 33405 21649 33408
rect 21683 33405 21695 33439
rect 21818 33436 21824 33448
rect 21779 33408 21824 33436
rect 21637 33399 21695 33405
rect 21818 33396 21824 33408
rect 21876 33396 21882 33448
rect 22738 33396 22744 33448
rect 22796 33436 22802 33448
rect 22925 33439 22983 33445
rect 22925 33436 22937 33439
rect 22796 33408 22937 33436
rect 22796 33396 22802 33408
rect 22925 33405 22937 33408
rect 22971 33436 22983 33439
rect 24486 33436 24492 33448
rect 22971 33408 24492 33436
rect 22971 33405 22983 33408
rect 22925 33399 22983 33405
rect 24486 33396 24492 33408
rect 24544 33396 24550 33448
rect 24765 33439 24823 33445
rect 24765 33405 24777 33439
rect 24811 33436 24823 33439
rect 24854 33436 24860 33448
rect 24811 33408 24860 33436
rect 24811 33405 24823 33408
rect 24765 33399 24823 33405
rect 24854 33396 24860 33408
rect 24912 33396 24918 33448
rect 24964 33445 24992 33544
rect 25590 33532 25596 33544
rect 25648 33532 25654 33584
rect 25961 33575 26019 33581
rect 25961 33541 25973 33575
rect 26007 33541 26019 33575
rect 25961 33535 26019 33541
rect 25041 33507 25099 33513
rect 25041 33473 25053 33507
rect 25087 33504 25099 33507
rect 25222 33504 25228 33516
rect 25087 33476 25228 33504
rect 25087 33473 25099 33476
rect 25041 33467 25099 33473
rect 25222 33464 25228 33476
rect 25280 33464 25286 33516
rect 25976 33504 26004 33535
rect 29086 33532 29092 33584
rect 29144 33572 29150 33584
rect 29730 33572 29736 33584
rect 29144 33544 29736 33572
rect 29144 33532 29150 33544
rect 29730 33532 29736 33544
rect 29788 33572 29794 33584
rect 29788 33544 29960 33572
rect 29788 33532 29794 33544
rect 25608 33476 26004 33504
rect 25608 33448 25636 33476
rect 28074 33464 28080 33516
rect 28132 33504 28138 33516
rect 28169 33507 28227 33513
rect 28169 33504 28181 33507
rect 28132 33476 28181 33504
rect 28132 33464 28138 33476
rect 28169 33473 28181 33476
rect 28215 33473 28227 33507
rect 28169 33467 28227 33473
rect 28261 33507 28319 33513
rect 28261 33473 28273 33507
rect 28307 33504 28319 33507
rect 29270 33504 29276 33516
rect 28307 33476 29276 33504
rect 28307 33473 28319 33476
rect 28261 33467 28319 33473
rect 29270 33464 29276 33476
rect 29328 33504 29334 33516
rect 29822 33504 29828 33516
rect 29328 33476 29828 33504
rect 29328 33464 29334 33476
rect 29822 33464 29828 33476
rect 29880 33464 29886 33516
rect 29932 33513 29960 33544
rect 29917 33507 29975 33513
rect 29917 33473 29929 33507
rect 29963 33473 29975 33507
rect 29917 33467 29975 33473
rect 24949 33439 25007 33445
rect 24949 33405 24961 33439
rect 24995 33405 25007 33439
rect 24949 33399 25007 33405
rect 25133 33439 25191 33445
rect 25133 33405 25145 33439
rect 25179 33405 25191 33439
rect 25133 33399 25191 33405
rect 25317 33439 25375 33445
rect 25317 33405 25329 33439
rect 25363 33436 25375 33439
rect 25590 33436 25596 33448
rect 25363 33408 25596 33436
rect 25363 33405 25375 33408
rect 25317 33399 25375 33405
rect 19249 33389 19307 33395
rect 16356 33340 16436 33368
rect 16356 33328 16362 33340
rect 16758 33328 16764 33380
rect 16816 33368 16822 33380
rect 17865 33371 17923 33377
rect 17865 33368 17877 33371
rect 16816 33340 17877 33368
rect 16816 33328 16822 33340
rect 17865 33337 17877 33340
rect 17911 33337 17923 33371
rect 17865 33331 17923 33337
rect 18601 33371 18659 33377
rect 18601 33337 18613 33371
rect 18647 33368 18659 33371
rect 20530 33368 20536 33380
rect 18647 33340 19104 33368
rect 18647 33337 18659 33340
rect 18601 33331 18659 33337
rect 14918 33300 14924 33312
rect 11072 33272 14924 33300
rect 14918 33260 14924 33272
rect 14976 33260 14982 33312
rect 15194 33260 15200 33312
rect 15252 33300 15258 33312
rect 15473 33303 15531 33309
rect 15473 33300 15485 33303
rect 15252 33272 15485 33300
rect 15252 33260 15258 33272
rect 15473 33269 15485 33272
rect 15519 33269 15531 33303
rect 17310 33300 17316 33312
rect 17271 33272 17316 33300
rect 15473 33263 15531 33269
rect 17310 33260 17316 33272
rect 17368 33260 17374 33312
rect 17770 33260 17776 33312
rect 17828 33300 17834 33312
rect 18782 33300 18788 33312
rect 17828 33272 18788 33300
rect 17828 33260 17834 33272
rect 18782 33260 18788 33272
rect 18840 33260 18846 33312
rect 19076 33300 19104 33340
rect 19812 33340 20536 33368
rect 19518 33300 19524 33312
rect 19076 33272 19524 33300
rect 19518 33260 19524 33272
rect 19576 33260 19582 33312
rect 19702 33260 19708 33312
rect 19760 33300 19766 33312
rect 19812 33300 19840 33340
rect 20530 33328 20536 33340
rect 20588 33328 20594 33380
rect 23198 33328 23204 33380
rect 23256 33368 23262 33380
rect 23382 33368 23388 33380
rect 23256 33340 23388 33368
rect 23256 33328 23262 33340
rect 23382 33328 23388 33340
rect 23440 33328 23446 33380
rect 25148 33368 25176 33399
rect 25590 33396 25596 33408
rect 25648 33396 25654 33448
rect 25893 33408 26197 33436
rect 25222 33368 25228 33380
rect 25148 33340 25228 33368
rect 25222 33328 25228 33340
rect 25280 33368 25286 33380
rect 25774 33368 25780 33380
rect 25280 33340 25780 33368
rect 25280 33328 25286 33340
rect 25774 33328 25780 33340
rect 25832 33328 25838 33380
rect 19760 33272 19840 33300
rect 19981 33303 20039 33309
rect 19760 33260 19766 33272
rect 19981 33269 19993 33303
rect 20027 33300 20039 33303
rect 20622 33300 20628 33312
rect 20027 33272 20628 33300
rect 20027 33269 20039 33272
rect 19981 33263 20039 33269
rect 20622 33260 20628 33272
rect 20680 33260 20686 33312
rect 20806 33300 20812 33312
rect 20767 33272 20812 33300
rect 20806 33260 20812 33272
rect 20864 33260 20870 33312
rect 20898 33260 20904 33312
rect 20956 33300 20962 33312
rect 20993 33303 21051 33309
rect 20993 33300 21005 33303
rect 20956 33272 21005 33300
rect 20956 33260 20962 33272
rect 20993 33269 21005 33272
rect 21039 33269 21051 33303
rect 20993 33263 21051 33269
rect 21174 33260 21180 33312
rect 21232 33300 21238 33312
rect 21450 33300 21456 33312
rect 21232 33272 21456 33300
rect 21232 33260 21238 33272
rect 21450 33260 21456 33272
rect 21508 33260 21514 33312
rect 21910 33260 21916 33312
rect 21968 33300 21974 33312
rect 23750 33300 23756 33312
rect 21968 33272 23756 33300
rect 21968 33260 21974 33272
rect 23750 33260 23756 33272
rect 23808 33300 23814 33312
rect 24578 33300 24584 33312
rect 23808 33272 24584 33300
rect 23808 33260 23814 33272
rect 24578 33260 24584 33272
rect 24636 33260 24642 33312
rect 25038 33260 25044 33312
rect 25096 33300 25102 33312
rect 25406 33300 25412 33312
rect 25096 33272 25412 33300
rect 25096 33260 25102 33272
rect 25406 33260 25412 33272
rect 25464 33260 25470 33312
rect 25501 33303 25559 33309
rect 25501 33269 25513 33303
rect 25547 33300 25559 33303
rect 25893 33300 25921 33408
rect 26169 33368 26197 33408
rect 26234 33396 26240 33448
rect 26292 33436 26298 33448
rect 27341 33439 27399 33445
rect 27341 33436 27353 33439
rect 26292 33408 27353 33436
rect 26292 33396 26298 33408
rect 27341 33405 27353 33408
rect 27387 33405 27399 33439
rect 27982 33436 27988 33448
rect 27943 33408 27988 33436
rect 27341 33399 27399 33405
rect 27982 33396 27988 33408
rect 28040 33396 28046 33448
rect 28350 33396 28356 33448
rect 28408 33436 28414 33448
rect 28537 33439 28595 33445
rect 28408 33408 28453 33436
rect 28408 33396 28414 33408
rect 28537 33405 28549 33439
rect 28583 33436 28595 33439
rect 28626 33436 28632 33448
rect 28583 33408 28632 33436
rect 28583 33405 28595 33408
rect 28537 33399 28595 33405
rect 28626 33396 28632 33408
rect 28684 33436 28690 33448
rect 28810 33436 28816 33448
rect 28684 33408 28816 33436
rect 28684 33396 28690 33408
rect 28810 33396 28816 33408
rect 28868 33436 28874 33448
rect 29549 33439 29607 33445
rect 29549 33436 29561 33439
rect 28868 33408 29561 33436
rect 28868 33396 28874 33408
rect 29549 33405 29561 33408
rect 29595 33405 29607 33439
rect 29549 33399 29607 33405
rect 29638 33396 29644 33448
rect 29696 33436 29702 33448
rect 29733 33439 29791 33445
rect 29733 33436 29745 33439
rect 29696 33408 29745 33436
rect 29696 33396 29702 33408
rect 29733 33405 29745 33408
rect 29779 33405 29791 33439
rect 29733 33399 29791 33405
rect 30006 33396 30012 33448
rect 30064 33436 30070 33448
rect 30101 33439 30159 33445
rect 30101 33436 30113 33439
rect 30064 33408 30113 33436
rect 30064 33396 30070 33408
rect 30101 33405 30113 33408
rect 30147 33405 30159 33439
rect 30101 33399 30159 33405
rect 27074 33371 27132 33377
rect 27074 33368 27086 33371
rect 26169 33340 27086 33368
rect 27074 33337 27086 33340
rect 27120 33337 27132 33371
rect 27074 33331 27132 33337
rect 25547 33272 25921 33300
rect 27801 33303 27859 33309
rect 25547 33269 25559 33272
rect 25501 33263 25559 33269
rect 27801 33269 27813 33303
rect 27847 33300 27859 33303
rect 28442 33300 28448 33312
rect 27847 33272 28448 33300
rect 27847 33269 27859 33272
rect 27801 33263 27859 33269
rect 28442 33260 28448 33272
rect 28500 33260 28506 33312
rect 30285 33303 30343 33309
rect 30285 33269 30297 33303
rect 30331 33300 30343 33303
rect 30650 33300 30656 33312
rect 30331 33272 30656 33300
rect 30331 33269 30343 33272
rect 30285 33263 30343 33269
rect 30650 33260 30656 33272
rect 30708 33260 30714 33312
rect 1104 33210 32016 33232
rect 1104 33158 11253 33210
rect 11305 33158 11317 33210
rect 11369 33158 11381 33210
rect 11433 33158 11445 33210
rect 11497 33158 11509 33210
rect 11561 33158 21557 33210
rect 21609 33158 21621 33210
rect 21673 33158 21685 33210
rect 21737 33158 21749 33210
rect 21801 33158 21813 33210
rect 21865 33158 32016 33210
rect 1104 33136 32016 33158
rect 2038 33096 2044 33108
rect 1596 33068 2044 33096
rect 1596 32960 1624 33068
rect 2038 33056 2044 33068
rect 2096 33056 2102 33108
rect 10413 33099 10471 33105
rect 3979 33068 7696 33096
rect 1670 32988 1676 33040
rect 1728 33028 1734 33040
rect 3979 33028 4007 33068
rect 1728 33000 1900 33028
rect 1728 32988 1734 33000
rect 1872 32969 1900 33000
rect 3344 33000 4007 33028
rect 1765 32963 1823 32969
rect 1765 32960 1777 32963
rect 1596 32932 1777 32960
rect 1765 32929 1777 32932
rect 1811 32929 1823 32963
rect 1765 32923 1823 32929
rect 1857 32963 1915 32969
rect 1857 32929 1869 32963
rect 1903 32929 1915 32963
rect 1857 32923 1915 32929
rect 1949 32963 2007 32969
rect 1949 32929 1961 32963
rect 1995 32929 2007 32963
rect 1949 32923 2007 32929
rect 2133 32963 2191 32969
rect 2133 32929 2145 32963
rect 2179 32960 2191 32963
rect 2222 32960 2228 32972
rect 2179 32932 2228 32960
rect 2179 32929 2191 32932
rect 2133 32923 2191 32929
rect 1489 32759 1547 32765
rect 1489 32725 1501 32759
rect 1535 32756 1547 32759
rect 1670 32756 1676 32768
rect 1535 32728 1676 32756
rect 1535 32725 1547 32728
rect 1489 32719 1547 32725
rect 1670 32716 1676 32728
rect 1728 32716 1734 32768
rect 1872 32756 1900 32923
rect 1964 32824 1992 32923
rect 2222 32920 2228 32932
rect 2280 32920 2286 32972
rect 2866 32960 2872 32972
rect 2827 32932 2872 32960
rect 2866 32920 2872 32932
rect 2924 32920 2930 32972
rect 2038 32852 2044 32904
rect 2096 32892 2102 32904
rect 3145 32895 3203 32901
rect 3145 32892 3157 32895
rect 2096 32864 3157 32892
rect 2096 32852 2102 32864
rect 3145 32861 3157 32864
rect 3191 32861 3203 32895
rect 3145 32855 3203 32861
rect 2130 32824 2136 32836
rect 1964 32796 2136 32824
rect 2130 32784 2136 32796
rect 2188 32824 2194 32836
rect 3344 32833 3372 33000
rect 6730 32988 6736 33040
rect 6788 33028 6794 33040
rect 6788 33000 6960 33028
rect 6788 32988 6794 33000
rect 3510 32960 3516 32972
rect 3471 32932 3516 32960
rect 3510 32920 3516 32932
rect 3568 32920 3574 32972
rect 3878 32960 3884 32972
rect 3839 32932 3884 32960
rect 3878 32920 3884 32932
rect 3936 32920 3942 32972
rect 4617 32963 4675 32969
rect 4617 32929 4629 32963
rect 4663 32960 4675 32963
rect 5353 32963 5411 32969
rect 5353 32960 5365 32963
rect 4663 32932 5365 32960
rect 4663 32929 4675 32932
rect 4617 32923 4675 32929
rect 5353 32929 5365 32932
rect 5399 32960 5411 32963
rect 5534 32960 5540 32972
rect 5399 32932 5540 32960
rect 5399 32929 5411 32932
rect 5353 32923 5411 32929
rect 5534 32920 5540 32932
rect 5592 32960 5598 32972
rect 6457 32963 6515 32969
rect 5592 32932 5764 32960
rect 5592 32920 5598 32932
rect 4890 32892 4896 32904
rect 4851 32864 4896 32892
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 5442 32892 5448 32904
rect 5403 32864 5448 32892
rect 5442 32852 5448 32864
rect 5500 32852 5506 32904
rect 5626 32892 5632 32904
rect 5587 32864 5632 32892
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 3329 32827 3387 32833
rect 2188 32796 3280 32824
rect 2188 32784 2194 32796
rect 3050 32756 3056 32768
rect 1872 32728 3056 32756
rect 3050 32716 3056 32728
rect 3108 32716 3114 32768
rect 3252 32756 3280 32796
rect 3329 32793 3341 32827
rect 3375 32793 3387 32827
rect 3329 32787 3387 32793
rect 3602 32784 3608 32836
rect 3660 32824 3666 32836
rect 3878 32824 3884 32836
rect 3660 32796 3884 32824
rect 3660 32784 3666 32796
rect 3878 32784 3884 32796
rect 3936 32784 3942 32836
rect 4982 32824 4988 32836
rect 4724 32796 4988 32824
rect 3970 32756 3976 32768
rect 3252 32728 3976 32756
rect 3970 32716 3976 32728
rect 4028 32716 4034 32768
rect 4338 32716 4344 32768
rect 4396 32756 4402 32768
rect 4724 32765 4752 32796
rect 4982 32784 4988 32796
rect 5040 32784 5046 32836
rect 5736 32824 5764 32932
rect 6457 32929 6469 32963
rect 6503 32960 6515 32963
rect 6822 32960 6828 32972
rect 6503 32932 6828 32960
rect 6503 32929 6515 32932
rect 6457 32923 6515 32929
rect 6822 32920 6828 32932
rect 6880 32920 6886 32972
rect 6638 32892 6644 32904
rect 6599 32864 6644 32892
rect 6638 32852 6644 32864
rect 6696 32852 6702 32904
rect 6733 32895 6791 32901
rect 6733 32861 6745 32895
rect 6779 32861 6791 32895
rect 6932 32892 6960 33000
rect 7098 32988 7104 33040
rect 7156 32988 7162 33040
rect 7116 32960 7144 32988
rect 7193 32963 7251 32969
rect 7193 32960 7205 32963
rect 7116 32932 7205 32960
rect 7193 32929 7205 32932
rect 7239 32929 7251 32963
rect 7668 32960 7696 33068
rect 10413 33065 10425 33099
rect 10459 33096 10471 33099
rect 10686 33096 10692 33108
rect 10459 33068 10692 33096
rect 10459 33065 10471 33068
rect 10413 33059 10471 33065
rect 10686 33056 10692 33068
rect 10744 33056 10750 33108
rect 11606 33096 11612 33108
rect 11567 33068 11612 33096
rect 11606 33056 11612 33068
rect 11664 33056 11670 33108
rect 11698 33056 11704 33108
rect 11756 33096 11762 33108
rect 12066 33096 12072 33108
rect 11756 33068 12072 33096
rect 11756 33056 11762 33068
rect 12066 33056 12072 33068
rect 12124 33056 12130 33108
rect 13814 33096 13820 33108
rect 12452 33068 13032 33096
rect 13775 33068 13820 33096
rect 7745 33031 7803 33037
rect 7745 32997 7757 33031
rect 7791 33028 7803 33031
rect 8294 33028 8300 33040
rect 7791 33000 8300 33028
rect 7791 32997 7803 33000
rect 7745 32991 7803 32997
rect 8294 32988 8300 33000
rect 8352 32988 8358 33040
rect 9858 33028 9864 33040
rect 8404 33000 9864 33028
rect 8404 32960 8432 33000
rect 9858 32988 9864 33000
rect 9916 32988 9922 33040
rect 9950 32988 9956 33040
rect 10008 33028 10014 33040
rect 10597 33031 10655 33037
rect 10597 33028 10609 33031
rect 10008 33000 10609 33028
rect 10008 32988 10014 33000
rect 10428 32972 10456 33000
rect 10597 32997 10609 33000
rect 10643 33028 10655 33031
rect 12452 33028 12480 33068
rect 10643 33000 12480 33028
rect 10643 32997 10655 33000
rect 10597 32991 10655 32997
rect 12526 32988 12532 33040
rect 12584 33028 12590 33040
rect 13004 33028 13032 33068
rect 13814 33056 13820 33068
rect 13872 33056 13878 33108
rect 15746 33096 15752 33108
rect 13924 33068 15516 33096
rect 15707 33068 15752 33096
rect 13924 33028 13952 33068
rect 15488 33028 15516 33068
rect 15746 33056 15752 33068
rect 15804 33056 15810 33108
rect 17681 33099 17739 33105
rect 17681 33065 17693 33099
rect 17727 33096 17739 33099
rect 18506 33096 18512 33108
rect 17727 33068 18512 33096
rect 17727 33065 17739 33068
rect 17681 33059 17739 33065
rect 18506 33056 18512 33068
rect 18564 33056 18570 33108
rect 22278 33096 22284 33108
rect 18616 33068 22284 33096
rect 16022 33028 16028 33040
rect 12584 33000 12940 33028
rect 13004 33000 13952 33028
rect 14200 33000 15424 33028
rect 15488 33000 16028 33028
rect 12584 32988 12590 33000
rect 7668 32932 8432 32960
rect 8481 32963 8539 32969
rect 7193 32923 7251 32929
rect 8481 32929 8493 32963
rect 8527 32929 8539 32963
rect 9306 32960 9312 32972
rect 9267 32932 9312 32960
rect 8481 32923 8539 32929
rect 8496 32892 8524 32923
rect 9306 32920 9312 32932
rect 9364 32920 9370 32972
rect 10410 32920 10416 32972
rect 10468 32920 10474 32972
rect 10965 32963 11023 32969
rect 10965 32929 10977 32963
rect 11011 32960 11023 32963
rect 11606 32960 11612 32972
rect 11011 32932 11612 32960
rect 11011 32929 11023 32932
rect 10965 32923 11023 32929
rect 11606 32920 11612 32932
rect 11664 32960 11670 32972
rect 12250 32960 12256 32972
rect 11664 32932 12256 32960
rect 11664 32920 11670 32932
rect 12250 32920 12256 32932
rect 12308 32920 12314 32972
rect 12621 32963 12679 32969
rect 12621 32929 12633 32963
rect 12667 32929 12679 32963
rect 12621 32923 12679 32929
rect 8754 32892 8760 32904
rect 6932 32864 8524 32892
rect 8715 32864 8760 32892
rect 6733 32855 6791 32861
rect 6748 32824 6776 32855
rect 8754 32852 8760 32864
rect 8812 32852 8818 32904
rect 9493 32895 9551 32901
rect 9493 32861 9505 32895
rect 9539 32892 9551 32895
rect 9674 32892 9680 32904
rect 9539 32864 9680 32892
rect 9539 32861 9551 32864
rect 9493 32855 9551 32861
rect 9674 32852 9680 32864
rect 9732 32852 9738 32904
rect 5736 32796 6776 32824
rect 6822 32784 6828 32836
rect 6880 32824 6886 32836
rect 7101 32827 7159 32833
rect 7101 32824 7113 32827
rect 6880 32796 7113 32824
rect 6880 32784 6886 32796
rect 7101 32793 7113 32796
rect 7147 32793 7159 32827
rect 7101 32787 7159 32793
rect 8941 32827 8999 32833
rect 8941 32793 8953 32827
rect 8987 32824 8999 32827
rect 12526 32824 12532 32836
rect 8987 32796 12532 32824
rect 8987 32793 8999 32796
rect 8941 32787 8999 32793
rect 12526 32784 12532 32796
rect 12584 32784 12590 32836
rect 12636 32824 12664 32923
rect 12710 32920 12716 32972
rect 12768 32960 12774 32972
rect 12912 32969 12940 33000
rect 12805 32963 12863 32969
rect 12805 32960 12817 32963
rect 12768 32932 12817 32960
rect 12768 32920 12774 32932
rect 12805 32929 12817 32932
rect 12851 32929 12863 32963
rect 12805 32923 12863 32929
rect 12897 32963 12955 32969
rect 12897 32929 12909 32963
rect 12943 32960 12955 32963
rect 13173 32963 13231 32969
rect 12943 32932 13124 32960
rect 12943 32929 12955 32932
rect 12897 32923 12955 32929
rect 12989 32895 13047 32901
rect 12989 32861 13001 32895
rect 13035 32861 13047 32895
rect 13096 32892 13124 32932
rect 13173 32929 13185 32963
rect 13219 32960 13231 32963
rect 13814 32960 13820 32972
rect 13219 32932 13820 32960
rect 13219 32929 13231 32932
rect 13173 32923 13231 32929
rect 13814 32920 13820 32932
rect 13872 32920 13878 32972
rect 14200 32969 14228 33000
rect 15396 32972 15424 33000
rect 16022 32988 16028 33000
rect 16080 32988 16086 33040
rect 17129 33031 17187 33037
rect 17129 32997 17141 33031
rect 17175 33028 17187 33031
rect 17586 33028 17592 33040
rect 17175 33000 17592 33028
rect 17175 32997 17187 33000
rect 17129 32991 17187 32997
rect 17586 32988 17592 33000
rect 17644 32988 17650 33040
rect 18322 32988 18328 33040
rect 18380 33028 18386 33040
rect 18616 33028 18644 33068
rect 22278 33056 22284 33068
rect 22336 33056 22342 33108
rect 22373 33099 22431 33105
rect 22373 33065 22385 33099
rect 22419 33096 22431 33099
rect 22554 33096 22560 33108
rect 22419 33068 22560 33096
rect 22419 33065 22431 33068
rect 22373 33059 22431 33065
rect 22554 33056 22560 33068
rect 22612 33096 22618 33108
rect 22738 33096 22744 33108
rect 22612 33068 22744 33096
rect 22612 33056 22618 33068
rect 22738 33056 22744 33068
rect 22796 33056 22802 33108
rect 23658 33056 23664 33108
rect 23716 33096 23722 33108
rect 24305 33099 24363 33105
rect 24305 33096 24317 33099
rect 23716 33068 24317 33096
rect 23716 33056 23722 33068
rect 24305 33065 24317 33068
rect 24351 33065 24363 33099
rect 24305 33059 24363 33065
rect 24578 33056 24584 33108
rect 24636 33096 24642 33108
rect 24762 33096 24768 33108
rect 24636 33068 24768 33096
rect 24636 33056 24642 33068
rect 24762 33056 24768 33068
rect 24820 33096 24826 33108
rect 24857 33099 24915 33105
rect 24857 33096 24869 33099
rect 24820 33068 24869 33096
rect 24820 33056 24826 33068
rect 24857 33065 24869 33068
rect 24903 33065 24915 33099
rect 24857 33059 24915 33065
rect 25317 33099 25375 33105
rect 25317 33065 25329 33099
rect 25363 33096 25375 33099
rect 25498 33096 25504 33108
rect 25363 33068 25504 33096
rect 25363 33065 25375 33068
rect 25317 33059 25375 33065
rect 25498 33056 25504 33068
rect 25556 33056 25562 33108
rect 25866 33056 25872 33108
rect 25924 33096 25930 33108
rect 26326 33096 26332 33108
rect 25924 33068 26332 33096
rect 25924 33056 25930 33068
rect 26326 33056 26332 33068
rect 26384 33056 26390 33108
rect 26602 33056 26608 33108
rect 26660 33096 26666 33108
rect 30466 33096 30472 33108
rect 26660 33068 30472 33096
rect 26660 33056 26666 33068
rect 30466 33056 30472 33068
rect 30524 33056 30530 33108
rect 18380 33000 18644 33028
rect 18816 33031 18874 33037
rect 18380 32988 18386 33000
rect 18816 32997 18828 33031
rect 18862 33028 18874 33031
rect 19521 33031 19579 33037
rect 19521 33028 19533 33031
rect 18862 33000 19533 33028
rect 18862 32997 18874 33000
rect 18816 32991 18874 32997
rect 19521 32997 19533 33000
rect 19567 32997 19579 33031
rect 19521 32991 19579 32997
rect 19610 32988 19616 33040
rect 19668 33028 19674 33040
rect 21266 33028 21272 33040
rect 19668 33000 21272 33028
rect 19668 32988 19674 33000
rect 21266 32988 21272 33000
rect 21324 32988 21330 33040
rect 24946 33028 24952 33040
rect 22388 33000 24952 33028
rect 14001 32963 14059 32969
rect 14001 32929 14013 32963
rect 14047 32929 14059 32963
rect 14001 32923 14059 32929
rect 14185 32963 14243 32969
rect 14185 32929 14197 32963
rect 14231 32929 14243 32963
rect 14366 32960 14372 32972
rect 14327 32932 14372 32960
rect 14185 32923 14243 32929
rect 13096 32864 13216 32892
rect 12989 32855 13047 32861
rect 12894 32824 12900 32836
rect 12636 32796 12900 32824
rect 12894 32784 12900 32796
rect 12952 32784 12958 32836
rect 13004 32768 13032 32855
rect 13188 32824 13216 32864
rect 13262 32852 13268 32904
rect 13320 32892 13326 32904
rect 14016 32892 14044 32923
rect 14366 32920 14372 32932
rect 14424 32920 14430 32972
rect 14553 32963 14611 32969
rect 14553 32929 14565 32963
rect 14599 32960 14611 32963
rect 15010 32960 15016 32972
rect 14599 32932 15016 32960
rect 14599 32929 14611 32932
rect 14553 32923 14611 32929
rect 15010 32920 15016 32932
rect 15068 32920 15074 32972
rect 15102 32920 15108 32972
rect 15160 32960 15166 32972
rect 15197 32963 15255 32969
rect 15197 32960 15209 32963
rect 15160 32932 15209 32960
rect 15160 32920 15166 32932
rect 15197 32929 15209 32932
rect 15243 32929 15255 32963
rect 15378 32960 15384 32972
rect 15339 32932 15384 32960
rect 15197 32923 15255 32929
rect 15378 32920 15384 32932
rect 15436 32920 15442 32972
rect 15470 32920 15476 32972
rect 15528 32960 15534 32972
rect 15565 32963 15623 32969
rect 15565 32960 15577 32963
rect 15528 32932 15577 32960
rect 15528 32920 15534 32932
rect 15565 32929 15577 32932
rect 15611 32929 15623 32963
rect 15565 32923 15623 32929
rect 15746 32920 15752 32972
rect 15804 32960 15810 32972
rect 16853 32963 16911 32969
rect 16853 32960 16865 32963
rect 15804 32932 16865 32960
rect 15804 32920 15810 32932
rect 16853 32929 16865 32932
rect 16899 32929 16911 32963
rect 17218 32960 17224 32972
rect 17179 32932 17224 32960
rect 16853 32923 16911 32929
rect 17218 32920 17224 32932
rect 17276 32920 17282 32972
rect 18506 32920 18512 32972
rect 18564 32960 18570 32972
rect 19334 32960 19340 32972
rect 18564 32932 19340 32960
rect 18564 32920 18570 32932
rect 19334 32920 19340 32932
rect 19392 32960 19398 32972
rect 19702 32960 19708 32972
rect 19392 32932 19708 32960
rect 19392 32920 19398 32932
rect 19702 32920 19708 32932
rect 19760 32920 19766 32972
rect 19794 32920 19800 32972
rect 19852 32970 19858 32972
rect 19852 32963 19923 32970
rect 19852 32929 19855 32963
rect 19889 32932 19923 32963
rect 20073 32963 20131 32969
rect 19889 32929 19901 32932
rect 19852 32923 19901 32929
rect 20073 32929 20085 32963
rect 20119 32929 20131 32963
rect 20073 32923 20131 32929
rect 19852 32920 19858 32923
rect 13320 32864 14044 32892
rect 13320 32852 13326 32864
rect 14016 32824 14044 32864
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32892 14335 32895
rect 15289 32895 15347 32901
rect 15289 32892 15301 32895
rect 14323 32864 15301 32892
rect 14323 32861 14335 32864
rect 14277 32855 14335 32861
rect 15289 32861 15301 32864
rect 15335 32892 15347 32895
rect 15654 32892 15660 32904
rect 15335 32864 15660 32892
rect 15335 32861 15347 32864
rect 15289 32855 15347 32861
rect 15654 32852 15660 32864
rect 15712 32852 15718 32904
rect 16206 32852 16212 32904
rect 16264 32892 16270 32904
rect 16669 32895 16727 32901
rect 16669 32892 16681 32895
rect 16264 32864 16681 32892
rect 16264 32852 16270 32864
rect 16669 32861 16681 32864
rect 16715 32861 16727 32895
rect 16669 32855 16727 32861
rect 19061 32895 19119 32901
rect 19061 32861 19073 32895
rect 19107 32861 19119 32895
rect 19061 32855 19119 32861
rect 14458 32824 14464 32836
rect 13188 32796 13492 32824
rect 14016 32796 14464 32824
rect 4709 32759 4767 32765
rect 4709 32756 4721 32759
rect 4396 32728 4721 32756
rect 4396 32716 4402 32728
rect 4709 32725 4721 32728
rect 4755 32725 4767 32759
rect 4709 32719 4767 32725
rect 4801 32759 4859 32765
rect 4801 32725 4813 32759
rect 4847 32756 4859 32759
rect 5350 32756 5356 32768
rect 4847 32728 5356 32756
rect 4847 32725 4859 32728
rect 4801 32719 4859 32725
rect 5350 32716 5356 32728
rect 5408 32716 5414 32768
rect 5537 32759 5595 32765
rect 5537 32725 5549 32759
rect 5583 32756 5595 32759
rect 5994 32756 6000 32768
rect 5583 32728 6000 32756
rect 5583 32725 5595 32728
rect 5537 32719 5595 32725
rect 5994 32716 6000 32728
rect 6052 32716 6058 32768
rect 6638 32716 6644 32768
rect 6696 32756 6702 32768
rect 8110 32756 8116 32768
rect 6696 32728 8116 32756
rect 6696 32716 6702 32728
rect 8110 32716 8116 32728
rect 8168 32716 8174 32768
rect 8294 32716 8300 32768
rect 8352 32756 8358 32768
rect 9398 32756 9404 32768
rect 8352 32728 9404 32756
rect 8352 32716 8358 32728
rect 9398 32716 9404 32728
rect 9456 32716 9462 32768
rect 10597 32759 10655 32765
rect 10597 32725 10609 32759
rect 10643 32756 10655 32759
rect 10778 32756 10784 32768
rect 10643 32728 10784 32756
rect 10643 32725 10655 32728
rect 10597 32719 10655 32725
rect 10778 32716 10784 32728
rect 10836 32756 10842 32768
rect 11146 32756 11152 32768
rect 10836 32728 11152 32756
rect 10836 32716 10842 32728
rect 11146 32716 11152 32728
rect 11204 32716 11210 32768
rect 12161 32759 12219 32765
rect 12161 32725 12173 32759
rect 12207 32756 12219 32759
rect 12986 32756 12992 32768
rect 12207 32728 12992 32756
rect 12207 32725 12219 32728
rect 12161 32719 12219 32725
rect 12986 32716 12992 32728
rect 13044 32716 13050 32768
rect 13354 32756 13360 32768
rect 13315 32728 13360 32756
rect 13354 32716 13360 32728
rect 13412 32716 13418 32768
rect 13464 32756 13492 32796
rect 14458 32784 14464 32796
rect 14516 32824 14522 32836
rect 15194 32824 15200 32836
rect 14516 32796 15200 32824
rect 14516 32784 14522 32796
rect 15194 32784 15200 32796
rect 15252 32784 15258 32836
rect 19076 32824 19104 32855
rect 19150 32852 19156 32904
rect 19208 32892 19214 32904
rect 19426 32892 19432 32904
rect 19208 32864 19432 32892
rect 19208 32852 19214 32864
rect 19426 32852 19432 32864
rect 19484 32892 19490 32904
rect 19981 32895 20039 32901
rect 19981 32892 19993 32895
rect 19484 32864 19993 32892
rect 19484 32852 19490 32864
rect 19981 32861 19993 32864
rect 20027 32861 20039 32895
rect 19981 32855 20039 32861
rect 19242 32824 19248 32836
rect 19076 32796 19248 32824
rect 17402 32756 17408 32768
rect 13464 32728 17408 32756
rect 17402 32716 17408 32728
rect 17460 32716 17466 32768
rect 17954 32716 17960 32768
rect 18012 32756 18018 32768
rect 19076 32756 19104 32796
rect 19242 32784 19248 32796
rect 19300 32784 19306 32836
rect 18012 32728 19104 32756
rect 18012 32716 18018 32728
rect 19150 32716 19156 32768
rect 19208 32756 19214 32768
rect 19610 32756 19616 32768
rect 19208 32728 19616 32756
rect 19208 32716 19214 32728
rect 19610 32716 19616 32728
rect 19668 32716 19674 32768
rect 19978 32716 19984 32768
rect 20036 32756 20042 32768
rect 20088 32756 20116 32923
rect 20162 32920 20168 32972
rect 20220 32960 20226 32972
rect 20257 32963 20315 32969
rect 20257 32960 20269 32963
rect 20220 32932 20269 32960
rect 20220 32920 20226 32932
rect 20257 32929 20269 32932
rect 20303 32960 20315 32963
rect 20530 32960 20536 32972
rect 20303 32932 20536 32960
rect 20303 32929 20315 32932
rect 20257 32923 20315 32929
rect 20530 32920 20536 32932
rect 20588 32920 20594 32972
rect 20714 32960 20720 32972
rect 20675 32932 20720 32960
rect 20714 32920 20720 32932
rect 20772 32920 20778 32972
rect 20898 32960 20904 32972
rect 20859 32932 20904 32960
rect 20898 32920 20904 32932
rect 20956 32920 20962 32972
rect 22186 32960 22192 32972
rect 22147 32932 22192 32960
rect 22186 32920 22192 32932
rect 22244 32920 22250 32972
rect 20438 32784 20444 32836
rect 20496 32824 20502 32836
rect 21177 32827 21235 32833
rect 20496 32796 20944 32824
rect 20496 32784 20502 32796
rect 20036 32728 20116 32756
rect 20036 32716 20042 32728
rect 20162 32716 20168 32768
rect 20220 32756 20226 32768
rect 20806 32756 20812 32768
rect 20220 32728 20812 32756
rect 20220 32716 20226 32728
rect 20806 32716 20812 32728
rect 20864 32716 20870 32768
rect 20916 32756 20944 32796
rect 21177 32793 21189 32827
rect 21223 32824 21235 32827
rect 22388 32824 22416 33000
rect 24946 32988 24952 33000
rect 25004 32988 25010 33040
rect 25038 32988 25044 33040
rect 25096 33028 25102 33040
rect 26050 33028 26056 33040
rect 25096 33000 26056 33028
rect 25096 32988 25102 33000
rect 26050 32988 26056 33000
rect 26108 33028 26114 33040
rect 26108 33000 27200 33028
rect 26108 32988 26114 33000
rect 22462 32920 22468 32972
rect 22520 32960 22526 32972
rect 22925 32963 22983 32969
rect 22925 32960 22937 32963
rect 22520 32932 22937 32960
rect 22520 32920 22526 32932
rect 22925 32929 22937 32932
rect 22971 32929 22983 32963
rect 22925 32923 22983 32929
rect 23192 32963 23250 32969
rect 23192 32929 23204 32963
rect 23238 32960 23250 32963
rect 23566 32960 23572 32972
rect 23238 32932 23572 32960
rect 23238 32929 23250 32932
rect 23192 32923 23250 32929
rect 23566 32920 23572 32932
rect 23624 32920 23630 32972
rect 24854 32920 24860 32972
rect 24912 32960 24918 32972
rect 25409 32963 25467 32969
rect 25409 32960 25421 32963
rect 24912 32932 25421 32960
rect 24912 32920 24918 32932
rect 25409 32929 25421 32932
rect 25455 32929 25467 32963
rect 25590 32960 25596 32972
rect 25551 32932 25596 32960
rect 25409 32923 25467 32929
rect 25590 32920 25596 32932
rect 25648 32920 25654 32972
rect 25774 32960 25780 32972
rect 25735 32932 25780 32960
rect 25774 32920 25780 32932
rect 25832 32920 25838 32972
rect 25961 32963 26019 32969
rect 25961 32929 25973 32963
rect 26007 32929 26019 32963
rect 26142 32960 26148 32972
rect 26103 32932 26148 32960
rect 25961 32923 26019 32929
rect 24946 32852 24952 32904
rect 25004 32892 25010 32904
rect 25317 32895 25375 32901
rect 25317 32892 25329 32895
rect 25004 32864 25329 32892
rect 25004 32852 25010 32864
rect 25317 32861 25329 32864
rect 25363 32861 25375 32895
rect 25317 32855 25375 32861
rect 25685 32895 25743 32901
rect 25685 32861 25697 32895
rect 25731 32892 25743 32895
rect 25866 32892 25872 32904
rect 25731 32864 25872 32892
rect 25731 32861 25743 32864
rect 25685 32855 25743 32861
rect 25866 32852 25872 32864
rect 25924 32852 25930 32904
rect 25976 32892 26004 32923
rect 26142 32920 26148 32932
rect 26200 32920 26206 32972
rect 27172 32969 27200 33000
rect 28350 32988 28356 33040
rect 28408 32988 28414 33040
rect 28626 32988 28632 33040
rect 28684 33028 28690 33040
rect 28684 33000 30144 33028
rect 28684 32988 28690 33000
rect 27157 32963 27215 32969
rect 27157 32929 27169 32963
rect 27203 32929 27215 32963
rect 27157 32923 27215 32929
rect 28077 32963 28135 32969
rect 28077 32929 28089 32963
rect 28123 32960 28135 32963
rect 28166 32960 28172 32972
rect 28123 32932 28172 32960
rect 28123 32929 28135 32932
rect 28077 32923 28135 32929
rect 28166 32920 28172 32932
rect 28224 32920 28230 32972
rect 28368 32960 28396 32988
rect 28810 32960 28816 32972
rect 28368 32932 28816 32960
rect 28810 32920 28816 32932
rect 28868 32960 28874 32972
rect 29549 32963 29607 32969
rect 29549 32960 29561 32963
rect 28868 32932 29561 32960
rect 28868 32920 28874 32932
rect 29549 32929 29561 32932
rect 29595 32929 29607 32963
rect 29730 32960 29736 32972
rect 29691 32932 29736 32960
rect 29549 32923 29607 32929
rect 29730 32920 29736 32932
rect 29788 32920 29794 32972
rect 29914 32960 29920 32972
rect 29875 32932 29920 32960
rect 29914 32920 29920 32932
rect 29972 32920 29978 32972
rect 30116 32969 30144 33000
rect 30101 32963 30159 32969
rect 30101 32929 30113 32963
rect 30147 32929 30159 32963
rect 30101 32923 30159 32929
rect 26050 32892 26056 32904
rect 25976 32864 26056 32892
rect 26050 32852 26056 32864
rect 26108 32892 26114 32904
rect 27341 32895 27399 32901
rect 27341 32892 27353 32895
rect 26108 32864 27353 32892
rect 26108 32852 26114 32864
rect 27341 32861 27353 32864
rect 27387 32861 27399 32895
rect 27341 32855 27399 32861
rect 28353 32895 28411 32901
rect 28353 32861 28365 32895
rect 28399 32892 28411 32895
rect 28626 32892 28632 32904
rect 28399 32864 28632 32892
rect 28399 32861 28411 32864
rect 28353 32855 28411 32861
rect 28626 32852 28632 32864
rect 28684 32852 28690 32904
rect 29822 32852 29828 32904
rect 29880 32892 29886 32904
rect 29880 32864 29925 32892
rect 29880 32852 29886 32864
rect 21223 32796 22416 32824
rect 21223 32793 21235 32796
rect 21177 32787 21235 32793
rect 23934 32784 23940 32836
rect 23992 32824 23998 32836
rect 26973 32827 27031 32833
rect 26973 32824 26985 32827
rect 23992 32796 26985 32824
rect 23992 32784 23998 32796
rect 26973 32793 26985 32796
rect 27019 32793 27031 32827
rect 26973 32787 27031 32793
rect 28994 32784 29000 32836
rect 29052 32824 29058 32836
rect 31113 32827 31171 32833
rect 31113 32824 31125 32827
rect 29052 32796 31125 32824
rect 29052 32784 29058 32796
rect 31113 32793 31125 32796
rect 31159 32793 31171 32827
rect 31113 32787 31171 32793
rect 21910 32756 21916 32768
rect 20916 32728 21916 32756
rect 21910 32716 21916 32728
rect 21968 32716 21974 32768
rect 22094 32716 22100 32768
rect 22152 32756 22158 32768
rect 27614 32756 27620 32768
rect 22152 32728 27620 32756
rect 22152 32716 22158 32728
rect 27614 32716 27620 32728
rect 27672 32716 27678 32768
rect 29362 32756 29368 32768
rect 29323 32728 29368 32756
rect 29362 32716 29368 32728
rect 29420 32716 29426 32768
rect 29822 32716 29828 32768
rect 29880 32756 29886 32768
rect 30561 32759 30619 32765
rect 30561 32756 30573 32759
rect 29880 32728 30573 32756
rect 29880 32716 29886 32728
rect 30561 32725 30573 32728
rect 30607 32725 30619 32759
rect 30561 32719 30619 32725
rect 1104 32666 32016 32688
rect 1104 32614 6102 32666
rect 6154 32614 6166 32666
rect 6218 32614 6230 32666
rect 6282 32614 6294 32666
rect 6346 32614 6358 32666
rect 6410 32614 16405 32666
rect 16457 32614 16469 32666
rect 16521 32614 16533 32666
rect 16585 32614 16597 32666
rect 16649 32614 16661 32666
rect 16713 32614 26709 32666
rect 26761 32614 26773 32666
rect 26825 32614 26837 32666
rect 26889 32614 26901 32666
rect 26953 32614 26965 32666
rect 27017 32614 32016 32666
rect 1104 32592 32016 32614
rect 1765 32555 1823 32561
rect 1765 32521 1777 32555
rect 1811 32552 1823 32555
rect 2038 32552 2044 32564
rect 1811 32524 2044 32552
rect 1811 32521 1823 32524
rect 1765 32515 1823 32521
rect 2038 32512 2044 32524
rect 2096 32512 2102 32564
rect 2498 32552 2504 32564
rect 2332 32524 2504 32552
rect 2222 32484 2228 32496
rect 1780 32456 2228 32484
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 1780 32348 1808 32456
rect 2222 32444 2228 32456
rect 2280 32444 2286 32496
rect 1857 32419 1915 32425
rect 1857 32385 1869 32419
rect 1903 32416 1915 32419
rect 2038 32416 2044 32428
rect 1903 32388 2044 32416
rect 1903 32385 1915 32388
rect 1857 32379 1915 32385
rect 2038 32376 2044 32388
rect 2096 32376 2102 32428
rect 2332 32416 2360 32524
rect 2498 32512 2504 32524
rect 2556 32512 2562 32564
rect 3326 32512 3332 32564
rect 3384 32552 3390 32564
rect 3789 32555 3847 32561
rect 3789 32552 3801 32555
rect 3384 32524 3801 32552
rect 3384 32512 3390 32524
rect 3789 32521 3801 32524
rect 3835 32521 3847 32555
rect 3789 32515 3847 32521
rect 4890 32512 4896 32564
rect 4948 32552 4954 32564
rect 5166 32552 5172 32564
rect 4948 32524 5172 32552
rect 4948 32512 4954 32524
rect 5166 32512 5172 32524
rect 5224 32512 5230 32564
rect 6730 32552 6736 32564
rect 5506 32524 6736 32552
rect 2406 32444 2412 32496
rect 2464 32484 2470 32496
rect 3145 32487 3203 32493
rect 2464 32456 2820 32484
rect 2464 32444 2470 32456
rect 2792 32425 2820 32456
rect 3145 32453 3157 32487
rect 3191 32484 3203 32487
rect 3510 32484 3516 32496
rect 3191 32456 3516 32484
rect 3191 32453 3203 32456
rect 3145 32447 3203 32453
rect 3510 32444 3516 32456
rect 3568 32444 3574 32496
rect 4525 32487 4583 32493
rect 4525 32453 4537 32487
rect 4571 32484 4583 32487
rect 5258 32484 5264 32496
rect 4571 32456 5264 32484
rect 4571 32453 4583 32456
rect 4525 32447 4583 32453
rect 5258 32444 5264 32456
rect 5316 32444 5322 32496
rect 2501 32419 2559 32425
rect 2501 32416 2513 32419
rect 2332 32388 2513 32416
rect 2501 32385 2513 32388
rect 2547 32385 2559 32419
rect 2501 32379 2559 32385
rect 2777 32419 2835 32425
rect 2777 32385 2789 32419
rect 2823 32385 2835 32419
rect 3234 32416 3240 32428
rect 3195 32388 3240 32416
rect 2777 32379 2835 32385
rect 3234 32376 3240 32388
rect 3292 32376 3298 32428
rect 3326 32376 3332 32428
rect 3384 32416 3390 32428
rect 5506 32416 5534 32524
rect 6730 32512 6736 32524
rect 6788 32512 6794 32564
rect 7650 32512 7656 32564
rect 7708 32552 7714 32564
rect 7745 32555 7803 32561
rect 7745 32552 7757 32555
rect 7708 32524 7757 32552
rect 7708 32512 7714 32524
rect 7745 32521 7757 32524
rect 7791 32521 7803 32555
rect 9122 32552 9128 32564
rect 9083 32524 9128 32552
rect 7745 32515 7803 32521
rect 9122 32512 9128 32524
rect 9180 32512 9186 32564
rect 9674 32552 9680 32564
rect 9635 32524 9680 32552
rect 9674 32512 9680 32524
rect 9732 32512 9738 32564
rect 14090 32552 14096 32564
rect 11808 32524 14096 32552
rect 6454 32444 6460 32496
rect 6512 32484 6518 32496
rect 6549 32487 6607 32493
rect 6549 32484 6561 32487
rect 6512 32456 6561 32484
rect 6512 32444 6518 32456
rect 6549 32453 6561 32456
rect 6595 32453 6607 32487
rect 6549 32447 6607 32453
rect 7374 32444 7380 32496
rect 7432 32484 7438 32496
rect 8110 32484 8116 32496
rect 7432 32456 8116 32484
rect 7432 32444 7438 32456
rect 8110 32444 8116 32456
rect 8168 32484 8174 32496
rect 8168 32456 8616 32484
rect 8168 32444 8174 32456
rect 3384 32388 5534 32416
rect 3384 32376 3390 32388
rect 5994 32376 6000 32428
rect 6052 32416 6058 32428
rect 6365 32419 6423 32425
rect 6365 32416 6377 32419
rect 6052 32388 6377 32416
rect 6052 32376 6058 32388
rect 6365 32385 6377 32388
rect 6411 32385 6423 32419
rect 6365 32379 6423 32385
rect 1688 32320 1808 32348
rect 1949 32351 2007 32357
rect 1688 32292 1716 32320
rect 1949 32317 1961 32351
rect 1995 32317 2007 32351
rect 1949 32311 2007 32317
rect 1670 32240 1676 32292
rect 1728 32240 1734 32292
rect 1964 32212 1992 32311
rect 2590 32308 2596 32360
rect 2648 32348 2654 32360
rect 2685 32351 2743 32357
rect 2685 32348 2697 32351
rect 2648 32320 2697 32348
rect 2648 32308 2654 32320
rect 2685 32317 2697 32320
rect 2731 32348 2743 32351
rect 2731 32320 3112 32348
rect 2731 32317 2743 32320
rect 2685 32311 2743 32317
rect 2222 32212 2228 32224
rect 1964 32184 2228 32212
rect 2222 32172 2228 32184
rect 2280 32212 2286 32224
rect 2774 32212 2780 32224
rect 2280 32184 2780 32212
rect 2280 32172 2286 32184
rect 2774 32172 2780 32184
rect 2832 32172 2838 32224
rect 3084 32212 3112 32320
rect 3142 32308 3148 32360
rect 3200 32348 3206 32360
rect 3789 32351 3847 32357
rect 3789 32348 3801 32351
rect 3200 32320 3801 32348
rect 3200 32308 3206 32320
rect 3789 32317 3801 32320
rect 3835 32317 3847 32351
rect 3970 32348 3976 32360
rect 3931 32320 3976 32348
rect 3789 32311 3847 32317
rect 3970 32308 3976 32320
rect 4028 32308 4034 32360
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32317 4491 32351
rect 4433 32311 4491 32317
rect 3602 32240 3608 32292
rect 3660 32280 3666 32292
rect 4448 32280 4476 32311
rect 4522 32308 4528 32360
rect 4580 32348 4586 32360
rect 5077 32351 5135 32357
rect 5077 32348 5089 32351
rect 4580 32320 5089 32348
rect 4580 32308 4586 32320
rect 5077 32317 5089 32320
rect 5123 32317 5135 32351
rect 5077 32311 5135 32317
rect 5350 32308 5356 32360
rect 5408 32348 5414 32360
rect 6089 32351 6147 32357
rect 6089 32348 6101 32351
rect 5408 32320 6101 32348
rect 5408 32308 5414 32320
rect 6089 32317 6101 32320
rect 6135 32317 6147 32351
rect 6822 32348 6828 32360
rect 6783 32320 6828 32348
rect 6089 32311 6147 32317
rect 6822 32308 6828 32320
rect 6880 32308 6886 32360
rect 7190 32348 7196 32360
rect 7151 32320 7196 32348
rect 7190 32308 7196 32320
rect 7248 32308 7254 32360
rect 8018 32348 8024 32360
rect 7979 32320 8024 32348
rect 8018 32308 8024 32320
rect 8076 32308 8082 32360
rect 8113 32351 8171 32357
rect 8113 32317 8125 32351
rect 8159 32317 8171 32351
rect 8113 32311 8171 32317
rect 8226 32348 8284 32354
rect 8226 32314 8238 32348
rect 8272 32345 8284 32348
rect 8312 32345 8340 32456
rect 8272 32317 8340 32345
rect 8389 32351 8447 32357
rect 8389 32317 8401 32351
rect 8435 32317 8447 32351
rect 8588 32348 8616 32456
rect 8662 32444 8668 32496
rect 8720 32484 8726 32496
rect 10502 32484 10508 32496
rect 8720 32456 9168 32484
rect 8720 32444 8726 32456
rect 9140 32357 9168 32456
rect 9646 32456 10508 32484
rect 9646 32416 9674 32456
rect 10502 32444 10508 32456
rect 10560 32444 10566 32496
rect 11054 32444 11060 32496
rect 11112 32444 11118 32496
rect 10962 32416 10968 32428
rect 9232 32388 9674 32416
rect 10923 32388 10968 32416
rect 9232 32360 9260 32388
rect 10962 32376 10968 32388
rect 11020 32376 11026 32428
rect 11072 32416 11100 32444
rect 11808 32425 11836 32524
rect 14090 32512 14096 32524
rect 14148 32512 14154 32564
rect 14550 32552 14556 32564
rect 14511 32524 14556 32552
rect 14550 32512 14556 32524
rect 14608 32512 14614 32564
rect 14918 32512 14924 32564
rect 14976 32552 14982 32564
rect 15102 32552 15108 32564
rect 14976 32524 15108 32552
rect 14976 32512 14982 32524
rect 15102 32512 15108 32524
rect 15160 32552 15166 32564
rect 15565 32555 15623 32561
rect 15565 32552 15577 32555
rect 15160 32524 15577 32552
rect 15160 32512 15166 32524
rect 15565 32521 15577 32524
rect 15611 32552 15623 32555
rect 15611 32524 15985 32552
rect 15611 32521 15623 32524
rect 15565 32515 15623 32521
rect 12894 32444 12900 32496
rect 12952 32484 12958 32496
rect 13173 32487 13231 32493
rect 13173 32484 13185 32487
rect 12952 32456 13185 32484
rect 12952 32444 12958 32456
rect 13173 32453 13185 32456
rect 13219 32453 13231 32487
rect 13173 32447 13231 32453
rect 15197 32487 15255 32493
rect 15197 32453 15209 32487
rect 15243 32484 15255 32487
rect 15470 32484 15476 32496
rect 15243 32456 15476 32484
rect 15243 32453 15255 32456
rect 15197 32447 15255 32453
rect 15470 32444 15476 32456
rect 15528 32444 15534 32496
rect 15746 32444 15752 32496
rect 15804 32484 15810 32496
rect 15957 32484 15985 32524
rect 16022 32512 16028 32564
rect 16080 32552 16086 32564
rect 17218 32552 17224 32564
rect 16080 32524 17224 32552
rect 16080 32512 16086 32524
rect 17218 32512 17224 32524
rect 17276 32512 17282 32564
rect 17402 32512 17408 32564
rect 17460 32552 17466 32564
rect 18966 32552 18972 32564
rect 17460 32524 18972 32552
rect 17460 32512 17466 32524
rect 18966 32512 18972 32524
rect 19024 32512 19030 32564
rect 19702 32512 19708 32564
rect 19760 32552 19766 32564
rect 21361 32555 21419 32561
rect 19760 32524 20760 32552
rect 19760 32512 19766 32524
rect 16298 32484 16304 32496
rect 15804 32456 15849 32484
rect 15957 32456 16304 32484
rect 15804 32444 15810 32456
rect 16298 32444 16304 32456
rect 16356 32444 16362 32496
rect 16574 32444 16580 32496
rect 16632 32484 16638 32496
rect 16632 32456 17724 32484
rect 16632 32444 16638 32456
rect 11793 32419 11851 32425
rect 11793 32416 11805 32419
rect 11072 32388 11805 32416
rect 11793 32385 11805 32388
rect 11839 32385 11851 32419
rect 11793 32379 11851 32385
rect 13354 32376 13360 32428
rect 13412 32416 13418 32428
rect 14093 32419 14151 32425
rect 14093 32416 14105 32419
rect 13412 32388 14105 32416
rect 13412 32376 13418 32388
rect 14093 32385 14105 32388
rect 14139 32385 14151 32419
rect 15488 32416 15516 32444
rect 17310 32416 17316 32428
rect 15488 32388 17316 32416
rect 14093 32379 14151 32385
rect 8941 32351 8999 32357
rect 8941 32348 8953 32351
rect 8588 32320 8953 32348
rect 8272 32314 8284 32317
rect 3660 32252 4476 32280
rect 3660 32240 3666 32252
rect 5534 32240 5540 32292
rect 5592 32280 5598 32292
rect 5994 32280 6000 32292
rect 5592 32252 6000 32280
rect 5592 32240 5598 32252
rect 5994 32240 6000 32252
rect 6052 32240 6058 32292
rect 6914 32240 6920 32292
rect 6972 32280 6978 32292
rect 6972 32252 7328 32280
rect 6972 32240 6978 32252
rect 4338 32212 4344 32224
rect 3084 32184 4344 32212
rect 4338 32172 4344 32184
rect 4396 32172 4402 32224
rect 5166 32212 5172 32224
rect 5127 32184 5172 32212
rect 5166 32172 5172 32184
rect 5224 32172 5230 32224
rect 7190 32172 7196 32224
rect 7248 32212 7254 32224
rect 7300 32212 7328 32252
rect 7374 32240 7380 32292
rect 7432 32280 7438 32292
rect 8125 32280 8153 32311
rect 8226 32308 8284 32314
rect 8389 32311 8447 32317
rect 8941 32317 8953 32320
rect 8987 32317 8999 32351
rect 8941 32311 8999 32317
rect 9125 32351 9183 32357
rect 9125 32317 9137 32351
rect 9171 32317 9183 32351
rect 9125 32311 9183 32317
rect 8404 32280 8432 32311
rect 9214 32308 9220 32360
rect 9272 32308 9278 32360
rect 9582 32348 9588 32360
rect 9543 32320 9588 32348
rect 9582 32308 9588 32320
rect 9640 32308 9646 32360
rect 10778 32348 10784 32360
rect 10739 32320 10784 32348
rect 10778 32308 10784 32320
rect 10836 32308 10842 32360
rect 10870 32308 10876 32360
rect 10928 32348 10934 32360
rect 11057 32351 11115 32357
rect 11057 32348 11069 32351
rect 10928 32320 11069 32348
rect 10928 32308 10934 32320
rect 11057 32317 11069 32320
rect 11103 32317 11115 32351
rect 11057 32311 11115 32317
rect 11146 32308 11152 32360
rect 11204 32348 11210 32360
rect 11333 32351 11391 32357
rect 11204 32320 11249 32348
rect 11204 32308 11210 32320
rect 11333 32317 11345 32351
rect 11379 32348 11391 32351
rect 12618 32348 12624 32360
rect 11379 32320 12624 32348
rect 11379 32317 11391 32320
rect 11333 32311 11391 32317
rect 12618 32308 12624 32320
rect 12676 32308 12682 32360
rect 14274 32348 14280 32360
rect 14235 32320 14280 32348
rect 14274 32308 14280 32320
rect 14332 32308 14338 32360
rect 14826 32308 14832 32360
rect 14884 32348 14890 32360
rect 16022 32348 16028 32360
rect 14884 32320 16028 32348
rect 14884 32308 14890 32320
rect 16022 32308 16028 32320
rect 16080 32308 16086 32360
rect 16206 32348 16212 32360
rect 16167 32320 16212 32348
rect 16206 32308 16212 32320
rect 16264 32308 16270 32360
rect 16298 32308 16304 32360
rect 16356 32348 16362 32360
rect 16393 32351 16451 32357
rect 16393 32348 16405 32351
rect 16356 32320 16405 32348
rect 16356 32308 16362 32320
rect 16393 32317 16405 32320
rect 16439 32317 16451 32351
rect 16574 32348 16580 32360
rect 16535 32320 16580 32348
rect 16393 32311 16451 32317
rect 16574 32308 16580 32320
rect 16632 32308 16638 32360
rect 16669 32351 16727 32357
rect 16669 32317 16681 32351
rect 16715 32317 16727 32351
rect 16669 32311 16727 32317
rect 7432 32252 8153 32280
rect 7432 32240 7438 32252
rect 8018 32212 8024 32224
rect 7248 32184 8024 32212
rect 7248 32172 7254 32184
rect 8018 32172 8024 32184
rect 8076 32172 8082 32224
rect 8125 32212 8153 32252
rect 8312 32252 8432 32280
rect 8312 32224 8340 32252
rect 9858 32240 9864 32292
rect 9916 32280 9922 32292
rect 9916 32252 11836 32280
rect 9916 32240 9922 32252
rect 8202 32212 8208 32224
rect 8125 32184 8208 32212
rect 8202 32172 8208 32184
rect 8260 32172 8266 32224
rect 8294 32172 8300 32224
rect 8352 32172 8358 32224
rect 10594 32212 10600 32224
rect 10555 32184 10600 32212
rect 10594 32172 10600 32184
rect 10652 32172 10658 32224
rect 11808 32212 11836 32252
rect 11882 32240 11888 32292
rect 11940 32280 11946 32292
rect 12038 32283 12096 32289
rect 12038 32280 12050 32283
rect 11940 32252 12050 32280
rect 11940 32240 11946 32252
rect 12038 32249 12050 32252
rect 12084 32249 12096 32283
rect 12038 32243 12096 32249
rect 14645 32283 14703 32289
rect 14645 32249 14657 32283
rect 14691 32280 14703 32283
rect 15286 32280 15292 32292
rect 14691 32252 15292 32280
rect 14691 32249 14703 32252
rect 14645 32243 14703 32249
rect 15286 32240 15292 32252
rect 15344 32240 15350 32292
rect 16482 32280 16488 32292
rect 15488 32252 16488 32280
rect 15488 32212 15516 32252
rect 16482 32240 16488 32252
rect 16540 32240 16546 32292
rect 16684 32280 16712 32311
rect 16758 32308 16764 32360
rect 16816 32348 16822 32360
rect 16960 32357 16988 32388
rect 17310 32376 17316 32388
rect 17368 32376 17374 32428
rect 17696 32416 17724 32456
rect 18046 32444 18052 32496
rect 18104 32484 18110 32496
rect 20162 32484 20168 32496
rect 18104 32456 20168 32484
rect 18104 32444 18110 32456
rect 20162 32444 20168 32456
rect 20220 32444 20226 32496
rect 20622 32484 20628 32496
rect 20272 32456 20628 32484
rect 18325 32419 18383 32425
rect 18325 32416 18337 32419
rect 17696 32388 18337 32416
rect 18325 32385 18337 32388
rect 18371 32416 18383 32419
rect 19061 32419 19119 32425
rect 19061 32416 19073 32419
rect 18371 32388 19073 32416
rect 18371 32385 18383 32388
rect 18325 32379 18383 32385
rect 19061 32385 19073 32388
rect 19107 32385 19119 32419
rect 20070 32416 20076 32428
rect 19061 32379 19119 32385
rect 19628 32388 20076 32416
rect 16945 32351 17003 32357
rect 16816 32320 16861 32348
rect 16816 32308 16822 32320
rect 16945 32317 16957 32351
rect 16991 32317 17003 32351
rect 16945 32311 17003 32317
rect 17218 32308 17224 32360
rect 17276 32348 17282 32360
rect 19628 32348 19656 32388
rect 20070 32376 20076 32388
rect 20128 32376 20134 32428
rect 17276 32320 19656 32348
rect 17276 32308 17282 32320
rect 19702 32308 19708 32360
rect 19760 32348 19766 32360
rect 20165 32351 20223 32357
rect 19760 32320 19805 32348
rect 19760 32308 19766 32320
rect 20165 32317 20177 32351
rect 20211 32348 20223 32351
rect 20272 32348 20300 32456
rect 20622 32444 20628 32456
rect 20680 32444 20686 32496
rect 20438 32416 20444 32428
rect 20399 32388 20444 32416
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 20732 32357 20760 32524
rect 21361 32521 21373 32555
rect 21407 32552 21419 32555
rect 22094 32552 22100 32564
rect 21407 32524 22100 32552
rect 21407 32521 21419 32524
rect 21361 32515 21419 32521
rect 22094 32512 22100 32524
rect 22152 32512 22158 32564
rect 22186 32512 22192 32564
rect 22244 32552 22250 32564
rect 22649 32555 22707 32561
rect 22649 32552 22661 32555
rect 22244 32524 22661 32552
rect 22244 32512 22250 32524
rect 22649 32521 22661 32524
rect 22695 32521 22707 32555
rect 23566 32552 23572 32564
rect 23527 32524 23572 32552
rect 22649 32515 22707 32521
rect 23566 32512 23572 32524
rect 23624 32512 23630 32564
rect 24857 32555 24915 32561
rect 24857 32521 24869 32555
rect 24903 32552 24915 32555
rect 26602 32552 26608 32564
rect 24903 32524 26608 32552
rect 24903 32521 24915 32524
rect 24857 32515 24915 32521
rect 26602 32512 26608 32524
rect 26660 32512 26666 32564
rect 27341 32555 27399 32561
rect 27341 32521 27353 32555
rect 27387 32552 27399 32555
rect 27982 32552 27988 32564
rect 27387 32524 27988 32552
rect 27387 32521 27399 32524
rect 27341 32515 27399 32521
rect 27982 32512 27988 32524
rect 28040 32512 28046 32564
rect 29549 32555 29607 32561
rect 29549 32521 29561 32555
rect 29595 32552 29607 32555
rect 29914 32552 29920 32564
rect 29595 32524 29920 32552
rect 29595 32521 29607 32524
rect 29549 32515 29607 32521
rect 29914 32512 29920 32524
rect 29972 32512 29978 32564
rect 21266 32444 21272 32496
rect 21324 32484 21330 32496
rect 25038 32484 25044 32496
rect 21324 32456 24932 32484
rect 24999 32456 25044 32484
rect 21324 32444 21330 32456
rect 20901 32419 20959 32425
rect 20901 32385 20913 32419
rect 20947 32416 20959 32419
rect 23474 32416 23480 32428
rect 20947 32388 23480 32416
rect 20947 32385 20959 32388
rect 20901 32379 20959 32385
rect 23474 32376 23480 32388
rect 23532 32376 23538 32428
rect 24904 32416 24932 32456
rect 25038 32444 25044 32456
rect 25096 32444 25102 32496
rect 30926 32416 30932 32428
rect 24904 32388 25636 32416
rect 30887 32388 30932 32416
rect 20211 32320 20300 32348
rect 20349 32351 20407 32357
rect 20211 32317 20223 32320
rect 20165 32311 20223 32317
rect 20349 32317 20361 32351
rect 20395 32317 20407 32351
rect 20349 32311 20407 32317
rect 20533 32351 20591 32357
rect 20533 32317 20545 32351
rect 20579 32317 20591 32351
rect 20533 32311 20591 32317
rect 20717 32351 20775 32357
rect 20717 32317 20729 32351
rect 20763 32348 20775 32351
rect 20990 32348 20996 32360
rect 20763 32320 20996 32348
rect 20763 32317 20775 32320
rect 20717 32311 20775 32317
rect 17497 32283 17555 32289
rect 17497 32280 17509 32283
rect 16684 32252 17509 32280
rect 17497 32249 17509 32252
rect 17543 32280 17555 32283
rect 17862 32280 17868 32292
rect 17543 32252 17868 32280
rect 17543 32249 17555 32252
rect 17497 32243 17555 32249
rect 17862 32240 17868 32252
rect 17920 32240 17926 32292
rect 17954 32240 17960 32292
rect 18012 32280 18018 32292
rect 19150 32280 19156 32292
rect 18012 32252 19156 32280
rect 18012 32240 18018 32252
rect 19150 32240 19156 32252
rect 19208 32240 19214 32292
rect 19613 32283 19671 32289
rect 19613 32249 19625 32283
rect 19659 32280 19671 32283
rect 20364 32280 20392 32311
rect 19659 32252 20392 32280
rect 19659 32249 19671 32252
rect 19613 32243 19671 32249
rect 20438 32240 20444 32292
rect 20496 32280 20502 32292
rect 20548 32280 20576 32311
rect 20990 32308 20996 32320
rect 21048 32308 21054 32360
rect 21266 32308 21272 32360
rect 21324 32348 21330 32360
rect 21453 32351 21511 32357
rect 21453 32348 21465 32351
rect 21324 32320 21465 32348
rect 21324 32308 21330 32320
rect 21453 32317 21465 32320
rect 21499 32317 21511 32351
rect 21453 32311 21511 32317
rect 21637 32351 21695 32357
rect 21637 32317 21649 32351
rect 21683 32317 21695 32351
rect 21637 32311 21695 32317
rect 21729 32351 21787 32357
rect 21729 32317 21741 32351
rect 21775 32317 21787 32351
rect 21729 32311 21787 32317
rect 21821 32351 21879 32357
rect 21821 32317 21833 32351
rect 21867 32348 21879 32351
rect 21910 32348 21916 32360
rect 21867 32320 21916 32348
rect 21867 32317 21879 32320
rect 21821 32311 21879 32317
rect 20496 32252 20576 32280
rect 20496 32240 20502 32252
rect 20622 32240 20628 32292
rect 20680 32280 20686 32292
rect 21652 32280 21680 32311
rect 20680 32252 21680 32280
rect 21744 32280 21772 32311
rect 21910 32308 21916 32320
rect 21968 32308 21974 32360
rect 22005 32351 22063 32357
rect 22005 32317 22017 32351
rect 22051 32348 22063 32351
rect 23382 32348 23388 32360
rect 22051 32320 23388 32348
rect 22051 32317 22063 32320
rect 22005 32311 22063 32317
rect 23382 32308 23388 32320
rect 23440 32308 23446 32360
rect 23753 32351 23811 32357
rect 23753 32317 23765 32351
rect 23799 32348 23811 32351
rect 23934 32348 23940 32360
rect 23799 32320 23940 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 23934 32308 23940 32320
rect 23992 32308 23998 32360
rect 24762 32308 24768 32360
rect 24820 32348 24826 32360
rect 25222 32348 25228 32360
rect 24820 32320 25228 32348
rect 24820 32308 24826 32320
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 25498 32348 25504 32360
rect 25459 32320 25504 32348
rect 25498 32308 25504 32320
rect 25556 32308 25562 32360
rect 24673 32283 24731 32289
rect 21744 32252 22048 32280
rect 20680 32240 20686 32252
rect 22020 32224 22048 32252
rect 24673 32249 24685 32283
rect 24719 32249 24731 32283
rect 24673 32243 24731 32249
rect 11808 32184 15516 32212
rect 15565 32215 15623 32221
rect 15565 32181 15577 32215
rect 15611 32212 15623 32215
rect 16942 32212 16948 32224
rect 15611 32184 16948 32212
rect 15611 32181 15623 32184
rect 15565 32175 15623 32181
rect 16942 32172 16948 32184
rect 17000 32172 17006 32224
rect 17310 32172 17316 32224
rect 17368 32212 17374 32224
rect 17589 32215 17647 32221
rect 17589 32212 17601 32215
rect 17368 32184 17601 32212
rect 17368 32172 17374 32184
rect 17589 32181 17601 32184
rect 17635 32212 17647 32215
rect 18322 32212 18328 32224
rect 17635 32184 18328 32212
rect 17635 32181 17647 32184
rect 17589 32175 17647 32181
rect 18322 32172 18328 32184
rect 18380 32172 18386 32224
rect 18782 32172 18788 32224
rect 18840 32212 18846 32224
rect 18966 32212 18972 32224
rect 18840 32184 18972 32212
rect 18840 32172 18846 32184
rect 18966 32172 18972 32184
rect 19024 32172 19030 32224
rect 19061 32215 19119 32221
rect 19061 32181 19073 32215
rect 19107 32212 19119 32215
rect 21361 32215 21419 32221
rect 21361 32212 21373 32215
rect 19107 32184 21373 32212
rect 19107 32181 19119 32184
rect 19061 32175 19119 32181
rect 21361 32181 21373 32184
rect 21407 32181 21419 32215
rect 21361 32175 21419 32181
rect 22002 32172 22008 32224
rect 22060 32172 22066 32224
rect 22189 32215 22247 32221
rect 22189 32181 22201 32215
rect 22235 32212 22247 32215
rect 22278 32212 22284 32224
rect 22235 32184 22284 32212
rect 22235 32181 22247 32184
rect 22189 32175 22247 32181
rect 22278 32172 22284 32184
rect 22336 32172 22342 32224
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 23750 32212 23756 32224
rect 23072 32184 23756 32212
rect 23072 32172 23078 32184
rect 23750 32172 23756 32184
rect 23808 32172 23814 32224
rect 24688 32212 24716 32243
rect 24854 32240 24860 32292
rect 24912 32289 24918 32292
rect 24912 32283 24931 32289
rect 24919 32249 24931 32283
rect 25608 32280 25636 32388
rect 30926 32376 30932 32388
rect 30984 32376 30990 32428
rect 25768 32351 25826 32357
rect 25768 32317 25780 32351
rect 25814 32348 25826 32351
rect 26142 32348 26148 32360
rect 25814 32320 26148 32348
rect 25814 32317 25826 32320
rect 25768 32311 25826 32317
rect 26142 32308 26148 32320
rect 26200 32308 26206 32360
rect 28442 32308 28448 32360
rect 28500 32357 28506 32360
rect 28500 32348 28512 32357
rect 28721 32351 28779 32357
rect 28500 32320 28545 32348
rect 28500 32311 28512 32320
rect 28721 32317 28733 32351
rect 28767 32348 28779 32351
rect 30374 32348 30380 32360
rect 28767 32320 30380 32348
rect 28767 32317 28779 32320
rect 28721 32311 28779 32317
rect 28500 32308 28506 32311
rect 30374 32308 30380 32320
rect 30432 32348 30438 32360
rect 30944 32348 30972 32376
rect 30432 32320 30972 32348
rect 30432 32308 30438 32320
rect 27522 32280 27528 32292
rect 25608 32252 27528 32280
rect 24912 32243 24931 32249
rect 24912 32240 24918 32243
rect 27522 32240 27528 32252
rect 27580 32240 27586 32292
rect 27982 32240 27988 32292
rect 28040 32280 28046 32292
rect 29086 32280 29092 32292
rect 28040 32252 29092 32280
rect 28040 32240 28046 32252
rect 29086 32240 29092 32252
rect 29144 32240 29150 32292
rect 30650 32240 30656 32292
rect 30708 32289 30714 32292
rect 30708 32280 30720 32289
rect 30708 32252 30753 32280
rect 30708 32243 30720 32252
rect 30708 32240 30714 32243
rect 25406 32212 25412 32224
rect 24688 32184 25412 32212
rect 25406 32172 25412 32184
rect 25464 32172 25470 32224
rect 25774 32172 25780 32224
rect 25832 32212 25838 32224
rect 25958 32212 25964 32224
rect 25832 32184 25964 32212
rect 25832 32172 25838 32184
rect 25958 32172 25964 32184
rect 26016 32172 26022 32224
rect 26050 32172 26056 32224
rect 26108 32212 26114 32224
rect 26881 32215 26939 32221
rect 26881 32212 26893 32215
rect 26108 32184 26893 32212
rect 26108 32172 26114 32184
rect 26881 32181 26893 32184
rect 26927 32181 26939 32215
rect 26881 32175 26939 32181
rect 1104 32122 32016 32144
rect 1104 32070 11253 32122
rect 11305 32070 11317 32122
rect 11369 32070 11381 32122
rect 11433 32070 11445 32122
rect 11497 32070 11509 32122
rect 11561 32070 21557 32122
rect 21609 32070 21621 32122
rect 21673 32070 21685 32122
rect 21737 32070 21749 32122
rect 21801 32070 21813 32122
rect 21865 32070 32016 32122
rect 1104 32048 32016 32070
rect 1949 32011 2007 32017
rect 1949 31977 1961 32011
rect 1995 32008 2007 32011
rect 2866 32008 2872 32020
rect 1995 31980 2872 32008
rect 1995 31977 2007 31980
rect 1949 31971 2007 31977
rect 2866 31968 2872 31980
rect 2924 31968 2930 32020
rect 3510 31968 3516 32020
rect 3568 32008 3574 32020
rect 5166 32008 5172 32020
rect 3568 31980 5172 32008
rect 3568 31968 3574 31980
rect 1489 31943 1547 31949
rect 1489 31909 1501 31943
rect 1535 31940 1547 31943
rect 2590 31940 2596 31952
rect 1535 31912 2596 31940
rect 1535 31909 1547 31912
rect 1489 31903 1547 31909
rect 2590 31900 2596 31912
rect 2648 31900 2654 31952
rect 2777 31943 2835 31949
rect 2777 31909 2789 31943
rect 2823 31940 2835 31943
rect 3142 31940 3148 31952
rect 2823 31912 3148 31940
rect 2823 31909 2835 31912
rect 2777 31903 2835 31909
rect 3142 31900 3148 31912
rect 3200 31900 3206 31952
rect 3789 31943 3847 31949
rect 3789 31909 3801 31943
rect 3835 31940 3847 31943
rect 4430 31940 4436 31952
rect 3835 31912 4436 31940
rect 3835 31909 3847 31912
rect 3789 31903 3847 31909
rect 4430 31900 4436 31912
rect 4488 31900 4494 31952
rect 4540 31949 4568 31980
rect 5166 31968 5172 31980
rect 5224 31968 5230 32020
rect 5810 31968 5816 32020
rect 5868 32008 5874 32020
rect 6914 32008 6920 32020
rect 5868 31980 6920 32008
rect 5868 31968 5874 31980
rect 6914 31968 6920 31980
rect 6972 31968 6978 32020
rect 7561 32011 7619 32017
rect 7561 31977 7573 32011
rect 7607 32008 7619 32011
rect 8754 32008 8760 32020
rect 7607 31980 8760 32008
rect 7607 31977 7619 31980
rect 7561 31971 7619 31977
rect 8754 31968 8760 31980
rect 8812 31968 8818 32020
rect 10778 31968 10784 32020
rect 10836 32008 10842 32020
rect 10965 32011 11023 32017
rect 10965 32008 10977 32011
rect 10836 31980 10977 32008
rect 10836 31968 10842 31980
rect 10965 31977 10977 31980
rect 11011 32008 11023 32011
rect 11054 32008 11060 32020
rect 11011 31980 11060 32008
rect 11011 31977 11023 31980
rect 10965 31971 11023 31977
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 11882 32008 11888 32020
rect 11843 31980 11888 32008
rect 11882 31968 11888 31980
rect 11940 31968 11946 32020
rect 13170 31968 13176 32020
rect 13228 32008 13234 32020
rect 13449 32011 13507 32017
rect 13449 32008 13461 32011
rect 13228 31980 13461 32008
rect 13228 31968 13234 31980
rect 13449 31977 13461 31980
rect 13495 31977 13507 32011
rect 13449 31971 13507 31977
rect 13633 32011 13691 32017
rect 13633 31977 13645 32011
rect 13679 32008 13691 32011
rect 14274 32008 14280 32020
rect 13679 31980 14280 32008
rect 13679 31977 13691 31980
rect 13633 31971 13691 31977
rect 14274 31968 14280 31980
rect 14332 31968 14338 32020
rect 19794 32008 19800 32020
rect 15672 31980 19800 32008
rect 4525 31943 4583 31949
rect 4525 31909 4537 31943
rect 4571 31909 4583 31943
rect 4525 31903 4583 31909
rect 4741 31943 4799 31949
rect 4741 31909 4753 31943
rect 4787 31940 4799 31943
rect 5534 31940 5540 31952
rect 4787 31912 5540 31940
rect 4787 31909 4799 31912
rect 4741 31903 4799 31909
rect 5534 31900 5540 31912
rect 5592 31900 5598 31952
rect 5718 31900 5724 31952
rect 5776 31940 5782 31952
rect 6730 31940 6736 31952
rect 5776 31912 6736 31940
rect 5776 31900 5782 31912
rect 6730 31900 6736 31912
rect 6788 31900 6794 31952
rect 7834 31900 7840 31952
rect 7892 31940 7898 31952
rect 8113 31943 8171 31949
rect 8113 31940 8125 31943
rect 7892 31912 8125 31940
rect 7892 31900 7898 31912
rect 8113 31909 8125 31912
rect 8159 31940 8171 31943
rect 8938 31940 8944 31952
rect 8159 31912 8708 31940
rect 8159 31909 8171 31912
rect 8113 31903 8171 31909
rect 1670 31832 1676 31884
rect 1728 31872 1734 31884
rect 2222 31872 2228 31884
rect 1728 31844 2084 31872
rect 2183 31844 2228 31872
rect 1728 31832 1734 31844
rect 1946 31804 1952 31816
rect 1907 31776 1952 31804
rect 1946 31764 1952 31776
rect 2004 31764 2010 31816
rect 2056 31804 2084 31844
rect 2222 31832 2228 31844
rect 2280 31832 2286 31884
rect 2685 31875 2743 31881
rect 2685 31872 2697 31875
rect 2332 31844 2697 31872
rect 2332 31804 2360 31844
rect 2685 31841 2697 31844
rect 2731 31841 2743 31875
rect 4065 31875 4123 31881
rect 4065 31872 4077 31875
rect 2685 31835 2743 31841
rect 3988 31844 4077 31872
rect 3326 31804 3332 31816
rect 2056 31776 2360 31804
rect 2424 31776 3332 31804
rect 1302 31696 1308 31748
rect 1360 31736 1366 31748
rect 2424 31736 2452 31776
rect 3326 31764 3332 31776
rect 3384 31764 3390 31816
rect 3786 31804 3792 31816
rect 3747 31776 3792 31804
rect 3786 31764 3792 31776
rect 3844 31764 3850 31816
rect 3988 31736 4016 31844
rect 4065 31841 4077 31844
rect 4111 31841 4123 31875
rect 5350 31872 5356 31884
rect 5311 31844 5356 31872
rect 4065 31835 4123 31841
rect 5350 31832 5356 31844
rect 5408 31832 5414 31884
rect 6638 31832 6644 31884
rect 6696 31872 6702 31884
rect 7285 31875 7343 31881
rect 7285 31872 7297 31875
rect 6696 31844 7297 31872
rect 6696 31832 6702 31844
rect 7285 31841 7297 31844
rect 7331 31841 7343 31875
rect 8202 31872 8208 31884
rect 8163 31844 8208 31872
rect 7285 31835 7343 31841
rect 8202 31832 8208 31844
rect 8260 31832 8266 31884
rect 8680 31881 8708 31912
rect 8772 31912 8944 31940
rect 8772 31881 8800 31912
rect 8938 31900 8944 31912
rect 8996 31900 9002 31952
rect 9852 31943 9910 31949
rect 9852 31909 9864 31943
rect 9898 31940 9910 31943
rect 10594 31940 10600 31952
rect 9898 31912 10600 31940
rect 9898 31909 9910 31912
rect 9852 31903 9910 31909
rect 10594 31900 10600 31912
rect 10652 31900 10658 31952
rect 12084 31912 12940 31940
rect 8665 31875 8723 31881
rect 8665 31841 8677 31875
rect 8711 31841 8723 31875
rect 8665 31835 8723 31841
rect 8757 31875 8815 31881
rect 8757 31841 8769 31875
rect 8803 31841 8815 31875
rect 8757 31835 8815 31841
rect 8849 31875 8907 31881
rect 8849 31841 8861 31875
rect 8895 31841 8907 31875
rect 8849 31835 8907 31841
rect 4246 31764 4252 31816
rect 4304 31804 4310 31816
rect 4706 31804 4712 31816
rect 4304 31776 4712 31804
rect 4304 31764 4310 31776
rect 4706 31764 4712 31776
rect 4764 31764 4770 31816
rect 5442 31804 5448 31816
rect 5092 31776 5448 31804
rect 5092 31736 5120 31776
rect 5442 31764 5448 31776
rect 5500 31804 5506 31816
rect 6365 31807 6423 31813
rect 6365 31804 6377 31807
rect 5500 31776 6377 31804
rect 5500 31764 5506 31776
rect 6365 31773 6377 31776
rect 6411 31773 6423 31807
rect 7558 31804 7564 31816
rect 7519 31776 7564 31804
rect 6365 31767 6423 31773
rect 7558 31764 7564 31776
rect 7616 31764 7622 31816
rect 7650 31764 7656 31816
rect 7708 31804 7714 31816
rect 8294 31804 8300 31816
rect 7708 31776 8300 31804
rect 7708 31764 7714 31776
rect 8294 31764 8300 31776
rect 8352 31804 8358 31816
rect 8864 31804 8892 31835
rect 10318 31832 10324 31884
rect 10376 31872 10382 31884
rect 10376 31844 10732 31872
rect 10376 31832 10382 31844
rect 10704 31816 10732 31844
rect 11146 31832 11152 31884
rect 11204 31872 11210 31884
rect 12084 31881 12112 31912
rect 12912 31884 12940 31912
rect 13814 31900 13820 31952
rect 13872 31940 13878 31952
rect 14185 31943 14243 31949
rect 14185 31940 14197 31943
rect 13872 31912 14197 31940
rect 13872 31900 13878 31912
rect 14185 31909 14197 31912
rect 14231 31909 14243 31943
rect 14185 31903 14243 31909
rect 12069 31875 12127 31881
rect 12069 31872 12081 31875
rect 11204 31844 12081 31872
rect 11204 31832 11210 31844
rect 12069 31841 12081 31844
rect 12115 31841 12127 31875
rect 12069 31835 12127 31841
rect 12437 31875 12495 31881
rect 12437 31841 12449 31875
rect 12483 31872 12495 31875
rect 12483 31844 12572 31872
rect 12483 31841 12495 31844
rect 12437 31835 12495 31841
rect 8352 31776 8892 31804
rect 8352 31764 8358 31776
rect 9490 31764 9496 31816
rect 9548 31804 9554 31816
rect 9585 31807 9643 31813
rect 9585 31804 9597 31807
rect 9548 31776 9597 31804
rect 9548 31764 9554 31776
rect 9585 31773 9597 31776
rect 9631 31773 9643 31807
rect 9585 31767 9643 31773
rect 10686 31764 10692 31816
rect 10744 31764 10750 31816
rect 10962 31764 10968 31816
rect 11020 31804 11026 31816
rect 11698 31804 11704 31816
rect 11020 31776 11704 31804
rect 11020 31764 11026 31776
rect 11698 31764 11704 31776
rect 11756 31804 11762 31816
rect 12253 31807 12311 31813
rect 12253 31804 12265 31807
rect 11756 31776 12265 31804
rect 11756 31764 11762 31776
rect 12253 31773 12265 31776
rect 12299 31773 12311 31807
rect 12253 31767 12311 31773
rect 12345 31807 12403 31813
rect 12345 31773 12357 31807
rect 12391 31773 12403 31807
rect 12345 31767 12403 31773
rect 1360 31708 2452 31736
rect 2976 31708 4016 31736
rect 4724 31708 5120 31736
rect 1360 31696 1366 31708
rect 0 31668 800 31682
rect 2976 31680 3004 31708
rect 4724 31680 4752 31708
rect 6454 31696 6460 31748
rect 6512 31736 6518 31748
rect 9214 31736 9220 31748
rect 6512 31708 9220 31736
rect 6512 31696 6518 31708
rect 9214 31696 9220 31708
rect 9272 31696 9278 31748
rect 12360 31736 12388 31767
rect 12176 31708 12388 31736
rect 12176 31680 12204 31708
rect 1578 31668 1584 31680
rect 0 31640 1584 31668
rect 0 31626 800 31640
rect 1578 31628 1584 31640
rect 1636 31628 1642 31680
rect 2133 31671 2191 31677
rect 2133 31637 2145 31671
rect 2179 31668 2191 31671
rect 2314 31668 2320 31680
rect 2179 31640 2320 31668
rect 2179 31637 2191 31640
rect 2133 31631 2191 31637
rect 2314 31628 2320 31640
rect 2372 31628 2378 31680
rect 2958 31628 2964 31680
rect 3016 31628 3022 31680
rect 3973 31671 4031 31677
rect 3973 31637 3985 31671
rect 4019 31668 4031 31671
rect 4154 31668 4160 31680
rect 4019 31640 4160 31668
rect 4019 31637 4031 31640
rect 3973 31631 4031 31637
rect 4154 31628 4160 31640
rect 4212 31628 4218 31680
rect 4706 31668 4712 31680
rect 4667 31640 4712 31668
rect 4706 31628 4712 31640
rect 4764 31628 4770 31680
rect 4893 31671 4951 31677
rect 4893 31637 4905 31671
rect 4939 31668 4951 31671
rect 4982 31668 4988 31680
rect 4939 31640 4988 31668
rect 4939 31637 4951 31640
rect 4893 31631 4951 31637
rect 4982 31628 4988 31640
rect 5040 31628 5046 31680
rect 5442 31668 5448 31680
rect 5403 31640 5448 31668
rect 5442 31628 5448 31640
rect 5500 31628 5506 31680
rect 6638 31628 6644 31680
rect 6696 31668 6702 31680
rect 7377 31671 7435 31677
rect 7377 31668 7389 31671
rect 6696 31640 7389 31668
rect 6696 31628 6702 31640
rect 7377 31637 7389 31640
rect 7423 31637 7435 31671
rect 7377 31631 7435 31637
rect 8110 31628 8116 31680
rect 8168 31668 8174 31680
rect 8478 31668 8484 31680
rect 8168 31640 8484 31668
rect 8168 31628 8174 31640
rect 8478 31628 8484 31640
rect 8536 31628 8542 31680
rect 12158 31628 12164 31680
rect 12216 31628 12222 31680
rect 12544 31668 12572 31844
rect 12618 31832 12624 31884
rect 12676 31872 12682 31884
rect 12676 31844 12721 31872
rect 12676 31832 12682 31844
rect 12894 31832 12900 31884
rect 12952 31872 12958 31884
rect 13081 31875 13139 31881
rect 13081 31872 13093 31875
rect 12952 31844 13093 31872
rect 12952 31832 12958 31844
rect 13081 31841 13093 31844
rect 13127 31841 13139 31875
rect 13081 31835 13139 31841
rect 13354 31832 13360 31884
rect 13412 31872 13418 31884
rect 14093 31875 14151 31881
rect 14093 31872 14105 31875
rect 13412 31844 14105 31872
rect 13412 31832 13418 31844
rect 14093 31841 14105 31844
rect 14139 31841 14151 31875
rect 14093 31835 14151 31841
rect 14918 31832 14924 31884
rect 14976 31872 14982 31884
rect 15197 31875 15255 31881
rect 15197 31872 15209 31875
rect 14976 31844 15209 31872
rect 14976 31832 14982 31844
rect 15197 31841 15209 31844
rect 15243 31841 15255 31875
rect 15378 31872 15384 31884
rect 15339 31844 15384 31872
rect 15197 31835 15255 31841
rect 15378 31832 15384 31844
rect 15436 31832 15442 31884
rect 15577 31881 15635 31887
rect 15577 31847 15589 31881
rect 15623 31878 15635 31881
rect 15672 31878 15700 31980
rect 19794 31968 19800 31980
rect 19852 31968 19858 32020
rect 20530 31968 20536 32020
rect 20588 32008 20594 32020
rect 20714 32008 20720 32020
rect 20588 31980 20720 32008
rect 20588 31968 20594 31980
rect 20714 31968 20720 31980
rect 20772 31968 20778 32020
rect 20990 31968 20996 32020
rect 21048 32008 21054 32020
rect 21910 32008 21916 32020
rect 21048 31980 21916 32008
rect 21048 31968 21054 31980
rect 21910 31968 21916 31980
rect 21968 31968 21974 32020
rect 22112 31980 23152 32008
rect 16482 31900 16488 31952
rect 16540 31940 16546 31952
rect 16574 31940 16580 31952
rect 16540 31912 16580 31940
rect 16540 31900 16546 31912
rect 16574 31900 16580 31912
rect 16632 31900 16638 31952
rect 18233 31943 18291 31949
rect 18233 31940 18245 31943
rect 17144 31912 18245 31940
rect 15623 31850 15700 31878
rect 15749 31875 15807 31881
rect 15623 31847 15635 31850
rect 15577 31841 15635 31847
rect 15749 31841 15761 31875
rect 15795 31872 15807 31875
rect 15838 31872 15844 31884
rect 15795 31844 15844 31872
rect 15795 31841 15807 31844
rect 15749 31835 15807 31841
rect 15838 31832 15844 31844
rect 15896 31832 15902 31884
rect 16114 31872 16120 31884
rect 15957 31844 16120 31872
rect 15102 31764 15108 31816
rect 15160 31804 15166 31816
rect 15396 31804 15424 31832
rect 15160 31776 15424 31804
rect 15473 31807 15531 31813
rect 15160 31764 15166 31776
rect 15473 31773 15485 31807
rect 15519 31804 15531 31807
rect 15654 31804 15660 31816
rect 15519 31776 15660 31804
rect 15519 31773 15531 31776
rect 15473 31767 15531 31773
rect 15654 31764 15660 31776
rect 15712 31804 15718 31816
rect 15957 31804 15985 31844
rect 16114 31832 16120 31844
rect 16172 31832 16178 31884
rect 16758 31832 16764 31884
rect 16816 31872 16822 31884
rect 17144 31881 17172 31912
rect 18233 31909 18245 31912
rect 18279 31909 18291 31943
rect 18233 31903 18291 31909
rect 18598 31900 18604 31952
rect 18656 31940 18662 31952
rect 18782 31940 18788 31952
rect 18656 31912 18788 31940
rect 18656 31900 18662 31912
rect 18782 31900 18788 31912
rect 18840 31940 18846 31952
rect 22112 31940 22140 31980
rect 23124 31940 23152 31980
rect 23198 31968 23204 32020
rect 23256 32008 23262 32020
rect 23753 32011 23811 32017
rect 23753 32008 23765 32011
rect 23256 31980 23765 32008
rect 23256 31968 23262 31980
rect 23753 31977 23765 31980
rect 23799 32008 23811 32011
rect 26234 32008 26240 32020
rect 23799 31980 26240 32008
rect 23799 31977 23811 31980
rect 23753 31971 23811 31977
rect 26234 31968 26240 31980
rect 26292 31968 26298 32020
rect 26602 31968 26608 32020
rect 26660 32008 26666 32020
rect 26973 32011 27031 32017
rect 26973 32008 26985 32011
rect 26660 31980 26985 32008
rect 26660 31968 26666 31980
rect 26973 31977 26985 31980
rect 27019 31977 27031 32011
rect 27522 32008 27528 32020
rect 27483 31980 27528 32008
rect 26973 31971 27031 31977
rect 27522 31968 27528 31980
rect 27580 31968 27586 32020
rect 28810 32008 28816 32020
rect 28771 31980 28816 32008
rect 28810 31968 28816 31980
rect 28868 31968 28874 32020
rect 24486 31940 24492 31952
rect 18840 31912 22140 31940
rect 22204 31912 23076 31940
rect 23124 31912 24492 31940
rect 18840 31900 18846 31912
rect 16945 31875 17003 31881
rect 16945 31872 16957 31875
rect 16816 31844 16957 31872
rect 16816 31832 16822 31844
rect 16945 31841 16957 31844
rect 16991 31841 17003 31875
rect 16945 31835 17003 31841
rect 17129 31875 17187 31881
rect 17129 31841 17141 31875
rect 17175 31841 17187 31875
rect 17494 31872 17500 31884
rect 17455 31844 17500 31872
rect 17129 31835 17187 31841
rect 17494 31832 17500 31844
rect 17552 31872 17558 31884
rect 18141 31875 18199 31881
rect 18141 31872 18153 31875
rect 17552 31844 18153 31872
rect 17552 31832 17558 31844
rect 18141 31841 18153 31844
rect 18187 31841 18199 31875
rect 18141 31835 18199 31841
rect 19702 31832 19708 31884
rect 19760 31872 19766 31884
rect 20162 31872 20168 31884
rect 19760 31844 20168 31872
rect 19760 31832 19766 31844
rect 20162 31832 20168 31844
rect 20220 31872 20226 31884
rect 20622 31872 20628 31884
rect 20220 31844 20628 31872
rect 20220 31832 20226 31844
rect 20622 31832 20628 31844
rect 20680 31832 20686 31884
rect 20990 31872 20996 31884
rect 20951 31844 20996 31872
rect 20990 31832 20996 31844
rect 21048 31832 21054 31884
rect 21174 31872 21180 31884
rect 21135 31844 21180 31872
rect 21174 31832 21180 31844
rect 21232 31832 21238 31884
rect 22002 31832 22008 31884
rect 22060 31832 22066 31884
rect 15712 31776 15985 31804
rect 15712 31764 15718 31776
rect 16022 31764 16028 31816
rect 16080 31804 16086 31816
rect 17218 31804 17224 31816
rect 16080 31776 17224 31804
rect 16080 31764 16086 31776
rect 17218 31764 17224 31776
rect 17276 31764 17282 31816
rect 17313 31807 17371 31813
rect 17313 31773 17325 31807
rect 17359 31804 17371 31807
rect 17402 31804 17408 31816
rect 17359 31776 17408 31804
rect 17359 31773 17371 31776
rect 17313 31767 17371 31773
rect 17402 31764 17408 31776
rect 17460 31764 17466 31816
rect 17681 31807 17739 31813
rect 17681 31773 17693 31807
rect 17727 31804 17739 31807
rect 17954 31804 17960 31816
rect 17727 31776 17960 31804
rect 17727 31773 17739 31776
rect 17681 31767 17739 31773
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18966 31764 18972 31816
rect 19024 31804 19030 31816
rect 19153 31807 19211 31813
rect 19153 31804 19165 31807
rect 19024 31776 19165 31804
rect 19024 31764 19030 31776
rect 19153 31773 19165 31776
rect 19199 31773 19211 31807
rect 19153 31767 19211 31773
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31804 19487 31807
rect 19886 31804 19892 31816
rect 19475 31776 19892 31804
rect 19475 31773 19487 31776
rect 19429 31767 19487 31773
rect 19886 31764 19892 31776
rect 19944 31804 19950 31816
rect 20809 31807 20867 31813
rect 20809 31804 20821 31807
rect 19944 31776 20821 31804
rect 19944 31764 19950 31776
rect 20809 31773 20821 31776
rect 20855 31773 20867 31807
rect 20809 31767 20867 31773
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31804 20959 31807
rect 22020 31804 22048 31832
rect 20947 31776 22048 31804
rect 20947 31773 20959 31776
rect 20901 31767 20959 31773
rect 12986 31696 12992 31748
rect 13044 31736 13050 31748
rect 13044 31708 20576 31736
rect 13044 31696 13050 31708
rect 12710 31668 12716 31680
rect 12544 31640 12716 31668
rect 12710 31628 12716 31640
rect 12768 31668 12774 31680
rect 13446 31668 13452 31680
rect 12768 31640 13452 31668
rect 12768 31628 12774 31640
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 13538 31628 13544 31680
rect 13596 31668 13602 31680
rect 13906 31668 13912 31680
rect 13596 31640 13912 31668
rect 13596 31628 13602 31640
rect 13906 31628 13912 31640
rect 13964 31628 13970 31680
rect 15010 31668 15016 31680
rect 14971 31640 15016 31668
rect 15010 31628 15016 31640
rect 15068 31628 15074 31680
rect 20438 31668 20444 31680
rect 20399 31640 20444 31668
rect 20438 31628 20444 31640
rect 20496 31628 20502 31680
rect 20548 31668 20576 31708
rect 20622 31696 20628 31748
rect 20680 31736 20686 31748
rect 21174 31736 21180 31748
rect 20680 31708 21180 31736
rect 20680 31696 20686 31708
rect 21174 31696 21180 31708
rect 21232 31696 21238 31748
rect 21821 31739 21879 31745
rect 21821 31705 21833 31739
rect 21867 31736 21879 31739
rect 21910 31736 21916 31748
rect 21867 31708 21916 31736
rect 21867 31705 21879 31708
rect 21821 31699 21879 31705
rect 21910 31696 21916 31708
rect 21968 31696 21974 31748
rect 22002 31696 22008 31748
rect 22060 31736 22066 31748
rect 22204 31736 22232 31912
rect 22554 31832 22560 31884
rect 22612 31872 22618 31884
rect 22934 31875 22992 31881
rect 22934 31872 22946 31875
rect 22612 31844 22946 31872
rect 22612 31832 22618 31844
rect 22934 31841 22946 31844
rect 22980 31841 22992 31875
rect 23048 31872 23076 31912
rect 24486 31900 24492 31912
rect 24544 31900 24550 31952
rect 25498 31940 25504 31952
rect 24780 31912 25504 31940
rect 23201 31875 23259 31881
rect 23201 31872 23213 31875
rect 23048 31844 23213 31872
rect 22934 31835 22992 31841
rect 23201 31841 23213 31844
rect 23247 31872 23259 31875
rect 24780 31872 24808 31912
rect 25148 31881 25176 31912
rect 25498 31900 25504 31912
rect 25556 31900 25562 31952
rect 23247 31844 24808 31872
rect 24877 31875 24935 31881
rect 23247 31841 23259 31844
rect 23201 31835 23259 31841
rect 24877 31841 24889 31875
rect 24923 31872 24935 31875
rect 25133 31875 25191 31881
rect 24923 31844 25084 31872
rect 24923 31841 24935 31844
rect 24877 31835 24935 31841
rect 25056 31804 25084 31844
rect 25133 31841 25145 31875
rect 25179 31841 25191 31875
rect 25133 31835 25191 31841
rect 25222 31832 25228 31884
rect 25280 31872 25286 31884
rect 25406 31872 25412 31884
rect 25280 31844 25412 31872
rect 25280 31832 25286 31844
rect 25406 31832 25412 31844
rect 25464 31872 25470 31884
rect 25593 31875 25651 31881
rect 25593 31872 25605 31875
rect 25464 31844 25605 31872
rect 25464 31832 25470 31844
rect 25593 31841 25605 31844
rect 25639 31841 25651 31875
rect 25593 31835 25651 31841
rect 25774 31832 25780 31884
rect 25832 31872 25838 31884
rect 25832 31844 25877 31872
rect 25832 31832 25838 31844
rect 25958 31832 25964 31884
rect 26016 31872 26022 31884
rect 26145 31875 26203 31881
rect 26016 31844 26061 31872
rect 26016 31832 26022 31844
rect 26145 31841 26157 31875
rect 26191 31870 26203 31875
rect 26252 31870 26280 31968
rect 29362 31900 29368 31952
rect 29420 31940 29426 31952
rect 29926 31943 29984 31949
rect 29926 31940 29938 31943
rect 29420 31912 29938 31940
rect 29420 31900 29426 31912
rect 29926 31909 29938 31912
rect 29972 31909 29984 31943
rect 29926 31903 29984 31909
rect 29638 31872 29644 31884
rect 26191 31842 26280 31870
rect 28966 31844 29644 31872
rect 26191 31841 26203 31842
rect 26145 31835 26203 31841
rect 25498 31804 25504 31816
rect 25056 31776 25504 31804
rect 25498 31764 25504 31776
rect 25556 31764 25562 31816
rect 25869 31807 25927 31813
rect 25869 31773 25881 31807
rect 25915 31804 25927 31807
rect 26326 31804 26332 31816
rect 25915 31776 26332 31804
rect 25915 31773 25927 31776
rect 25869 31767 25927 31773
rect 26326 31764 26332 31776
rect 26384 31764 26390 31816
rect 26510 31764 26516 31816
rect 26568 31804 26574 31816
rect 28077 31807 28135 31813
rect 28077 31804 28089 31807
rect 26568 31776 28089 31804
rect 26568 31764 26574 31776
rect 28077 31773 28089 31776
rect 28123 31773 28135 31807
rect 28077 31767 28135 31773
rect 22060 31708 22232 31736
rect 22060 31696 22066 31708
rect 25222 31696 25228 31748
rect 25280 31736 25286 31748
rect 25590 31736 25596 31748
rect 25280 31708 25596 31736
rect 25280 31696 25286 31708
rect 25590 31696 25596 31708
rect 25648 31696 25654 31748
rect 28966 31736 28994 31844
rect 29638 31832 29644 31844
rect 29696 31832 29702 31884
rect 30193 31875 30251 31881
rect 30193 31841 30205 31875
rect 30239 31872 30251 31875
rect 30374 31872 30380 31884
rect 30239 31844 30380 31872
rect 30239 31841 30251 31844
rect 30193 31835 30251 31841
rect 30374 31832 30380 31844
rect 30432 31832 30438 31884
rect 31113 31875 31171 31881
rect 31113 31841 31125 31875
rect 31159 31872 31171 31875
rect 31478 31872 31484 31884
rect 31159 31844 31484 31872
rect 31159 31841 31171 31844
rect 31113 31835 31171 31841
rect 31478 31832 31484 31844
rect 31536 31832 31542 31884
rect 26068 31708 28994 31736
rect 23934 31668 23940 31680
rect 20548 31640 23940 31668
rect 23934 31628 23940 31640
rect 23992 31628 23998 31680
rect 24486 31628 24492 31680
rect 24544 31668 24550 31680
rect 26068 31668 26096 31708
rect 26326 31668 26332 31680
rect 24544 31640 26096 31668
rect 26287 31640 26332 31668
rect 24544 31628 24550 31640
rect 26326 31628 26332 31640
rect 26384 31628 26390 31680
rect 31297 31671 31355 31677
rect 31297 31637 31309 31671
rect 31343 31668 31355 31671
rect 32320 31668 33120 31682
rect 31343 31640 33120 31668
rect 31343 31637 31355 31640
rect 31297 31631 31355 31637
rect 32320 31626 33120 31640
rect 1104 31578 32016 31600
rect 1104 31526 6102 31578
rect 6154 31526 6166 31578
rect 6218 31526 6230 31578
rect 6282 31526 6294 31578
rect 6346 31526 6358 31578
rect 6410 31526 16405 31578
rect 16457 31526 16469 31578
rect 16521 31526 16533 31578
rect 16585 31526 16597 31578
rect 16649 31526 16661 31578
rect 16713 31526 26709 31578
rect 26761 31526 26773 31578
rect 26825 31526 26837 31578
rect 26889 31526 26901 31578
rect 26953 31526 26965 31578
rect 27017 31526 32016 31578
rect 1104 31504 32016 31526
rect 2774 31424 2780 31476
rect 2832 31464 2838 31476
rect 3602 31464 3608 31476
rect 2832 31436 3608 31464
rect 2832 31424 2838 31436
rect 3602 31424 3608 31436
rect 3660 31424 3666 31476
rect 3881 31467 3939 31473
rect 3881 31433 3893 31467
rect 3927 31464 3939 31467
rect 4154 31464 4160 31476
rect 3927 31436 4160 31464
rect 3927 31433 3939 31436
rect 3881 31427 3939 31433
rect 4154 31424 4160 31436
rect 4212 31464 4218 31476
rect 4212 31436 5672 31464
rect 4212 31424 4218 31436
rect 2041 31399 2099 31405
rect 2041 31365 2053 31399
rect 2087 31396 2099 31399
rect 2314 31396 2320 31408
rect 2087 31368 2320 31396
rect 2087 31365 2099 31368
rect 2041 31359 2099 31365
rect 2314 31356 2320 31368
rect 2372 31356 2378 31408
rect 3418 31356 3424 31408
rect 3476 31396 3482 31408
rect 4062 31396 4068 31408
rect 3476 31368 4068 31396
rect 3476 31356 3482 31368
rect 4062 31356 4068 31368
rect 4120 31356 4126 31408
rect 5077 31399 5135 31405
rect 5077 31365 5089 31399
rect 5123 31396 5135 31399
rect 5644 31396 5672 31436
rect 5902 31424 5908 31476
rect 5960 31464 5966 31476
rect 6546 31464 6552 31476
rect 5960 31436 6552 31464
rect 5960 31424 5966 31436
rect 6546 31424 6552 31436
rect 6604 31424 6610 31476
rect 7006 31464 7012 31476
rect 6967 31436 7012 31464
rect 7006 31424 7012 31436
rect 7064 31424 7070 31476
rect 7650 31464 7656 31476
rect 7611 31436 7656 31464
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 8018 31424 8024 31476
rect 8076 31464 8082 31476
rect 8205 31467 8263 31473
rect 8205 31464 8217 31467
rect 8076 31436 8217 31464
rect 8076 31424 8082 31436
rect 8205 31433 8217 31436
rect 8251 31464 8263 31467
rect 8938 31464 8944 31476
rect 8251 31436 8944 31464
rect 8251 31433 8263 31436
rect 8205 31427 8263 31433
rect 8938 31424 8944 31436
rect 8996 31424 9002 31476
rect 13170 31464 13176 31476
rect 9508 31436 13032 31464
rect 13131 31436 13176 31464
rect 7024 31396 7052 31424
rect 9508 31396 9536 31436
rect 5123 31368 5589 31396
rect 5644 31368 7052 31396
rect 7484 31368 9536 31396
rect 10873 31399 10931 31405
rect 5123 31365 5135 31368
rect 5077 31359 5135 31365
rect 3234 31328 3240 31340
rect 3195 31300 3240 31328
rect 3234 31288 3240 31300
rect 3292 31288 3298 31340
rect 4430 31288 4436 31340
rect 4488 31328 4494 31340
rect 4893 31331 4951 31337
rect 4893 31328 4905 31331
rect 4488 31300 4905 31328
rect 4488 31288 4494 31300
rect 4893 31297 4905 31300
rect 4939 31297 4951 31331
rect 4893 31291 4951 31297
rect 5169 31331 5227 31337
rect 5169 31297 5181 31331
rect 5215 31328 5227 31331
rect 5442 31328 5448 31340
rect 5215 31300 5448 31328
rect 5215 31297 5227 31300
rect 5169 31291 5227 31297
rect 5442 31288 5448 31300
rect 5500 31288 5506 31340
rect 1578 31220 1584 31272
rect 1636 31260 1642 31272
rect 1857 31263 1915 31269
rect 1857 31260 1869 31263
rect 1636 31232 1869 31260
rect 1636 31220 1642 31232
rect 1857 31229 1869 31232
rect 1903 31229 1915 31263
rect 2958 31260 2964 31272
rect 2919 31232 2964 31260
rect 1857 31223 1915 31229
rect 2958 31220 2964 31232
rect 3016 31220 3022 31272
rect 3050 31220 3056 31272
rect 3108 31260 3114 31272
rect 4617 31263 4675 31269
rect 4617 31260 4629 31263
rect 3108 31232 3201 31260
rect 3252 31232 4629 31260
rect 3108 31220 3114 31232
rect 3160 31124 3188 31232
rect 3252 31201 3280 31232
rect 4617 31229 4629 31232
rect 4663 31229 4675 31263
rect 4617 31223 4675 31229
rect 5074 31220 5080 31272
rect 5132 31260 5138 31272
rect 5261 31263 5319 31269
rect 5261 31260 5273 31263
rect 5132 31232 5273 31260
rect 5132 31220 5138 31232
rect 5261 31229 5273 31232
rect 5307 31229 5319 31263
rect 5261 31223 5319 31229
rect 3237 31195 3295 31201
rect 3237 31161 3249 31195
rect 3283 31161 3295 31195
rect 3237 31155 3295 31161
rect 4246 31152 4252 31204
rect 4304 31192 4310 31204
rect 5442 31192 5448 31204
rect 4304 31164 5448 31192
rect 4304 31152 4310 31164
rect 5442 31152 5448 31164
rect 5500 31152 5506 31204
rect 5561 31192 5589 31368
rect 6457 31263 6515 31269
rect 6457 31229 6469 31263
rect 6503 31260 6515 31263
rect 6546 31260 6552 31272
rect 6503 31232 6552 31260
rect 6503 31229 6515 31232
rect 6457 31223 6515 31229
rect 6546 31220 6552 31232
rect 6604 31220 6610 31272
rect 7484 31260 7512 31368
rect 10873 31365 10885 31399
rect 10919 31396 10931 31399
rect 10962 31396 10968 31408
rect 10919 31368 10968 31396
rect 10919 31365 10931 31368
rect 10873 31359 10931 31365
rect 10962 31356 10968 31368
rect 11020 31396 11026 31408
rect 11606 31396 11612 31408
rect 11020 31368 11612 31396
rect 11020 31356 11026 31368
rect 7834 31288 7840 31340
rect 7892 31328 7898 31340
rect 8941 31331 8999 31337
rect 8941 31328 8953 31331
rect 7892 31300 8953 31328
rect 7892 31288 7898 31300
rect 8941 31297 8953 31300
rect 8987 31328 8999 31331
rect 9122 31328 9128 31340
rect 8987 31300 9128 31328
rect 8987 31297 8999 31300
rect 8941 31291 8999 31297
rect 9122 31288 9128 31300
rect 9180 31288 9186 31340
rect 6840 31232 7512 31260
rect 7561 31263 7619 31269
rect 6840 31192 6868 31232
rect 7561 31229 7573 31263
rect 7607 31260 7619 31263
rect 8662 31260 8668 31272
rect 7607 31232 8668 31260
rect 7607 31229 7619 31232
rect 7561 31223 7619 31229
rect 8662 31220 8668 31232
rect 8720 31220 8726 31272
rect 9398 31220 9404 31272
rect 9456 31260 9462 31272
rect 9493 31263 9551 31269
rect 9493 31260 9505 31263
rect 9456 31232 9505 31260
rect 9456 31220 9462 31232
rect 9493 31229 9505 31232
rect 9539 31229 9551 31263
rect 9493 31223 9551 31229
rect 11054 31220 11060 31272
rect 11112 31260 11118 31272
rect 11532 31269 11560 31368
rect 11606 31356 11612 31368
rect 11664 31356 11670 31408
rect 12526 31396 12532 31408
rect 12487 31368 12532 31396
rect 12526 31356 12532 31368
rect 12584 31356 12590 31408
rect 11793 31331 11851 31337
rect 11793 31297 11805 31331
rect 11839 31328 11851 31331
rect 12158 31328 12164 31340
rect 11839 31300 12164 31328
rect 11839 31297 11851 31300
rect 11793 31291 11851 31297
rect 12158 31288 12164 31300
rect 12216 31288 12222 31340
rect 11517 31263 11575 31269
rect 11112 31232 11468 31260
rect 11112 31220 11118 31232
rect 5561 31164 6868 31192
rect 7006 31152 7012 31204
rect 7064 31192 7070 31204
rect 8478 31192 8484 31204
rect 7064 31164 8484 31192
rect 7064 31152 7070 31164
rect 8478 31152 8484 31164
rect 8536 31152 8542 31204
rect 9760 31195 9818 31201
rect 9760 31161 9772 31195
rect 9806 31192 9818 31195
rect 11333 31195 11391 31201
rect 11333 31192 11345 31195
rect 9806 31164 11345 31192
rect 9806 31161 9818 31164
rect 9760 31155 9818 31161
rect 11333 31161 11345 31164
rect 11379 31161 11391 31195
rect 11440 31192 11468 31232
rect 11517 31229 11529 31263
rect 11563 31229 11575 31263
rect 11698 31260 11704 31272
rect 11659 31232 11704 31260
rect 11517 31223 11575 31229
rect 11698 31220 11704 31232
rect 11756 31220 11762 31272
rect 11885 31263 11943 31269
rect 11885 31229 11897 31263
rect 11931 31229 11943 31263
rect 11885 31223 11943 31229
rect 12069 31263 12127 31269
rect 12069 31229 12081 31263
rect 12115 31260 12127 31263
rect 12434 31260 12440 31272
rect 12115 31232 12440 31260
rect 12115 31229 12127 31232
rect 12069 31223 12127 31229
rect 11900 31192 11928 31223
rect 12434 31220 12440 31232
rect 12492 31260 12498 31272
rect 12618 31260 12624 31272
rect 12492 31232 12624 31260
rect 12492 31220 12498 31232
rect 12618 31220 12624 31232
rect 12676 31220 12682 31272
rect 13004 31204 13032 31436
rect 13170 31424 13176 31436
rect 13228 31424 13234 31476
rect 16945 31467 17003 31473
rect 16945 31433 16957 31467
rect 16991 31464 17003 31467
rect 16991 31436 17080 31464
rect 16991 31433 17003 31436
rect 16945 31427 17003 31433
rect 16577 31399 16635 31405
rect 16577 31365 16589 31399
rect 16623 31396 16635 31399
rect 16758 31396 16764 31408
rect 16623 31368 16764 31396
rect 16623 31365 16635 31368
rect 16577 31359 16635 31365
rect 16758 31356 16764 31368
rect 16816 31356 16822 31408
rect 14274 31220 14280 31272
rect 14332 31260 14338 31272
rect 14829 31263 14887 31269
rect 14829 31260 14841 31263
rect 14332 31232 14841 31260
rect 14332 31220 14338 31232
rect 14829 31229 14841 31232
rect 14875 31229 14887 31263
rect 15102 31260 15108 31272
rect 15063 31232 15108 31260
rect 14829 31223 14887 31229
rect 11440 31164 11928 31192
rect 11333 31155 11391 31161
rect 12986 31152 12992 31204
rect 13044 31192 13050 31204
rect 14734 31192 14740 31204
rect 13044 31164 14740 31192
rect 13044 31152 13050 31164
rect 14734 31152 14740 31164
rect 14792 31152 14798 31204
rect 14844 31192 14872 31223
rect 15102 31220 15108 31232
rect 15160 31220 15166 31272
rect 17052 31260 17080 31436
rect 20162 31424 20168 31476
rect 20220 31464 20226 31476
rect 21545 31467 21603 31473
rect 21545 31464 21557 31467
rect 20220 31436 21557 31464
rect 20220 31424 20226 31436
rect 21545 31433 21557 31436
rect 21591 31433 21603 31467
rect 21545 31427 21603 31433
rect 21634 31424 21640 31476
rect 21692 31464 21698 31476
rect 24854 31464 24860 31476
rect 21692 31436 24860 31464
rect 21692 31424 21698 31436
rect 24854 31424 24860 31436
rect 24912 31424 24918 31476
rect 24946 31424 24952 31476
rect 25004 31464 25010 31476
rect 26329 31467 26387 31473
rect 26329 31464 26341 31467
rect 25004 31436 26341 31464
rect 25004 31424 25010 31436
rect 26329 31433 26341 31436
rect 26375 31433 26387 31467
rect 26329 31427 26387 31433
rect 27614 31424 27620 31476
rect 27672 31464 27678 31476
rect 28721 31467 28779 31473
rect 28721 31464 28733 31467
rect 27672 31436 28733 31464
rect 27672 31424 27678 31436
rect 28721 31433 28733 31436
rect 28767 31433 28779 31467
rect 28721 31427 28779 31433
rect 30745 31467 30803 31473
rect 30745 31433 30757 31467
rect 30791 31464 30803 31467
rect 30834 31464 30840 31476
rect 30791 31436 30840 31464
rect 30791 31433 30803 31436
rect 30745 31427 30803 31433
rect 30834 31424 30840 31436
rect 30892 31424 30898 31476
rect 17129 31399 17187 31405
rect 17129 31365 17141 31399
rect 17175 31365 17187 31399
rect 23382 31396 23388 31408
rect 23343 31368 23388 31396
rect 17129 31359 17187 31365
rect 17144 31328 17172 31359
rect 23382 31356 23388 31368
rect 23440 31356 23446 31408
rect 23934 31356 23940 31408
rect 23992 31396 23998 31408
rect 29549 31399 29607 31405
rect 29549 31396 29561 31399
rect 23992 31368 29561 31396
rect 23992 31356 23998 31368
rect 29549 31365 29561 31368
rect 29595 31365 29607 31399
rect 29549 31359 29607 31365
rect 18693 31331 18751 31337
rect 17144 31300 18000 31328
rect 17494 31260 17500 31272
rect 17052 31232 17500 31260
rect 17494 31220 17500 31232
rect 17552 31260 17558 31272
rect 17678 31260 17684 31272
rect 17552 31232 17684 31260
rect 17552 31220 17558 31232
rect 17678 31220 17684 31232
rect 17736 31220 17742 31272
rect 17773 31263 17831 31269
rect 17773 31229 17785 31263
rect 17819 31260 17831 31263
rect 17862 31260 17868 31272
rect 17819 31232 17868 31260
rect 17819 31229 17831 31232
rect 17773 31223 17831 31229
rect 17862 31220 17868 31232
rect 17920 31220 17926 31272
rect 17972 31269 18000 31300
rect 18693 31297 18705 31331
rect 18739 31328 18751 31331
rect 18874 31328 18880 31340
rect 18739 31300 18880 31328
rect 18739 31297 18751 31300
rect 18693 31291 18751 31297
rect 18874 31288 18880 31300
rect 18932 31288 18938 31340
rect 19242 31288 19248 31340
rect 19300 31328 19306 31340
rect 20165 31331 20223 31337
rect 20165 31328 20177 31331
rect 19300 31300 20177 31328
rect 19300 31288 19306 31300
rect 20165 31297 20177 31300
rect 20211 31297 20223 31331
rect 20165 31291 20223 31297
rect 17957 31263 18015 31269
rect 17957 31229 17969 31263
rect 18003 31229 18015 31263
rect 17957 31223 18015 31229
rect 18138 31220 18144 31272
rect 18196 31260 18202 31272
rect 18417 31263 18475 31269
rect 18417 31260 18429 31263
rect 18196 31232 18429 31260
rect 18196 31220 18202 31232
rect 18417 31229 18429 31232
rect 18463 31260 18475 31263
rect 18506 31260 18512 31272
rect 18463 31232 18512 31260
rect 18463 31229 18475 31232
rect 18417 31223 18475 31229
rect 18506 31220 18512 31232
rect 18564 31260 18570 31272
rect 19702 31260 19708 31272
rect 18564 31232 19334 31260
rect 19663 31232 19708 31260
rect 18564 31220 18570 31232
rect 18966 31192 18972 31204
rect 14844 31164 18972 31192
rect 18966 31152 18972 31164
rect 19024 31152 19030 31204
rect 3602 31124 3608 31136
rect 3160 31096 3608 31124
rect 3602 31084 3608 31096
rect 3660 31084 3666 31136
rect 6365 31127 6423 31133
rect 6365 31093 6377 31127
rect 6411 31124 6423 31127
rect 6454 31124 6460 31136
rect 6411 31096 6460 31124
rect 6411 31093 6423 31096
rect 6365 31087 6423 31093
rect 6454 31084 6460 31096
rect 6512 31084 6518 31136
rect 6730 31084 6736 31136
rect 6788 31124 6794 31136
rect 8294 31124 8300 31136
rect 6788 31096 8300 31124
rect 6788 31084 6794 31096
rect 8294 31084 8300 31096
rect 8352 31084 8358 31136
rect 11606 31084 11612 31136
rect 11664 31124 11670 31136
rect 12342 31124 12348 31136
rect 11664 31096 12348 31124
rect 11664 31084 11670 31096
rect 12342 31084 12348 31096
rect 12400 31084 12406 31136
rect 13170 31084 13176 31136
rect 13228 31124 13234 31136
rect 13538 31124 13544 31136
rect 13228 31096 13544 31124
rect 13228 31084 13234 31096
rect 13538 31084 13544 31096
rect 13596 31084 13602 31136
rect 14366 31124 14372 31136
rect 14279 31096 14372 31124
rect 14366 31084 14372 31096
rect 14424 31124 14430 31136
rect 16942 31124 16948 31136
rect 14424 31096 16948 31124
rect 14424 31084 14430 31096
rect 16942 31084 16948 31096
rect 17000 31084 17006 31136
rect 17310 31084 17316 31136
rect 17368 31124 17374 31136
rect 17494 31124 17500 31136
rect 17368 31096 17500 31124
rect 17368 31084 17374 31096
rect 17494 31084 17500 31096
rect 17552 31084 17558 31136
rect 19306 31124 19334 31232
rect 19702 31220 19708 31232
rect 19760 31220 19766 31272
rect 20438 31269 20444 31272
rect 20432 31260 20444 31269
rect 20399 31232 20444 31260
rect 20432 31223 20444 31232
rect 20438 31220 20444 31223
rect 20496 31220 20502 31272
rect 22002 31260 22008 31272
rect 21560 31232 21772 31260
rect 21963 31232 22008 31260
rect 19613 31195 19671 31201
rect 19613 31161 19625 31195
rect 19659 31192 19671 31195
rect 21560 31192 21588 31232
rect 19659 31164 21588 31192
rect 19659 31161 19671 31164
rect 19613 31155 19671 31161
rect 21634 31152 21640 31204
rect 21692 31152 21698 31204
rect 21744 31192 21772 31232
rect 22002 31220 22008 31232
rect 22060 31220 22066 31272
rect 22278 31269 22284 31272
rect 22272 31223 22284 31269
rect 22336 31260 22342 31272
rect 22336 31232 22372 31260
rect 22278 31220 22284 31223
rect 22336 31220 22342 31232
rect 22738 31220 22744 31272
rect 22796 31260 22802 31272
rect 23400 31260 23428 31356
rect 24946 31328 24952 31340
rect 24907 31300 24952 31328
rect 24946 31288 24952 31300
rect 25004 31288 25010 31340
rect 25041 31331 25099 31337
rect 25041 31297 25053 31331
rect 25087 31328 25099 31331
rect 25590 31328 25596 31340
rect 25087 31300 25596 31328
rect 25087 31297 25099 31300
rect 25041 31291 25099 31297
rect 25590 31288 25596 31300
rect 25648 31288 25654 31340
rect 26326 31328 26332 31340
rect 25700 31300 26332 31328
rect 22796 31232 23428 31260
rect 24765 31263 24823 31269
rect 22796 31220 22802 31232
rect 24765 31229 24777 31263
rect 24811 31229 24823 31263
rect 24765 31223 24823 31229
rect 25133 31263 25191 31269
rect 25133 31229 25145 31263
rect 25179 31229 25191 31263
rect 25133 31223 25191 31229
rect 25317 31263 25375 31269
rect 25317 31229 25329 31263
rect 25363 31260 25375 31263
rect 25406 31260 25412 31272
rect 25363 31232 25412 31260
rect 25363 31229 25375 31232
rect 25317 31223 25375 31229
rect 23382 31192 23388 31204
rect 21744 31164 23388 31192
rect 23382 31152 23388 31164
rect 23440 31152 23446 31204
rect 24780 31192 24808 31223
rect 25038 31192 25044 31204
rect 24780 31164 25044 31192
rect 25038 31152 25044 31164
rect 25096 31152 25102 31204
rect 25148 31192 25176 31223
rect 25406 31220 25412 31232
rect 25464 31220 25470 31272
rect 25498 31220 25504 31272
rect 25556 31260 25562 31272
rect 25700 31260 25728 31300
rect 26326 31288 26332 31300
rect 26384 31288 26390 31340
rect 26697 31331 26755 31337
rect 26697 31297 26709 31331
rect 26743 31328 26755 31331
rect 27338 31328 27344 31340
rect 26743 31300 27344 31328
rect 26743 31297 26755 31300
rect 26697 31291 26755 31297
rect 27338 31288 27344 31300
rect 27396 31288 27402 31340
rect 27522 31288 27528 31340
rect 27580 31328 27586 31340
rect 28169 31331 28227 31337
rect 28169 31328 28181 31331
rect 27580 31300 28181 31328
rect 27580 31288 27586 31300
rect 28169 31297 28181 31300
rect 28215 31328 28227 31331
rect 28258 31328 28264 31340
rect 28215 31300 28264 31328
rect 28215 31297 28227 31300
rect 28169 31291 28227 31297
rect 28258 31288 28264 31300
rect 28316 31288 28322 31340
rect 25556 31232 25728 31260
rect 25556 31220 25562 31232
rect 26142 31220 26148 31272
rect 26200 31260 26206 31272
rect 26421 31263 26479 31269
rect 26421 31260 26433 31263
rect 26200 31232 26433 31260
rect 26200 31220 26206 31232
rect 26421 31229 26433 31232
rect 26467 31229 26479 31263
rect 26602 31260 26608 31272
rect 26563 31232 26608 31260
rect 26421 31223 26479 31229
rect 26602 31220 26608 31232
rect 26660 31220 26666 31272
rect 26789 31263 26847 31269
rect 26789 31229 26801 31263
rect 26835 31229 26847 31263
rect 26789 31223 26847 31229
rect 26973 31263 27031 31269
rect 26973 31229 26985 31263
rect 27019 31260 27031 31263
rect 27246 31260 27252 31272
rect 27019 31232 27252 31260
rect 27019 31229 27031 31232
rect 26973 31223 27031 31229
rect 25148 31164 25544 31192
rect 21652 31124 21680 31152
rect 25516 31136 25544 31164
rect 25590 31152 25596 31204
rect 25648 31192 25654 31204
rect 26234 31192 26240 31204
rect 25648 31164 26240 31192
rect 25648 31152 25654 31164
rect 26234 31152 26240 31164
rect 26292 31152 26298 31204
rect 26329 31195 26387 31201
rect 26329 31161 26341 31195
rect 26375 31192 26387 31195
rect 26804 31192 26832 31223
rect 27246 31220 27252 31232
rect 27304 31260 27310 31272
rect 28074 31260 28080 31272
rect 27304 31232 28080 31260
rect 27304 31220 27310 31232
rect 28074 31220 28080 31232
rect 28132 31220 28138 31272
rect 27430 31192 27436 31204
rect 26375 31164 27436 31192
rect 26375 31161 26387 31164
rect 26329 31155 26387 31161
rect 27430 31152 27436 31164
rect 27488 31152 27494 31204
rect 19306 31096 21680 31124
rect 22278 31084 22284 31136
rect 22336 31124 22342 31136
rect 22646 31124 22652 31136
rect 22336 31096 22652 31124
rect 22336 31084 22342 31096
rect 22646 31084 22652 31096
rect 22704 31084 22710 31136
rect 24578 31124 24584 31136
rect 24539 31096 24584 31124
rect 24578 31084 24584 31096
rect 24636 31084 24642 31136
rect 25498 31084 25504 31136
rect 25556 31124 25562 31136
rect 25777 31127 25835 31133
rect 25777 31124 25789 31127
rect 25556 31096 25789 31124
rect 25556 31084 25562 31096
rect 25777 31093 25789 31096
rect 25823 31093 25835 31127
rect 25777 31087 25835 31093
rect 27062 31084 27068 31136
rect 27120 31124 27126 31136
rect 27157 31127 27215 31133
rect 27157 31124 27169 31127
rect 27120 31096 27169 31124
rect 27120 31084 27126 31096
rect 27157 31093 27169 31096
rect 27203 31093 27215 31127
rect 27614 31124 27620 31136
rect 27575 31096 27620 31124
rect 27157 31087 27215 31093
rect 27614 31084 27620 31096
rect 27672 31084 27678 31136
rect 30190 31124 30196 31136
rect 30151 31096 30196 31124
rect 30190 31084 30196 31096
rect 30248 31084 30254 31136
rect 31018 31084 31024 31136
rect 31076 31124 31082 31136
rect 31205 31127 31263 31133
rect 31205 31124 31217 31127
rect 31076 31096 31217 31124
rect 31076 31084 31082 31096
rect 31205 31093 31217 31096
rect 31251 31093 31263 31127
rect 31205 31087 31263 31093
rect 1104 31034 32016 31056
rect 1104 30982 11253 31034
rect 11305 30982 11317 31034
rect 11369 30982 11381 31034
rect 11433 30982 11445 31034
rect 11497 30982 11509 31034
rect 11561 30982 21557 31034
rect 21609 30982 21621 31034
rect 21673 30982 21685 31034
rect 21737 30982 21749 31034
rect 21801 30982 21813 31034
rect 21865 30982 32016 31034
rect 1104 30960 32016 30982
rect 2130 30880 2136 30932
rect 2188 30920 2194 30932
rect 2593 30923 2651 30929
rect 2593 30920 2605 30923
rect 2188 30892 2605 30920
rect 2188 30880 2194 30892
rect 2593 30889 2605 30892
rect 2639 30889 2651 30923
rect 3786 30920 3792 30932
rect 3747 30892 3792 30920
rect 2593 30883 2651 30889
rect 3786 30880 3792 30892
rect 3844 30880 3850 30932
rect 5074 30920 5080 30932
rect 5035 30892 5080 30920
rect 5074 30880 5080 30892
rect 5132 30880 5138 30932
rect 6917 30923 6975 30929
rect 6917 30889 6929 30923
rect 6963 30920 6975 30923
rect 7282 30920 7288 30932
rect 6963 30892 7288 30920
rect 6963 30889 6975 30892
rect 6917 30883 6975 30889
rect 7282 30880 7288 30892
rect 7340 30920 7346 30932
rect 7742 30920 7748 30932
rect 7340 30892 7748 30920
rect 7340 30880 7346 30892
rect 7742 30880 7748 30892
rect 7800 30880 7806 30932
rect 8202 30880 8208 30932
rect 8260 30920 8266 30932
rect 8849 30923 8907 30929
rect 8849 30920 8861 30923
rect 8260 30892 8861 30920
rect 8260 30880 8266 30892
rect 8849 30889 8861 30892
rect 8895 30889 8907 30923
rect 8849 30883 8907 30889
rect 8938 30880 8944 30932
rect 8996 30920 9002 30932
rect 9309 30923 9367 30929
rect 9309 30920 9321 30923
rect 8996 30892 9321 30920
rect 8996 30880 9002 30892
rect 9309 30889 9321 30892
rect 9355 30889 9367 30923
rect 9309 30883 9367 30889
rect 10965 30923 11023 30929
rect 10965 30889 10977 30923
rect 11011 30920 11023 30923
rect 14366 30920 14372 30932
rect 11011 30892 14372 30920
rect 11011 30889 11023 30892
rect 10965 30883 11023 30889
rect 14366 30880 14372 30892
rect 14424 30880 14430 30932
rect 16117 30923 16175 30929
rect 16117 30889 16129 30923
rect 16163 30920 16175 30923
rect 16298 30920 16304 30932
rect 16163 30892 16304 30920
rect 16163 30889 16175 30892
rect 16117 30883 16175 30889
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 18046 30920 18052 30932
rect 16684 30892 18052 30920
rect 2038 30852 2044 30864
rect 1999 30824 2044 30852
rect 2038 30812 2044 30824
rect 2096 30812 2102 30864
rect 4430 30852 4436 30864
rect 3160 30824 4436 30852
rect 1762 30744 1768 30796
rect 1820 30784 1826 30796
rect 1857 30787 1915 30793
rect 1857 30784 1869 30787
rect 1820 30756 1869 30784
rect 1820 30744 1826 30756
rect 1857 30753 1869 30756
rect 1903 30753 1915 30787
rect 1857 30747 1915 30753
rect 2406 30744 2412 30796
rect 2464 30784 2470 30796
rect 3160 30793 3188 30824
rect 4430 30812 4436 30824
rect 4488 30852 4494 30864
rect 4488 30824 5580 30852
rect 4488 30812 4494 30824
rect 2685 30787 2743 30793
rect 2685 30784 2697 30787
rect 2464 30756 2697 30784
rect 2464 30744 2470 30756
rect 2685 30753 2697 30756
rect 2731 30753 2743 30787
rect 2685 30747 2743 30753
rect 3145 30787 3203 30793
rect 3145 30753 3157 30787
rect 3191 30753 3203 30787
rect 3326 30784 3332 30796
rect 3287 30756 3332 30784
rect 3145 30747 3203 30753
rect 3326 30744 3332 30756
rect 3384 30744 3390 30796
rect 3421 30787 3479 30793
rect 3421 30753 3433 30787
rect 3467 30753 3479 30787
rect 3421 30747 3479 30753
rect 2314 30676 2320 30728
rect 2372 30716 2378 30728
rect 3436 30716 3464 30747
rect 3510 30744 3516 30796
rect 3568 30784 3574 30796
rect 4062 30784 4068 30796
rect 3568 30756 4068 30784
rect 3568 30744 3574 30756
rect 4062 30744 4068 30756
rect 4120 30744 4126 30796
rect 4154 30744 4160 30796
rect 4212 30784 4218 30796
rect 4338 30784 4344 30796
rect 4212 30756 4344 30784
rect 4212 30744 4218 30756
rect 4338 30744 4344 30756
rect 4396 30784 4402 30796
rect 4525 30787 4583 30793
rect 4525 30784 4537 30787
rect 4396 30756 4537 30784
rect 4396 30744 4402 30756
rect 4525 30753 4537 30756
rect 4571 30753 4583 30787
rect 4982 30784 4988 30796
rect 4943 30756 4988 30784
rect 4525 30747 4583 30753
rect 4982 30744 4988 30756
rect 5040 30744 5046 30796
rect 5552 30793 5580 30824
rect 7374 30812 7380 30864
rect 7432 30852 7438 30864
rect 9861 30855 9919 30861
rect 9861 30852 9873 30855
rect 7432 30824 9873 30852
rect 7432 30812 7438 30824
rect 9861 30821 9873 30824
rect 9907 30821 9919 30855
rect 9861 30815 9919 30821
rect 13814 30812 13820 30864
rect 13872 30852 13878 30864
rect 14458 30852 14464 30864
rect 13872 30824 14464 30852
rect 13872 30812 13878 30824
rect 14458 30812 14464 30824
rect 14516 30812 14522 30864
rect 15010 30861 15016 30864
rect 15004 30852 15016 30861
rect 14971 30824 15016 30852
rect 15004 30815 15016 30824
rect 15010 30812 15016 30815
rect 15068 30812 15074 30864
rect 5537 30787 5595 30793
rect 5537 30753 5549 30787
rect 5583 30753 5595 30787
rect 5718 30784 5724 30796
rect 5679 30756 5724 30784
rect 5537 30747 5595 30753
rect 5718 30744 5724 30756
rect 5776 30744 5782 30796
rect 6546 30744 6552 30796
rect 6604 30784 6610 30796
rect 6733 30787 6791 30793
rect 6733 30784 6745 30787
rect 6604 30756 6745 30784
rect 6604 30744 6610 30756
rect 6733 30753 6745 30756
rect 6779 30753 6791 30787
rect 6733 30747 6791 30753
rect 7736 30787 7794 30793
rect 7736 30753 7748 30787
rect 7782 30784 7794 30787
rect 8018 30784 8024 30796
rect 7782 30756 8024 30784
rect 7782 30753 7794 30756
rect 7736 30747 7794 30753
rect 8018 30744 8024 30756
rect 8076 30744 8082 30796
rect 11698 30744 11704 30796
rect 11756 30784 11762 30796
rect 12342 30784 12348 30796
rect 11756 30756 12348 30784
rect 11756 30744 11762 30756
rect 12342 30744 12348 30756
rect 12400 30784 12406 30796
rect 14001 30787 14059 30793
rect 14001 30784 14013 30787
rect 12400 30756 14013 30784
rect 12400 30744 12406 30756
rect 14001 30753 14013 30756
rect 14047 30753 14059 30787
rect 14001 30747 14059 30753
rect 14090 30744 14096 30796
rect 14148 30784 14154 30796
rect 14734 30784 14740 30796
rect 14148 30756 14740 30784
rect 14148 30744 14154 30756
rect 14734 30744 14740 30756
rect 14792 30744 14798 30796
rect 16684 30784 16712 30892
rect 18046 30880 18052 30892
rect 18104 30880 18110 30932
rect 22554 30920 22560 30932
rect 22515 30892 22560 30920
rect 22554 30880 22560 30892
rect 22612 30880 22618 30932
rect 23017 30923 23075 30929
rect 23017 30889 23029 30923
rect 23063 30889 23075 30923
rect 27614 30920 27620 30932
rect 23017 30883 23075 30889
rect 24780 30892 27620 30920
rect 16758 30812 16764 30864
rect 16816 30852 16822 30864
rect 18138 30852 18144 30864
rect 16816 30824 18144 30852
rect 16816 30812 16822 30824
rect 17236 30793 17264 30824
rect 18138 30812 18144 30824
rect 18196 30812 18202 30864
rect 18233 30855 18291 30861
rect 18233 30821 18245 30855
rect 18279 30852 18291 30855
rect 19150 30852 19156 30864
rect 18279 30824 19156 30852
rect 18279 30821 18291 30824
rect 18233 30815 18291 30821
rect 19150 30812 19156 30824
rect 19208 30852 19214 30864
rect 21174 30852 21180 30864
rect 19208 30824 21180 30852
rect 19208 30812 19214 30824
rect 21174 30812 21180 30824
rect 21232 30812 21238 30864
rect 21358 30812 21364 30864
rect 21416 30852 21422 30864
rect 23032 30852 23060 30883
rect 21416 30824 23060 30852
rect 21416 30812 21422 30824
rect 14844 30756 16712 30784
rect 17037 30787 17095 30793
rect 4246 30716 4252 30728
rect 2372 30688 3556 30716
rect 4207 30688 4252 30716
rect 2372 30676 2378 30688
rect 3528 30648 3556 30688
rect 4246 30676 4252 30688
rect 4304 30676 4310 30728
rect 4709 30719 4767 30725
rect 4709 30685 4721 30719
rect 4755 30716 4767 30719
rect 5074 30716 5080 30728
rect 4755 30688 5080 30716
rect 4755 30685 4767 30688
rect 4709 30679 4767 30685
rect 5074 30676 5080 30688
rect 5132 30676 5138 30728
rect 7469 30719 7527 30725
rect 7469 30685 7481 30719
rect 7515 30685 7527 30719
rect 12434 30716 12440 30728
rect 12395 30688 12440 30716
rect 7469 30679 7527 30685
rect 5902 30648 5908 30660
rect 3528 30620 5908 30648
rect 5902 30608 5908 30620
rect 5960 30608 5966 30660
rect 2958 30540 2964 30592
rect 3016 30580 3022 30592
rect 5074 30580 5080 30592
rect 3016 30552 5080 30580
rect 3016 30540 3022 30552
rect 5074 30540 5080 30552
rect 5132 30540 5138 30592
rect 5534 30580 5540 30592
rect 5495 30552 5540 30580
rect 5534 30540 5540 30552
rect 5592 30540 5598 30592
rect 7484 30580 7512 30679
rect 12434 30676 12440 30688
rect 12492 30676 12498 30728
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30716 12771 30719
rect 13814 30716 13820 30728
rect 12759 30688 13820 30716
rect 12759 30685 12771 30688
rect 12713 30679 12771 30685
rect 13814 30676 13820 30688
rect 13872 30676 13878 30728
rect 14274 30716 14280 30728
rect 14235 30688 14280 30716
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 14844 30716 14872 30756
rect 17037 30753 17049 30787
rect 17083 30753 17095 30787
rect 17037 30747 17095 30753
rect 17221 30787 17279 30793
rect 17221 30753 17233 30787
rect 17267 30753 17279 30787
rect 17221 30747 17279 30753
rect 17589 30787 17647 30793
rect 17589 30753 17601 30787
rect 17635 30784 17647 30787
rect 18046 30784 18052 30796
rect 17635 30756 18052 30784
rect 17635 30753 17647 30756
rect 17589 30747 17647 30753
rect 14752 30688 14872 30716
rect 12452 30648 12480 30676
rect 13078 30648 13084 30660
rect 12452 30620 13084 30648
rect 13078 30608 13084 30620
rect 13136 30608 13142 30660
rect 13538 30608 13544 30660
rect 13596 30648 13602 30660
rect 14752 30648 14780 30688
rect 13596 30620 14780 30648
rect 13596 30608 13602 30620
rect 8386 30580 8392 30592
rect 7484 30552 8392 30580
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 12158 30540 12164 30592
rect 12216 30580 12222 30592
rect 13354 30580 13360 30592
rect 12216 30552 13360 30580
rect 12216 30540 12222 30552
rect 13354 30540 13360 30552
rect 13412 30540 13418 30592
rect 17052 30580 17080 30747
rect 18046 30744 18052 30756
rect 18104 30744 18110 30796
rect 20622 30744 20628 30796
rect 20680 30784 20686 30796
rect 20717 30787 20775 30793
rect 20717 30784 20729 30787
rect 20680 30756 20729 30784
rect 20680 30744 20686 30756
rect 20717 30753 20729 30756
rect 20763 30753 20775 30787
rect 21818 30784 21824 30796
rect 21779 30756 21824 30784
rect 20717 30747 20775 30753
rect 21818 30744 21824 30756
rect 21876 30744 21882 30796
rect 22005 30790 22063 30793
rect 22005 30787 22140 30790
rect 22005 30753 22017 30787
rect 22051 30784 22140 30787
rect 22278 30784 22284 30796
rect 22051 30762 22284 30784
rect 22051 30753 22063 30762
rect 22112 30756 22284 30762
rect 22005 30747 22063 30753
rect 22278 30744 22284 30756
rect 22336 30744 22342 30796
rect 22373 30787 22431 30793
rect 22373 30753 22385 30787
rect 22419 30784 22431 30787
rect 23293 30787 23351 30793
rect 23293 30784 23305 30787
rect 22419 30756 23305 30784
rect 22419 30753 22431 30756
rect 22373 30747 22431 30753
rect 23293 30753 23305 30756
rect 23339 30753 23351 30787
rect 23474 30784 23480 30796
rect 23435 30756 23480 30784
rect 23293 30747 23351 30753
rect 17313 30719 17371 30725
rect 17313 30685 17325 30719
rect 17359 30685 17371 30719
rect 17313 30679 17371 30685
rect 17405 30719 17463 30725
rect 17405 30685 17417 30719
rect 17451 30716 17463 30719
rect 17678 30716 17684 30728
rect 17451 30688 17684 30716
rect 17451 30685 17463 30688
rect 17405 30679 17463 30685
rect 17328 30648 17356 30679
rect 17678 30676 17684 30688
rect 17736 30676 17742 30728
rect 20441 30719 20499 30725
rect 20441 30685 20453 30719
rect 20487 30716 20499 30719
rect 22094 30716 22100 30728
rect 20487 30688 20760 30716
rect 22055 30688 22100 30716
rect 20487 30685 20499 30688
rect 20441 30679 20499 30685
rect 20732 30660 20760 30688
rect 22094 30676 22100 30688
rect 22152 30676 22158 30728
rect 22186 30676 22192 30728
rect 22244 30716 22250 30728
rect 22244 30688 22289 30716
rect 22244 30676 22250 30688
rect 18414 30648 18420 30660
rect 17328 30620 18420 30648
rect 18414 30608 18420 30620
rect 18472 30648 18478 30660
rect 19426 30648 19432 30660
rect 18472 30620 19432 30648
rect 18472 30608 18478 30620
rect 19426 30608 19432 30620
rect 19484 30608 19490 30660
rect 20714 30608 20720 30660
rect 20772 30608 20778 30660
rect 21910 30608 21916 30660
rect 21968 30648 21974 30660
rect 22388 30648 22416 30747
rect 23474 30744 23480 30756
rect 23532 30744 23538 30796
rect 24213 30787 24271 30793
rect 24213 30753 24225 30787
rect 24259 30784 24271 30787
rect 24486 30784 24492 30796
rect 24259 30756 24492 30784
rect 24259 30753 24271 30756
rect 24213 30747 24271 30753
rect 24486 30744 24492 30756
rect 24544 30784 24550 30796
rect 24780 30784 24808 30892
rect 27614 30880 27620 30892
rect 27672 30880 27678 30932
rect 29086 30880 29092 30932
rect 29144 30920 29150 30932
rect 29365 30923 29423 30929
rect 29365 30920 29377 30923
rect 29144 30892 29377 30920
rect 29144 30880 29150 30892
rect 29365 30889 29377 30892
rect 29411 30889 29423 30923
rect 29365 30883 29423 30889
rect 24854 30812 24860 30864
rect 24912 30852 24918 30864
rect 24912 30824 27844 30852
rect 24912 30812 24918 30824
rect 24544 30756 24808 30784
rect 25225 30787 25283 30793
rect 24544 30744 24550 30756
rect 25225 30753 25237 30787
rect 25271 30784 25283 30787
rect 25406 30784 25412 30796
rect 25271 30756 25412 30784
rect 25271 30753 25283 30756
rect 25225 30747 25283 30753
rect 25406 30744 25412 30756
rect 25464 30744 25470 30796
rect 25682 30744 25688 30796
rect 25740 30784 25746 30796
rect 26142 30784 26148 30796
rect 25740 30756 26148 30784
rect 25740 30744 25746 30756
rect 26142 30744 26148 30756
rect 26200 30784 26206 30796
rect 27065 30787 27123 30793
rect 27065 30784 27077 30787
rect 26200 30756 27077 30784
rect 26200 30744 26206 30756
rect 27065 30753 27077 30756
rect 27111 30753 27123 30787
rect 27246 30784 27252 30796
rect 27207 30756 27252 30784
rect 27065 30747 27123 30753
rect 27246 30744 27252 30756
rect 27304 30744 27310 30796
rect 27433 30787 27491 30793
rect 27433 30753 27445 30787
rect 27479 30753 27491 30787
rect 27433 30747 27491 30753
rect 23201 30719 23259 30725
rect 23201 30685 23213 30719
rect 23247 30685 23259 30719
rect 23382 30716 23388 30728
rect 23343 30688 23388 30716
rect 23201 30679 23259 30685
rect 21968 30620 22416 30648
rect 23216 30648 23244 30679
rect 23382 30676 23388 30688
rect 23440 30676 23446 30728
rect 23750 30676 23756 30728
rect 23808 30716 23814 30728
rect 25501 30719 25559 30725
rect 23808 30688 25452 30716
rect 23808 30676 23814 30688
rect 23290 30648 23296 30660
rect 23216 30620 23296 30648
rect 21968 30608 21974 30620
rect 23290 30608 23296 30620
rect 23348 30648 23354 30660
rect 24210 30648 24216 30660
rect 23348 30620 24216 30648
rect 23348 30608 23354 30620
rect 24210 30608 24216 30620
rect 24268 30608 24274 30660
rect 25424 30648 25452 30688
rect 25501 30685 25513 30719
rect 25547 30716 25559 30719
rect 25590 30716 25596 30728
rect 25547 30688 25596 30716
rect 25547 30685 25559 30688
rect 25501 30679 25559 30685
rect 25590 30676 25596 30688
rect 25648 30676 25654 30728
rect 27338 30716 27344 30728
rect 27299 30688 27344 30716
rect 27338 30676 27344 30688
rect 27396 30676 27402 30728
rect 27448 30660 27476 30747
rect 27614 30744 27620 30796
rect 27672 30784 27678 30796
rect 27816 30784 27844 30824
rect 28258 30812 28264 30864
rect 28316 30852 28322 30864
rect 31021 30855 31079 30861
rect 31021 30852 31033 30855
rect 28316 30824 31033 30852
rect 28316 30812 28322 30824
rect 31021 30821 31033 30824
rect 31067 30821 31079 30855
rect 31021 30815 31079 30821
rect 29917 30787 29975 30793
rect 29917 30784 29929 30787
rect 27672 30756 27717 30784
rect 27816 30756 29929 30784
rect 27672 30744 27678 30756
rect 29917 30753 29929 30756
rect 29963 30753 29975 30787
rect 29917 30747 29975 30753
rect 27706 30676 27712 30728
rect 27764 30716 27770 30728
rect 28261 30719 28319 30725
rect 28261 30716 28273 30719
rect 27764 30688 28273 30716
rect 27764 30676 27770 30688
rect 28261 30685 28273 30688
rect 28307 30685 28319 30719
rect 28261 30679 28319 30685
rect 28905 30719 28963 30725
rect 28905 30685 28917 30719
rect 28951 30716 28963 30719
rect 31018 30716 31024 30728
rect 28951 30688 31024 30716
rect 28951 30685 28963 30688
rect 28905 30679 28963 30685
rect 31018 30676 31024 30688
rect 31076 30676 31082 30728
rect 25424 30620 27384 30648
rect 17310 30580 17316 30592
rect 17052 30552 17316 30580
rect 17310 30540 17316 30552
rect 17368 30540 17374 30592
rect 17773 30583 17831 30589
rect 17773 30549 17785 30583
rect 17819 30580 17831 30583
rect 17954 30580 17960 30592
rect 17819 30552 17960 30580
rect 17819 30549 17831 30552
rect 17773 30543 17831 30549
rect 17954 30540 17960 30552
rect 18012 30540 18018 30592
rect 19242 30540 19248 30592
rect 19300 30580 19306 30592
rect 19521 30583 19579 30589
rect 19521 30580 19533 30583
rect 19300 30552 19533 30580
rect 19300 30540 19306 30552
rect 19521 30549 19533 30552
rect 19567 30549 19579 30583
rect 19521 30543 19579 30549
rect 23106 30540 23112 30592
rect 23164 30580 23170 30592
rect 24121 30583 24179 30589
rect 24121 30580 24133 30583
rect 23164 30552 24133 30580
rect 23164 30540 23170 30552
rect 24121 30549 24133 30552
rect 24167 30549 24179 30583
rect 24121 30543 24179 30549
rect 25314 30540 25320 30592
rect 25372 30580 25378 30592
rect 25961 30583 26019 30589
rect 25961 30580 25973 30583
rect 25372 30552 25973 30580
rect 25372 30540 25378 30552
rect 25961 30549 25973 30552
rect 26007 30549 26019 30583
rect 27356 30580 27384 30620
rect 27430 30608 27436 30660
rect 27488 30608 27494 30660
rect 30190 30648 30196 30660
rect 27540 30620 30196 30648
rect 27540 30580 27568 30620
rect 30190 30608 30196 30620
rect 30248 30608 30254 30660
rect 27798 30580 27804 30592
rect 27356 30552 27568 30580
rect 27759 30552 27804 30580
rect 25961 30543 26019 30549
rect 27798 30540 27804 30552
rect 27856 30540 27862 30592
rect 30558 30580 30564 30592
rect 30519 30552 30564 30580
rect 30558 30540 30564 30552
rect 30616 30540 30622 30592
rect 1104 30490 32016 30512
rect 1104 30438 6102 30490
rect 6154 30438 6166 30490
rect 6218 30438 6230 30490
rect 6282 30438 6294 30490
rect 6346 30438 6358 30490
rect 6410 30438 16405 30490
rect 16457 30438 16469 30490
rect 16521 30438 16533 30490
rect 16585 30438 16597 30490
rect 16649 30438 16661 30490
rect 16713 30438 26709 30490
rect 26761 30438 26773 30490
rect 26825 30438 26837 30490
rect 26889 30438 26901 30490
rect 26953 30438 26965 30490
rect 27017 30438 32016 30490
rect 1104 30416 32016 30438
rect 2038 30336 2044 30388
rect 2096 30376 2102 30388
rect 4338 30376 4344 30388
rect 2096 30348 4344 30376
rect 2096 30336 2102 30348
rect 4338 30336 4344 30348
rect 4396 30376 4402 30388
rect 6273 30379 6331 30385
rect 6273 30376 6285 30379
rect 4396 30348 6285 30376
rect 4396 30336 4402 30348
rect 6273 30345 6285 30348
rect 6319 30376 6331 30379
rect 6638 30376 6644 30388
rect 6319 30348 6644 30376
rect 6319 30345 6331 30348
rect 6273 30339 6331 30345
rect 6638 30336 6644 30348
rect 6696 30336 6702 30388
rect 7834 30376 7840 30388
rect 7392 30348 7840 30376
rect 3237 30311 3295 30317
rect 3237 30277 3249 30311
rect 3283 30308 3295 30311
rect 4246 30308 4252 30320
rect 3283 30280 4252 30308
rect 3283 30277 3295 30280
rect 3237 30271 3295 30277
rect 4246 30268 4252 30280
rect 4304 30308 4310 30320
rect 5077 30311 5135 30317
rect 4304 30280 4660 30308
rect 4304 30268 4310 30280
rect 2682 30240 2688 30252
rect 2056 30212 2688 30240
rect 1946 30172 1952 30184
rect 1907 30144 1952 30172
rect 1946 30132 1952 30144
rect 2004 30132 2010 30184
rect 2056 30181 2084 30212
rect 2682 30200 2688 30212
rect 2740 30200 2746 30252
rect 3326 30240 3332 30252
rect 3068 30212 3332 30240
rect 2041 30175 2099 30181
rect 2041 30141 2053 30175
rect 2087 30141 2099 30175
rect 2041 30135 2099 30141
rect 2133 30175 2191 30181
rect 2133 30141 2145 30175
rect 2179 30141 2191 30175
rect 2133 30135 2191 30141
rect 2317 30175 2375 30181
rect 2317 30141 2329 30175
rect 2363 30172 2375 30175
rect 2498 30172 2504 30184
rect 2363 30144 2504 30172
rect 2363 30141 2375 30144
rect 2317 30135 2375 30141
rect 2148 30104 2176 30135
rect 2498 30132 2504 30144
rect 2556 30132 2562 30184
rect 3068 30181 3096 30212
rect 3326 30200 3332 30212
rect 3384 30200 3390 30252
rect 4522 30240 4528 30252
rect 4483 30212 4528 30240
rect 4522 30200 4528 30212
rect 4580 30200 4586 30252
rect 4632 30249 4660 30280
rect 5077 30277 5089 30311
rect 5123 30308 5135 30311
rect 5350 30308 5356 30320
rect 5123 30280 5356 30308
rect 5123 30277 5135 30280
rect 5077 30271 5135 30277
rect 5350 30268 5356 30280
rect 5408 30268 5414 30320
rect 6178 30268 6184 30320
rect 6236 30308 6242 30320
rect 7282 30308 7288 30320
rect 6236 30280 7288 30308
rect 6236 30268 6242 30280
rect 7282 30268 7288 30280
rect 7340 30268 7346 30320
rect 4617 30243 4675 30249
rect 4617 30209 4629 30243
rect 4663 30209 4675 30243
rect 7392 30240 7420 30348
rect 7834 30336 7840 30348
rect 7892 30336 7898 30388
rect 8018 30376 8024 30388
rect 7979 30348 8024 30376
rect 8018 30336 8024 30348
rect 8076 30336 8082 30388
rect 8662 30336 8668 30388
rect 8720 30376 8726 30388
rect 8941 30379 8999 30385
rect 8941 30376 8953 30379
rect 8720 30348 8953 30376
rect 8720 30336 8726 30348
rect 8941 30345 8953 30348
rect 8987 30345 8999 30379
rect 8941 30339 8999 30345
rect 12434 30336 12440 30388
rect 12492 30376 12498 30388
rect 12894 30376 12900 30388
rect 12492 30348 12900 30376
rect 12492 30336 12498 30348
rect 12894 30336 12900 30348
rect 12952 30336 12958 30388
rect 13354 30336 13360 30388
rect 13412 30376 13418 30388
rect 16255 30379 16313 30385
rect 16255 30376 16267 30379
rect 13412 30348 16267 30376
rect 13412 30336 13418 30348
rect 16255 30345 16267 30348
rect 16301 30345 16313 30379
rect 16255 30339 16313 30345
rect 17586 30336 17592 30388
rect 17644 30376 17650 30388
rect 23106 30376 23112 30388
rect 17644 30348 23112 30376
rect 17644 30336 17650 30348
rect 23106 30336 23112 30348
rect 23164 30336 23170 30388
rect 27706 30376 27712 30388
rect 24044 30348 27712 30376
rect 7466 30268 7472 30320
rect 7524 30268 7530 30320
rect 18693 30311 18751 30317
rect 18693 30277 18705 30311
rect 18739 30308 18751 30311
rect 19058 30308 19064 30320
rect 18739 30280 19064 30308
rect 18739 30277 18751 30280
rect 18693 30271 18751 30277
rect 19058 30268 19064 30280
rect 19116 30308 19122 30320
rect 19978 30308 19984 30320
rect 19116 30280 19984 30308
rect 19116 30268 19122 30280
rect 19978 30268 19984 30280
rect 20036 30268 20042 30320
rect 20070 30268 20076 30320
rect 20128 30308 20134 30320
rect 20128 30280 22764 30308
rect 20128 30268 20134 30280
rect 4617 30203 4675 30209
rect 4715 30212 7420 30240
rect 7484 30240 7512 30268
rect 7561 30243 7619 30249
rect 7561 30240 7573 30243
rect 7484 30212 7573 30240
rect 3053 30175 3111 30181
rect 3053 30141 3065 30175
rect 3099 30141 3111 30175
rect 3053 30135 3111 30141
rect 3237 30175 3295 30181
rect 3237 30141 3249 30175
rect 3283 30172 3295 30175
rect 3510 30172 3516 30184
rect 3283 30144 3516 30172
rect 3283 30141 3295 30144
rect 3237 30135 3295 30141
rect 3510 30132 3516 30144
rect 3568 30132 3574 30184
rect 3786 30132 3792 30184
rect 3844 30172 3850 30184
rect 4715 30172 4743 30212
rect 7561 30209 7573 30212
rect 7607 30209 7619 30243
rect 7561 30203 7619 30209
rect 7653 30243 7711 30249
rect 7653 30209 7665 30243
rect 7699 30240 7711 30243
rect 7926 30240 7932 30252
rect 7699 30212 7932 30240
rect 7699 30209 7711 30212
rect 7653 30203 7711 30209
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 12158 30240 12164 30252
rect 10336 30212 12164 30240
rect 5534 30172 5540 30184
rect 3844 30144 4743 30172
rect 4816 30144 5540 30172
rect 3844 30132 3850 30144
rect 4709 30107 4767 30113
rect 2148 30076 4476 30104
rect 1670 30036 1676 30048
rect 1631 30008 1676 30036
rect 1670 29996 1676 30008
rect 1728 29996 1734 30048
rect 3881 30039 3939 30045
rect 3881 30005 3893 30039
rect 3927 30036 3939 30039
rect 4154 30036 4160 30048
rect 3927 30008 4160 30036
rect 3927 30005 3939 30008
rect 3881 29999 3939 30005
rect 4154 29996 4160 30008
rect 4212 29996 4218 30048
rect 4448 30036 4476 30076
rect 4709 30073 4721 30107
rect 4755 30104 4767 30107
rect 4816 30104 4844 30144
rect 5534 30132 5540 30144
rect 5592 30132 5598 30184
rect 5629 30175 5687 30181
rect 5629 30141 5641 30175
rect 5675 30172 5687 30175
rect 7006 30172 7012 30184
rect 5675 30144 7012 30172
rect 5675 30141 5687 30144
rect 5629 30135 5687 30141
rect 7006 30132 7012 30144
rect 7064 30132 7070 30184
rect 7098 30132 7104 30184
rect 7156 30172 7162 30184
rect 7285 30175 7343 30181
rect 7285 30172 7297 30175
rect 7156 30144 7297 30172
rect 7156 30132 7162 30144
rect 7285 30141 7297 30144
rect 7331 30141 7343 30175
rect 7285 30135 7343 30141
rect 7469 30175 7527 30181
rect 7469 30141 7481 30175
rect 7515 30141 7527 30175
rect 7469 30135 7527 30141
rect 7837 30175 7895 30181
rect 7837 30141 7849 30175
rect 7883 30172 7895 30175
rect 8202 30172 8208 30184
rect 7883 30144 8208 30172
rect 7883 30141 7895 30144
rect 7837 30135 7895 30141
rect 4755 30076 4844 30104
rect 4755 30073 4767 30076
rect 4709 30067 4767 30073
rect 4890 30064 4896 30116
rect 4948 30104 4954 30116
rect 6270 30113 6276 30116
rect 6241 30107 6276 30113
rect 6241 30104 6253 30107
rect 4948 30076 6253 30104
rect 4948 30064 4954 30076
rect 6241 30073 6253 30076
rect 6241 30067 6276 30073
rect 6270 30064 6276 30067
rect 6328 30064 6334 30116
rect 6454 30104 6460 30116
rect 6415 30076 6460 30104
rect 6454 30064 6460 30076
rect 6512 30064 6518 30116
rect 5258 30036 5264 30048
rect 4448 30008 5264 30036
rect 5258 29996 5264 30008
rect 5316 29996 5322 30048
rect 5350 29996 5356 30048
rect 5408 30036 5414 30048
rect 5718 30036 5724 30048
rect 5408 30008 5724 30036
rect 5408 29996 5414 30008
rect 5718 29996 5724 30008
rect 5776 29996 5782 30048
rect 6086 30036 6092 30048
rect 6047 30008 6092 30036
rect 6086 29996 6092 30008
rect 6144 29996 6150 30048
rect 7300 30036 7328 30135
rect 7484 30104 7512 30135
rect 8202 30132 8208 30144
rect 8260 30132 8266 30184
rect 10336 30181 10364 30212
rect 12158 30200 12164 30212
rect 12216 30200 12222 30252
rect 16025 30243 16083 30249
rect 16025 30209 16037 30243
rect 16071 30240 16083 30243
rect 16574 30240 16580 30252
rect 16071 30212 16580 30240
rect 16071 30209 16083 30212
rect 16025 30203 16083 30209
rect 16574 30200 16580 30212
rect 16632 30200 16638 30252
rect 18966 30200 18972 30252
rect 19024 30240 19030 30252
rect 19705 30243 19763 30249
rect 19705 30240 19717 30243
rect 19024 30212 19717 30240
rect 19024 30200 19030 30212
rect 19705 30209 19717 30212
rect 19751 30209 19763 30243
rect 22186 30240 22192 30252
rect 19705 30203 19763 30209
rect 20364 30212 22192 30240
rect 20364 30184 20392 30212
rect 22186 30200 22192 30212
rect 22244 30240 22250 30252
rect 22649 30243 22707 30249
rect 22649 30240 22661 30243
rect 22244 30212 22661 30240
rect 22244 30200 22250 30212
rect 22649 30209 22661 30212
rect 22695 30209 22707 30243
rect 22736 30240 22764 30280
rect 23198 30268 23204 30320
rect 23256 30308 23262 30320
rect 23934 30308 23940 30320
rect 23256 30280 23940 30308
rect 23256 30268 23262 30280
rect 23934 30268 23940 30280
rect 23992 30268 23998 30320
rect 24044 30240 24072 30348
rect 27706 30336 27712 30348
rect 27764 30336 27770 30388
rect 27908 30348 28212 30376
rect 24210 30268 24216 30320
rect 24268 30308 24274 30320
rect 24762 30308 24768 30320
rect 24268 30280 24768 30308
rect 24268 30268 24274 30280
rect 24762 30268 24768 30280
rect 24820 30268 24826 30320
rect 24949 30311 25007 30317
rect 24949 30277 24961 30311
rect 24995 30308 25007 30311
rect 25590 30308 25596 30320
rect 24995 30280 25596 30308
rect 24995 30277 25007 30280
rect 24949 30271 25007 30277
rect 25590 30268 25596 30280
rect 25648 30268 25654 30320
rect 22736 30212 24072 30240
rect 22649 30203 22707 30209
rect 10321 30175 10379 30181
rect 10321 30172 10333 30175
rect 9416 30144 10333 30172
rect 9416 30116 9444 30144
rect 10321 30141 10333 30144
rect 10367 30141 10379 30175
rect 10321 30135 10379 30141
rect 11146 30132 11152 30184
rect 11204 30172 11210 30184
rect 11333 30175 11391 30181
rect 11333 30172 11345 30175
rect 11204 30144 11345 30172
rect 11204 30132 11210 30144
rect 11333 30141 11345 30144
rect 11379 30141 11391 30175
rect 12894 30172 12900 30184
rect 11333 30135 11391 30141
rect 11440 30144 12900 30172
rect 8662 30104 8668 30116
rect 7484 30076 8668 30104
rect 8662 30064 8668 30076
rect 8720 30064 8726 30116
rect 9398 30064 9404 30116
rect 9456 30064 9462 30116
rect 9490 30064 9496 30116
rect 9548 30104 9554 30116
rect 10054 30107 10112 30113
rect 10054 30104 10066 30107
rect 9548 30076 10066 30104
rect 9548 30064 9554 30076
rect 10054 30073 10066 30076
rect 10100 30073 10112 30107
rect 10054 30067 10112 30073
rect 10502 30064 10508 30116
rect 10560 30104 10566 30116
rect 11440 30104 11468 30144
rect 12894 30132 12900 30144
rect 12952 30132 12958 30184
rect 14734 30132 14740 30184
rect 14792 30172 14798 30184
rect 15565 30175 15623 30181
rect 15565 30172 15577 30175
rect 14792 30144 15577 30172
rect 14792 30132 14798 30144
rect 15565 30141 15577 30144
rect 15611 30141 15623 30175
rect 15565 30135 15623 30141
rect 16666 30132 16672 30184
rect 16724 30172 16730 30184
rect 17313 30175 17371 30181
rect 17313 30172 17325 30175
rect 16724 30144 17325 30172
rect 16724 30132 16730 30144
rect 17313 30141 17325 30144
rect 17359 30172 17371 30175
rect 19242 30172 19248 30184
rect 17359 30144 19248 30172
rect 17359 30141 17371 30144
rect 17313 30135 17371 30141
rect 19242 30132 19248 30144
rect 19300 30132 19306 30184
rect 19981 30175 20039 30181
rect 19981 30141 19993 30175
rect 20027 30172 20039 30175
rect 20346 30172 20352 30184
rect 20027 30144 20352 30172
rect 20027 30141 20039 30144
rect 19981 30135 20039 30141
rect 20346 30132 20352 30144
rect 20404 30132 20410 30184
rect 20714 30132 20720 30184
rect 20772 30172 20778 30184
rect 20993 30175 21051 30181
rect 20993 30172 21005 30175
rect 20772 30144 21005 30172
rect 20772 30132 20778 30144
rect 20993 30141 21005 30144
rect 21039 30141 21051 30175
rect 21266 30172 21272 30184
rect 21227 30144 21272 30172
rect 20993 30135 21051 30141
rect 21266 30132 21272 30144
rect 21324 30172 21330 30184
rect 21818 30172 21824 30184
rect 21324 30144 21824 30172
rect 21324 30132 21330 30144
rect 21818 30132 21824 30144
rect 21876 30172 21882 30184
rect 22281 30175 22339 30181
rect 22281 30172 22293 30175
rect 21876 30144 22293 30172
rect 21876 30132 21882 30144
rect 22281 30141 22293 30144
rect 22327 30141 22339 30175
rect 22462 30172 22468 30184
rect 22423 30144 22468 30172
rect 22281 30135 22339 30141
rect 22462 30132 22468 30144
rect 22520 30132 22526 30184
rect 22557 30175 22615 30181
rect 22557 30141 22569 30175
rect 22603 30141 22615 30175
rect 22557 30135 22615 30141
rect 22833 30175 22891 30181
rect 22833 30141 22845 30175
rect 22879 30172 22891 30175
rect 23290 30172 23296 30184
rect 22879 30144 23296 30172
rect 22879 30141 22891 30144
rect 22833 30135 22891 30141
rect 10560 30076 11468 30104
rect 12428 30107 12486 30113
rect 10560 30064 10566 30076
rect 12428 30073 12440 30107
rect 12474 30104 12486 30107
rect 12526 30104 12532 30116
rect 12474 30076 12532 30104
rect 12474 30073 12486 30076
rect 12428 30067 12486 30073
rect 12526 30064 12532 30076
rect 12584 30064 12590 30116
rect 15010 30064 15016 30116
rect 15068 30104 15074 30116
rect 15298 30107 15356 30113
rect 15298 30104 15310 30107
rect 15068 30076 15310 30104
rect 15068 30064 15074 30076
rect 15298 30073 15310 30076
rect 15344 30073 15356 30107
rect 15298 30067 15356 30073
rect 17580 30107 17638 30113
rect 17580 30073 17592 30107
rect 17626 30104 17638 30107
rect 18598 30104 18604 30116
rect 17626 30076 18604 30104
rect 17626 30073 17638 30076
rect 17580 30067 17638 30073
rect 18598 30064 18604 30076
rect 18656 30064 18662 30116
rect 22572 30104 22600 30135
rect 23290 30132 23296 30144
rect 23348 30132 23354 30184
rect 24765 30175 24823 30181
rect 24765 30141 24777 30175
rect 24811 30172 24823 30175
rect 25314 30172 25320 30184
rect 24811 30144 25320 30172
rect 24811 30141 24823 30144
rect 24765 30135 24823 30141
rect 25314 30132 25320 30144
rect 25372 30132 25378 30184
rect 25409 30175 25467 30181
rect 25409 30141 25421 30175
rect 25455 30141 25467 30175
rect 25682 30172 25688 30184
rect 25643 30144 25688 30172
rect 25409 30135 25467 30141
rect 25424 30104 25452 30135
rect 25682 30132 25688 30144
rect 25740 30132 25746 30184
rect 26142 30132 26148 30184
rect 26200 30172 26206 30184
rect 26697 30175 26755 30181
rect 26697 30172 26709 30175
rect 26200 30144 26709 30172
rect 26200 30132 26206 30144
rect 26697 30141 26709 30144
rect 26743 30141 26755 30175
rect 26697 30135 26755 30141
rect 27338 30132 27344 30184
rect 27396 30172 27402 30184
rect 27908 30172 27936 30348
rect 28074 30308 28080 30320
rect 28035 30280 28080 30308
rect 28074 30268 28080 30280
rect 28132 30268 28138 30320
rect 28184 30308 28212 30348
rect 28629 30311 28687 30317
rect 28629 30308 28641 30311
rect 28184 30280 28641 30308
rect 28629 30277 28641 30280
rect 28675 30277 28687 30311
rect 28629 30271 28687 30277
rect 30374 30268 30380 30320
rect 30432 30308 30438 30320
rect 30650 30308 30656 30320
rect 30432 30280 30656 30308
rect 30432 30268 30438 30280
rect 30650 30268 30656 30280
rect 30708 30308 30714 30320
rect 30837 30311 30895 30317
rect 30837 30308 30849 30311
rect 30708 30280 30849 30308
rect 30708 30268 30714 30280
rect 30837 30277 30849 30280
rect 30883 30277 30895 30311
rect 30837 30271 30895 30277
rect 27396 30144 27936 30172
rect 28092 30172 28120 30268
rect 28442 30200 28448 30252
rect 28500 30240 28506 30252
rect 30558 30240 30564 30252
rect 28500 30212 30564 30240
rect 28500 30200 28506 30212
rect 30558 30200 30564 30212
rect 30616 30200 30622 30252
rect 28537 30175 28595 30181
rect 28537 30172 28549 30175
rect 28092 30144 28549 30172
rect 27396 30132 27402 30144
rect 28537 30141 28549 30144
rect 28583 30141 28595 30175
rect 28537 30135 28595 30141
rect 25590 30104 25596 30116
rect 18708 30076 22600 30104
rect 22949 30076 23612 30104
rect 25424 30076 25596 30104
rect 7558 30036 7564 30048
rect 7300 30008 7564 30036
rect 7558 29996 7564 30008
rect 7616 30036 7622 30048
rect 8110 30036 8116 30048
rect 7616 30008 8116 30036
rect 7616 29996 7622 30008
rect 8110 29996 8116 30008
rect 8168 29996 8174 30048
rect 8294 29996 8300 30048
rect 8352 30036 8358 30048
rect 10781 30039 10839 30045
rect 10781 30036 10793 30039
rect 8352 30008 10793 30036
rect 8352 29996 8358 30008
rect 10781 30005 10793 30008
rect 10827 30005 10839 30039
rect 10781 29999 10839 30005
rect 11425 30039 11483 30045
rect 11425 30005 11437 30039
rect 11471 30036 11483 30039
rect 11882 30036 11888 30048
rect 11471 30008 11888 30036
rect 11471 30005 11483 30008
rect 11425 29999 11483 30005
rect 11882 29996 11888 30008
rect 11940 29996 11946 30048
rect 12710 29996 12716 30048
rect 12768 30036 12774 30048
rect 13446 30036 13452 30048
rect 12768 30008 13452 30036
rect 12768 29996 12774 30008
rect 13446 29996 13452 30008
rect 13504 30036 13510 30048
rect 13541 30039 13599 30045
rect 13541 30036 13553 30039
rect 13504 30008 13553 30036
rect 13504 29996 13510 30008
rect 13541 30005 13553 30008
rect 13587 30005 13599 30039
rect 13541 29999 13599 30005
rect 14185 30039 14243 30045
rect 14185 30005 14197 30039
rect 14231 30036 14243 30039
rect 14826 30036 14832 30048
rect 14231 30008 14832 30036
rect 14231 30005 14243 30008
rect 14185 29999 14243 30005
rect 14826 29996 14832 30008
rect 14884 29996 14890 30048
rect 16114 29996 16120 30048
rect 16172 30036 16178 30048
rect 18708 30036 18736 30076
rect 16172 30008 18736 30036
rect 16172 29996 16178 30008
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 22949 30036 22977 30076
rect 19392 30008 22977 30036
rect 23017 30039 23075 30045
rect 19392 29996 19398 30008
rect 23017 30005 23029 30039
rect 23063 30036 23075 30039
rect 23198 30036 23204 30048
rect 23063 30008 23204 30036
rect 23063 30005 23075 30008
rect 23017 29999 23075 30005
rect 23198 29996 23204 30008
rect 23256 29996 23262 30048
rect 23584 30045 23612 30076
rect 25590 30064 25596 30076
rect 25648 30064 25654 30116
rect 26970 30113 26976 30116
rect 26964 30104 26976 30113
rect 26931 30076 26976 30104
rect 26964 30067 26976 30076
rect 26970 30064 26976 30067
rect 27028 30064 27034 30116
rect 27154 30064 27160 30116
rect 27212 30104 27218 30116
rect 29549 30107 29607 30113
rect 29549 30104 29561 30107
rect 27212 30076 29561 30104
rect 27212 30064 27218 30076
rect 29549 30073 29561 30076
rect 29595 30073 29607 30107
rect 29549 30067 29607 30073
rect 23569 30039 23627 30045
rect 23569 30005 23581 30039
rect 23615 30036 23627 30039
rect 23658 30036 23664 30048
rect 23615 30008 23664 30036
rect 23615 30005 23627 30008
rect 23569 29999 23627 30005
rect 23658 29996 23664 30008
rect 23716 29996 23722 30048
rect 1104 29946 32016 29968
rect 1104 29894 11253 29946
rect 11305 29894 11317 29946
rect 11369 29894 11381 29946
rect 11433 29894 11445 29946
rect 11497 29894 11509 29946
rect 11561 29894 21557 29946
rect 21609 29894 21621 29946
rect 21673 29894 21685 29946
rect 21737 29894 21749 29946
rect 21801 29894 21813 29946
rect 21865 29894 32016 29946
rect 1104 29872 32016 29894
rect 3234 29792 3240 29844
rect 3292 29832 3298 29844
rect 3789 29835 3847 29841
rect 3789 29832 3801 29835
rect 3292 29804 3801 29832
rect 3292 29792 3298 29804
rect 3789 29801 3801 29804
rect 3835 29801 3847 29835
rect 4338 29832 4344 29844
rect 3789 29795 3847 29801
rect 4172 29804 4344 29832
rect 1210 29724 1216 29776
rect 1268 29764 1274 29776
rect 2774 29764 2780 29776
rect 1268 29736 2268 29764
rect 1268 29724 1274 29736
rect 1578 29656 1584 29708
rect 1636 29696 1642 29708
rect 1946 29696 1952 29708
rect 1636 29668 1952 29696
rect 1636 29656 1642 29668
rect 1946 29656 1952 29668
rect 2004 29696 2010 29708
rect 2240 29705 2268 29736
rect 2332 29736 2780 29764
rect 2332 29705 2360 29736
rect 2774 29724 2780 29736
rect 2832 29724 2838 29776
rect 2133 29699 2191 29705
rect 2133 29696 2145 29699
rect 2004 29668 2145 29696
rect 2004 29656 2010 29668
rect 2133 29665 2145 29668
rect 2179 29665 2191 29699
rect 2133 29659 2191 29665
rect 2225 29699 2283 29705
rect 2225 29665 2237 29699
rect 2271 29665 2283 29699
rect 2225 29659 2283 29665
rect 2317 29699 2375 29705
rect 2317 29665 2329 29699
rect 2363 29665 2375 29699
rect 2317 29659 2375 29665
rect 2501 29699 2559 29705
rect 2501 29665 2513 29699
rect 2547 29696 2559 29699
rect 3234 29696 3240 29708
rect 2547 29668 3096 29696
rect 3195 29668 3240 29696
rect 2547 29665 2559 29668
rect 2501 29659 2559 29665
rect 0 29628 800 29642
rect 1762 29628 1768 29640
rect 0 29600 1768 29628
rect 0 29586 800 29600
rect 1762 29588 1768 29600
rect 1820 29588 1826 29640
rect 1946 29520 1952 29572
rect 2004 29560 2010 29572
rect 2332 29560 2360 29659
rect 2961 29631 3019 29637
rect 2961 29628 2973 29631
rect 2004 29532 2360 29560
rect 2746 29600 2973 29628
rect 2004 29520 2010 29532
rect 1857 29495 1915 29501
rect 1857 29461 1869 29495
rect 1903 29492 1915 29495
rect 2746 29492 2774 29600
rect 2961 29597 2973 29600
rect 3007 29597 3019 29631
rect 3068 29628 3096 29668
rect 3234 29656 3240 29668
rect 3292 29656 3298 29708
rect 4062 29696 4068 29708
rect 4023 29668 4068 29696
rect 4062 29656 4068 29668
rect 4120 29656 4126 29708
rect 4172 29705 4200 29804
rect 4338 29792 4344 29804
rect 4396 29792 4402 29844
rect 5537 29835 5595 29841
rect 5537 29801 5549 29835
rect 5583 29801 5595 29835
rect 5537 29795 5595 29801
rect 5350 29764 5356 29776
rect 4264 29736 5356 29764
rect 4264 29708 4292 29736
rect 5350 29724 5356 29736
rect 5408 29724 5414 29776
rect 5552 29764 5580 29795
rect 6270 29792 6276 29844
rect 6328 29832 6334 29844
rect 6733 29835 6791 29841
rect 6733 29832 6745 29835
rect 6328 29804 6745 29832
rect 6328 29792 6334 29804
rect 6733 29801 6745 29804
rect 6779 29801 6791 29835
rect 6733 29795 6791 29801
rect 8297 29835 8355 29841
rect 8297 29801 8309 29835
rect 8343 29832 8355 29835
rect 9490 29832 9496 29844
rect 8343 29804 9496 29832
rect 8343 29801 8355 29804
rect 8297 29795 8355 29801
rect 9490 29792 9496 29804
rect 9548 29792 9554 29844
rect 10318 29792 10324 29844
rect 10376 29832 10382 29844
rect 10594 29832 10600 29844
rect 10376 29804 10600 29832
rect 10376 29792 10382 29804
rect 10594 29792 10600 29804
rect 10652 29792 10658 29844
rect 10781 29835 10839 29841
rect 10781 29801 10793 29835
rect 10827 29832 10839 29835
rect 11146 29832 11152 29844
rect 10827 29804 11152 29832
rect 10827 29801 10839 29804
rect 10781 29795 10839 29801
rect 11146 29792 11152 29804
rect 11204 29792 11210 29844
rect 12621 29835 12679 29841
rect 12621 29832 12633 29835
rect 11716 29804 12633 29832
rect 5902 29764 5908 29776
rect 5552 29736 5908 29764
rect 5902 29724 5908 29736
rect 5960 29724 5966 29776
rect 7834 29724 7840 29776
rect 7892 29764 7898 29776
rect 9582 29764 9588 29776
rect 7892 29736 9588 29764
rect 7892 29724 7898 29736
rect 9582 29724 9588 29736
rect 9640 29764 9646 29776
rect 11716 29764 11744 29804
rect 12621 29801 12633 29804
rect 12667 29832 12679 29835
rect 14550 29832 14556 29844
rect 12667 29804 14556 29832
rect 12667 29801 12679 29804
rect 12621 29795 12679 29801
rect 14550 29792 14556 29804
rect 14608 29792 14614 29844
rect 15933 29835 15991 29841
rect 15933 29801 15945 29835
rect 15979 29832 15991 29835
rect 16114 29832 16120 29844
rect 15979 29804 16120 29832
rect 15979 29801 15991 29804
rect 15933 29795 15991 29801
rect 16114 29792 16120 29804
rect 16172 29792 16178 29844
rect 16942 29792 16948 29844
rect 17000 29832 17006 29844
rect 18049 29835 18107 29841
rect 17000 29804 17632 29832
rect 17000 29792 17006 29804
rect 9640 29736 11744 29764
rect 9640 29724 9646 29736
rect 11790 29724 11796 29776
rect 11848 29764 11854 29776
rect 11977 29767 12035 29773
rect 11977 29764 11989 29767
rect 11848 29736 11989 29764
rect 11848 29724 11854 29736
rect 11977 29733 11989 29736
rect 12023 29733 12035 29767
rect 11977 29727 12035 29733
rect 14274 29724 14280 29776
rect 14332 29764 14338 29776
rect 16025 29767 16083 29773
rect 14332 29736 14872 29764
rect 14332 29724 14338 29736
rect 4157 29699 4215 29705
rect 4157 29665 4169 29699
rect 4203 29665 4215 29699
rect 4157 29659 4215 29665
rect 4246 29656 4252 29708
rect 4304 29696 4310 29708
rect 4433 29699 4491 29705
rect 4304 29668 4397 29696
rect 4304 29656 4310 29668
rect 4433 29665 4445 29699
rect 4479 29665 4491 29699
rect 4433 29659 4491 29665
rect 5445 29699 5503 29705
rect 5445 29665 5457 29699
rect 5491 29665 5503 29699
rect 5445 29659 5503 29665
rect 5813 29699 5871 29705
rect 5813 29665 5825 29699
rect 5859 29696 5871 29699
rect 6086 29696 6092 29708
rect 5859 29668 6092 29696
rect 5859 29665 5871 29668
rect 5813 29659 5871 29665
rect 4338 29628 4344 29640
rect 3068 29600 4344 29628
rect 2961 29591 3019 29597
rect 4338 29588 4344 29600
rect 4396 29588 4402 29640
rect 4062 29520 4068 29572
rect 4120 29560 4126 29572
rect 4448 29560 4476 29659
rect 4120 29532 4476 29560
rect 5460 29560 5488 29659
rect 6086 29656 6092 29668
rect 6144 29656 6150 29708
rect 6546 29696 6552 29708
rect 6472 29668 6552 29696
rect 5629 29631 5687 29637
rect 5629 29597 5641 29631
rect 5675 29628 5687 29631
rect 6178 29628 6184 29640
rect 5675 29600 6184 29628
rect 5675 29597 5687 29600
rect 5629 29591 5687 29597
rect 6178 29588 6184 29600
rect 6236 29588 6242 29640
rect 6472 29637 6500 29668
rect 6546 29656 6552 29668
rect 6604 29656 6610 29708
rect 6641 29699 6699 29705
rect 6641 29665 6653 29699
rect 6687 29696 6699 29699
rect 7558 29696 7564 29708
rect 6687 29668 6776 29696
rect 7519 29668 7564 29696
rect 6687 29665 6699 29668
rect 6641 29659 6699 29665
rect 6457 29631 6515 29637
rect 6457 29597 6469 29631
rect 6503 29597 6515 29631
rect 6457 29591 6515 29597
rect 6748 29572 6776 29668
rect 7558 29656 7564 29668
rect 7616 29656 7622 29708
rect 7650 29656 7656 29708
rect 7708 29696 7714 29708
rect 7745 29699 7803 29705
rect 7745 29696 7757 29699
rect 7708 29668 7757 29696
rect 7708 29656 7714 29668
rect 7745 29665 7757 29668
rect 7791 29665 7803 29699
rect 7745 29659 7803 29665
rect 8113 29699 8171 29705
rect 8113 29665 8125 29699
rect 8159 29696 8171 29699
rect 8662 29696 8668 29708
rect 8159 29668 8668 29696
rect 8159 29665 8171 29668
rect 8113 29659 8171 29665
rect 8662 29656 8668 29668
rect 8720 29656 8726 29708
rect 8757 29699 8815 29705
rect 8757 29665 8769 29699
rect 8803 29665 8815 29699
rect 8757 29659 8815 29665
rect 9668 29699 9726 29705
rect 9668 29665 9680 29699
rect 9714 29696 9726 29699
rect 10502 29696 10508 29708
rect 9714 29668 10508 29696
rect 9714 29665 9726 29668
rect 9668 29659 9726 29665
rect 7466 29588 7472 29640
rect 7524 29628 7530 29640
rect 7837 29631 7895 29637
rect 7837 29628 7849 29631
rect 7524 29600 7849 29628
rect 7524 29588 7530 29600
rect 7837 29597 7849 29600
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 7926 29588 7932 29640
rect 7984 29628 7990 29640
rect 7984 29600 8029 29628
rect 7984 29588 7990 29600
rect 6730 29560 6736 29572
rect 5460 29532 6736 29560
rect 4120 29520 4126 29532
rect 6730 29520 6736 29532
rect 6788 29520 6794 29572
rect 7101 29563 7159 29569
rect 7101 29529 7113 29563
rect 7147 29560 7159 29563
rect 8772 29560 8800 29659
rect 10502 29656 10508 29668
rect 10560 29656 10566 29708
rect 10594 29656 10600 29708
rect 10652 29696 10658 29708
rect 11330 29696 11336 29708
rect 10652 29668 11336 29696
rect 10652 29656 10658 29668
rect 11330 29656 11336 29668
rect 11388 29656 11394 29708
rect 11698 29696 11704 29708
rect 11659 29668 11704 29696
rect 11698 29656 11704 29668
rect 11756 29656 11762 29708
rect 12069 29699 12127 29705
rect 12069 29665 12081 29699
rect 12115 29665 12127 29699
rect 13078 29696 13084 29708
rect 13039 29668 13084 29696
rect 12069 29659 12127 29665
rect 9398 29628 9404 29640
rect 9359 29600 9404 29628
rect 9398 29588 9404 29600
rect 9456 29588 9462 29640
rect 11606 29628 11612 29640
rect 11567 29600 11612 29628
rect 11606 29588 11612 29600
rect 11664 29588 11670 29640
rect 7147 29532 8800 29560
rect 7147 29529 7159 29532
rect 7101 29523 7159 29529
rect 10594 29520 10600 29572
rect 10652 29560 10658 29572
rect 10870 29560 10876 29572
rect 10652 29532 10876 29560
rect 10652 29520 10658 29532
rect 10870 29520 10876 29532
rect 10928 29520 10934 29572
rect 11422 29520 11428 29572
rect 11480 29560 11486 29572
rect 12084 29560 12112 29659
rect 13078 29656 13084 29668
rect 13136 29656 13142 29708
rect 13253 29696 13259 29708
rect 13214 29668 13259 29696
rect 13253 29656 13259 29668
rect 13311 29656 13317 29708
rect 13446 29696 13452 29708
rect 13407 29668 13452 29696
rect 13446 29656 13452 29668
rect 13504 29656 13510 29708
rect 13633 29699 13691 29705
rect 13633 29665 13645 29699
rect 13679 29696 13691 29699
rect 14458 29696 14464 29708
rect 13679 29668 14464 29696
rect 13679 29665 13691 29668
rect 13633 29659 13691 29665
rect 14458 29656 14464 29668
rect 14516 29656 14522 29708
rect 14844 29705 14872 29736
rect 16025 29733 16037 29767
rect 16071 29764 16083 29767
rect 16574 29764 16580 29776
rect 16071 29736 16580 29764
rect 16071 29733 16083 29736
rect 16025 29727 16083 29733
rect 16574 29724 16580 29736
rect 16632 29764 16638 29776
rect 17494 29764 17500 29776
rect 16632 29736 17500 29764
rect 16632 29724 16638 29736
rect 17494 29724 17500 29736
rect 17552 29724 17558 29776
rect 17604 29764 17632 29804
rect 18049 29801 18061 29835
rect 18095 29832 18107 29835
rect 18138 29832 18144 29844
rect 18095 29804 18144 29832
rect 18095 29801 18107 29804
rect 18049 29795 18107 29801
rect 18138 29792 18144 29804
rect 18196 29792 18202 29844
rect 18874 29792 18880 29844
rect 18932 29792 18938 29844
rect 21174 29792 21180 29844
rect 21232 29832 21238 29844
rect 21232 29804 23796 29832
rect 21232 29792 21238 29804
rect 18892 29764 18920 29792
rect 22738 29764 22744 29776
rect 17604 29736 18920 29764
rect 22020 29736 22744 29764
rect 14829 29699 14887 29705
rect 14829 29665 14841 29699
rect 14875 29696 14887 29699
rect 15838 29696 15844 29708
rect 14875 29668 15844 29696
rect 14875 29665 14887 29668
rect 14829 29659 14887 29665
rect 15838 29656 15844 29668
rect 15896 29656 15902 29708
rect 16666 29696 16672 29708
rect 16627 29668 16672 29696
rect 16666 29656 16672 29668
rect 16724 29656 16730 29708
rect 16942 29705 16948 29708
rect 16936 29659 16948 29705
rect 17000 29696 17006 29708
rect 18877 29699 18935 29705
rect 17000 29668 17036 29696
rect 16942 29656 16948 29659
rect 17000 29656 17006 29668
rect 18877 29665 18889 29699
rect 18923 29696 18935 29699
rect 19334 29696 19340 29708
rect 18923 29668 19340 29696
rect 18923 29665 18935 29668
rect 18877 29659 18935 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 21266 29656 21272 29708
rect 21324 29696 21330 29708
rect 22020 29707 22048 29736
rect 22738 29724 22744 29736
rect 22796 29724 22802 29776
rect 23768 29773 23796 29804
rect 25590 29792 25596 29844
rect 25648 29832 25654 29844
rect 28166 29832 28172 29844
rect 25648 29804 28172 29832
rect 25648 29792 25654 29804
rect 28166 29792 28172 29804
rect 28224 29792 28230 29844
rect 29178 29792 29184 29844
rect 29236 29832 29242 29844
rect 29236 29804 31156 29832
rect 29236 29792 29242 29804
rect 23753 29767 23811 29773
rect 23753 29733 23765 29767
rect 23799 29764 23811 29767
rect 27154 29764 27160 29776
rect 23799 29736 27160 29764
rect 23799 29733 23811 29736
rect 23753 29727 23811 29733
rect 27154 29724 27160 29736
rect 27212 29724 27218 29776
rect 27798 29724 27804 29776
rect 27856 29764 27862 29776
rect 28546 29767 28604 29773
rect 28546 29764 28558 29767
rect 27856 29736 28558 29764
rect 27856 29724 27862 29736
rect 28546 29733 28558 29736
rect 28592 29733 28604 29767
rect 28546 29727 28604 29733
rect 28828 29736 30696 29764
rect 21821 29699 21879 29705
rect 21821 29696 21833 29699
rect 21324 29668 21833 29696
rect 21324 29656 21330 29668
rect 21821 29665 21833 29668
rect 21867 29665 21879 29699
rect 21821 29659 21879 29665
rect 22005 29701 22063 29707
rect 22005 29667 22017 29701
rect 22051 29667 22063 29701
rect 22186 29696 22192 29708
rect 22147 29668 22192 29696
rect 22005 29661 22063 29667
rect 22186 29656 22192 29668
rect 22244 29656 22250 29708
rect 22373 29699 22431 29705
rect 22373 29665 22385 29699
rect 22419 29696 22431 29699
rect 22462 29696 22468 29708
rect 22419 29668 22468 29696
rect 22419 29665 22431 29668
rect 22373 29659 22431 29665
rect 22462 29656 22468 29668
rect 22520 29656 22526 29708
rect 24854 29656 24860 29708
rect 24912 29696 24918 29708
rect 25501 29699 25559 29705
rect 25501 29696 25513 29699
rect 24912 29668 25513 29696
rect 24912 29656 24918 29668
rect 25501 29665 25513 29668
rect 25547 29696 25559 29699
rect 26050 29696 26056 29708
rect 25547 29668 26056 29696
rect 25547 29665 25559 29668
rect 25501 29659 25559 29665
rect 26050 29656 26056 29668
rect 26108 29656 26114 29708
rect 26145 29699 26203 29705
rect 26145 29665 26157 29699
rect 26191 29696 26203 29699
rect 26234 29696 26240 29708
rect 26191 29668 26240 29696
rect 26191 29665 26203 29668
rect 26145 29659 26203 29665
rect 26234 29656 26240 29668
rect 26292 29696 26298 29708
rect 26602 29696 26608 29708
rect 26292 29668 26608 29696
rect 26292 29656 26298 29668
rect 26602 29656 26608 29668
rect 26660 29656 26666 29708
rect 27982 29696 27988 29708
rect 27816 29668 27988 29696
rect 13354 29637 13360 29640
rect 13351 29591 13360 29637
rect 13412 29628 13418 29640
rect 13412 29600 13451 29628
rect 13354 29588 13360 29591
rect 13412 29588 13418 29600
rect 13814 29588 13820 29640
rect 13872 29628 13878 29640
rect 14553 29631 14611 29637
rect 14553 29628 14565 29631
rect 13872 29600 14565 29628
rect 13872 29588 13878 29600
rect 14553 29597 14565 29600
rect 14599 29628 14611 29631
rect 15194 29628 15200 29640
rect 14599 29600 15200 29628
rect 14599 29597 14611 29600
rect 14553 29591 14611 29597
rect 15194 29588 15200 29600
rect 15252 29588 15258 29640
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19153 29631 19211 29637
rect 19153 29628 19165 29631
rect 19024 29600 19165 29628
rect 19024 29588 19030 29600
rect 19153 29597 19165 29600
rect 19199 29597 19211 29631
rect 20162 29628 20168 29640
rect 20123 29600 20168 29628
rect 19153 29591 19211 29597
rect 20162 29588 20168 29600
rect 20220 29588 20226 29640
rect 20438 29628 20444 29640
rect 20399 29600 20444 29628
rect 20438 29588 20444 29600
rect 20496 29628 20502 29640
rect 22094 29628 22100 29640
rect 20496 29600 22100 29628
rect 20496 29588 20502 29600
rect 22094 29588 22100 29600
rect 22152 29588 22158 29640
rect 22278 29588 22284 29640
rect 22336 29628 22342 29640
rect 27816 29628 27844 29668
rect 27982 29656 27988 29668
rect 28040 29656 28046 29708
rect 28828 29705 28856 29736
rect 30668 29708 30696 29736
rect 28813 29699 28871 29705
rect 28813 29665 28825 29699
rect 28859 29665 28871 29699
rect 30374 29696 30380 29708
rect 30432 29705 30438 29708
rect 30344 29668 30380 29696
rect 28813 29659 28871 29665
rect 30374 29656 30380 29668
rect 30432 29659 30444 29705
rect 30650 29696 30656 29708
rect 30611 29668 30656 29696
rect 30432 29656 30438 29659
rect 30650 29656 30656 29668
rect 30708 29656 30714 29708
rect 31128 29705 31156 29804
rect 31113 29699 31171 29705
rect 31113 29665 31125 29699
rect 31159 29665 31171 29699
rect 31113 29659 31171 29665
rect 32320 29628 33120 29642
rect 22336 29600 27844 29628
rect 31772 29600 33120 29628
rect 22336 29588 22342 29600
rect 11480 29532 12112 29560
rect 11480 29520 11486 29532
rect 12342 29520 12348 29572
rect 12400 29560 12406 29572
rect 13446 29560 13452 29572
rect 12400 29532 13452 29560
rect 12400 29520 12406 29532
rect 13446 29520 13452 29532
rect 13504 29520 13510 29572
rect 20714 29560 20720 29572
rect 17788 29532 20720 29560
rect 3050 29492 3056 29504
rect 1903 29464 2774 29492
rect 3011 29464 3056 29492
rect 1903 29461 1915 29464
rect 1857 29455 1915 29461
rect 3050 29452 3056 29464
rect 3108 29452 3114 29504
rect 3142 29452 3148 29504
rect 3200 29492 3206 29504
rect 3200 29464 3245 29492
rect 3200 29452 3206 29464
rect 3602 29452 3608 29504
rect 3660 29492 3666 29504
rect 4985 29495 5043 29501
rect 4985 29492 4997 29495
rect 3660 29464 4997 29492
rect 3660 29452 3666 29464
rect 4985 29461 4997 29464
rect 5031 29492 5043 29495
rect 5350 29492 5356 29504
rect 5031 29464 5356 29492
rect 5031 29461 5043 29464
rect 4985 29455 5043 29461
rect 5350 29452 5356 29464
rect 5408 29452 5414 29504
rect 5718 29452 5724 29504
rect 5776 29492 5782 29504
rect 5813 29495 5871 29501
rect 5813 29492 5825 29495
rect 5776 29464 5825 29492
rect 5776 29452 5782 29464
rect 5813 29461 5825 29464
rect 5859 29461 5871 29495
rect 5813 29455 5871 29461
rect 7006 29452 7012 29504
rect 7064 29492 7070 29504
rect 8018 29492 8024 29504
rect 7064 29464 8024 29492
rect 7064 29452 7070 29464
rect 8018 29452 8024 29464
rect 8076 29452 8082 29504
rect 8846 29492 8852 29504
rect 8807 29464 8852 29492
rect 8846 29452 8852 29464
rect 8904 29452 8910 29504
rect 12066 29452 12072 29504
rect 12124 29492 12130 29504
rect 13078 29492 13084 29504
rect 12124 29464 13084 29492
rect 12124 29452 12130 29464
rect 13078 29452 13084 29464
rect 13136 29452 13142 29504
rect 13262 29452 13268 29504
rect 13320 29492 13326 29504
rect 13817 29495 13875 29501
rect 13817 29492 13829 29495
rect 13320 29464 13829 29492
rect 13320 29452 13326 29464
rect 13817 29461 13829 29464
rect 13863 29461 13875 29495
rect 13817 29455 13875 29461
rect 15194 29452 15200 29504
rect 15252 29492 15258 29504
rect 17788 29492 17816 29532
rect 20714 29520 20720 29532
rect 20772 29520 20778 29572
rect 23017 29563 23075 29569
rect 23017 29560 23029 29563
rect 22066 29532 23029 29560
rect 15252 29464 17816 29492
rect 15252 29452 15258 29464
rect 17862 29452 17868 29504
rect 17920 29492 17926 29504
rect 21082 29492 21088 29504
rect 17920 29464 21088 29492
rect 17920 29452 17926 29464
rect 21082 29452 21088 29464
rect 21140 29452 21146 29504
rect 21174 29452 21180 29504
rect 21232 29492 21238 29504
rect 22066 29492 22094 29532
rect 23017 29529 23029 29532
rect 23063 29560 23075 29563
rect 23106 29560 23112 29572
rect 23063 29532 23112 29560
rect 23063 29529 23075 29532
rect 23017 29523 23075 29529
rect 23106 29520 23112 29532
rect 23164 29520 23170 29572
rect 22554 29492 22560 29504
rect 21232 29464 22094 29492
rect 22515 29464 22560 29492
rect 21232 29452 21238 29464
rect 22554 29452 22560 29464
rect 22612 29452 22618 29504
rect 26050 29492 26056 29504
rect 26011 29464 26056 29492
rect 26050 29452 26056 29464
rect 26108 29452 26114 29504
rect 27433 29495 27491 29501
rect 27433 29461 27445 29495
rect 27479 29492 27491 29495
rect 27614 29492 27620 29504
rect 27479 29464 27620 29492
rect 27479 29461 27491 29464
rect 27433 29455 27491 29461
rect 27614 29452 27620 29464
rect 27672 29452 27678 29504
rect 28810 29452 28816 29504
rect 28868 29492 28874 29504
rect 29273 29495 29331 29501
rect 29273 29492 29285 29495
rect 28868 29464 29285 29492
rect 28868 29452 28874 29464
rect 29273 29461 29285 29464
rect 29319 29461 29331 29495
rect 29273 29455 29331 29461
rect 31297 29495 31355 29501
rect 31297 29461 31309 29495
rect 31343 29492 31355 29495
rect 31772 29492 31800 29600
rect 32320 29586 33120 29600
rect 31343 29464 31800 29492
rect 31343 29461 31355 29464
rect 31297 29455 31355 29461
rect 1104 29402 32016 29424
rect 1104 29350 6102 29402
rect 6154 29350 6166 29402
rect 6218 29350 6230 29402
rect 6282 29350 6294 29402
rect 6346 29350 6358 29402
rect 6410 29350 16405 29402
rect 16457 29350 16469 29402
rect 16521 29350 16533 29402
rect 16585 29350 16597 29402
rect 16649 29350 16661 29402
rect 16713 29350 26709 29402
rect 26761 29350 26773 29402
rect 26825 29350 26837 29402
rect 26889 29350 26901 29402
rect 26953 29350 26965 29402
rect 27017 29350 32016 29402
rect 1104 29328 32016 29350
rect 1394 29248 1400 29300
rect 1452 29288 1458 29300
rect 1762 29288 1768 29300
rect 1452 29260 1768 29288
rect 1452 29248 1458 29260
rect 1762 29248 1768 29260
rect 1820 29288 1826 29300
rect 3786 29288 3792 29300
rect 1820 29260 3792 29288
rect 1820 29248 1826 29260
rect 3786 29248 3792 29260
rect 3844 29248 3850 29300
rect 3881 29291 3939 29297
rect 3881 29257 3893 29291
rect 3927 29288 3939 29291
rect 4246 29288 4252 29300
rect 3927 29260 4252 29288
rect 3927 29257 3939 29260
rect 3881 29251 3939 29257
rect 4246 29248 4252 29260
rect 4304 29248 4310 29300
rect 4430 29248 4436 29300
rect 4488 29288 4494 29300
rect 4525 29291 4583 29297
rect 4525 29288 4537 29291
rect 4488 29260 4537 29288
rect 4488 29248 4494 29260
rect 4525 29257 4537 29260
rect 4571 29257 4583 29291
rect 4525 29251 4583 29257
rect 5644 29260 6516 29288
rect 1949 29223 2007 29229
rect 1949 29189 1961 29223
rect 1995 29220 2007 29223
rect 2958 29220 2964 29232
rect 1995 29192 2964 29220
rect 1995 29189 2007 29192
rect 1949 29183 2007 29189
rect 2958 29180 2964 29192
rect 3016 29180 3022 29232
rect 4982 29220 4988 29232
rect 3068 29192 4988 29220
rect 2498 29152 2504 29164
rect 2459 29124 2504 29152
rect 2498 29112 2504 29124
rect 2556 29112 2562 29164
rect 2682 29112 2688 29164
rect 2740 29152 2746 29164
rect 3068 29152 3096 29192
rect 4982 29180 4988 29192
rect 5040 29180 5046 29232
rect 2740 29124 3096 29152
rect 2740 29112 2746 29124
rect 3510 29112 3516 29164
rect 3568 29152 3574 29164
rect 3568 29124 4016 29152
rect 3568 29112 3574 29124
rect 3326 29044 3332 29096
rect 3384 29084 3390 29096
rect 3602 29084 3608 29096
rect 3384 29056 3608 29084
rect 3384 29044 3390 29056
rect 3602 29044 3608 29056
rect 3660 29084 3666 29096
rect 3789 29087 3847 29093
rect 3789 29084 3801 29087
rect 3660 29056 3801 29084
rect 3660 29044 3666 29056
rect 3789 29053 3801 29056
rect 3835 29053 3847 29087
rect 3988 29084 4016 29124
rect 4338 29112 4344 29164
rect 4396 29152 4402 29164
rect 4396 29124 5120 29152
rect 4396 29112 4402 29124
rect 4062 29084 4068 29096
rect 3975 29056 4068 29084
rect 3789 29047 3847 29053
rect 4062 29044 4068 29056
rect 4120 29084 4126 29096
rect 5092 29093 5120 29124
rect 4433 29087 4491 29093
rect 4433 29084 4445 29087
rect 4120 29056 4445 29084
rect 4120 29044 4126 29056
rect 4433 29053 4445 29056
rect 4479 29053 4491 29087
rect 4433 29047 4491 29053
rect 5077 29087 5135 29093
rect 5077 29053 5089 29087
rect 5123 29053 5135 29087
rect 5258 29084 5264 29096
rect 5219 29056 5264 29084
rect 5077 29047 5135 29053
rect 5258 29044 5264 29056
rect 5316 29044 5322 29096
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 1797 29019 1855 29025
rect 1797 28985 1809 29019
rect 1843 29016 1855 29019
rect 2777 29019 2835 29025
rect 2777 29016 2789 29019
rect 1843 28988 2789 29016
rect 1843 28985 1855 28988
rect 1797 28979 1855 28985
rect 2777 28985 2789 28988
rect 2823 29016 2835 29019
rect 5169 29019 5227 29025
rect 5169 29016 5181 29019
rect 2823 28988 5181 29016
rect 2823 28985 2835 28988
rect 2777 28979 2835 28985
rect 5169 28985 5181 28988
rect 5215 28985 5227 29019
rect 5644 29016 5672 29260
rect 5718 29180 5724 29232
rect 5776 29180 5782 29232
rect 5810 29180 5816 29232
rect 5868 29220 5874 29232
rect 6086 29220 6092 29232
rect 5868 29192 6092 29220
rect 5868 29180 5874 29192
rect 6086 29180 6092 29192
rect 6144 29180 6150 29232
rect 6488 29220 6516 29260
rect 6638 29248 6644 29300
rect 6696 29288 6702 29300
rect 7009 29291 7067 29297
rect 7009 29288 7021 29291
rect 6696 29260 7021 29288
rect 6696 29248 6702 29260
rect 7009 29257 7021 29260
rect 7055 29257 7067 29291
rect 10318 29288 10324 29300
rect 7009 29251 7067 29257
rect 7396 29260 10324 29288
rect 7190 29220 7196 29232
rect 6488 29192 7196 29220
rect 7190 29180 7196 29192
rect 7248 29180 7254 29232
rect 5736 29152 5764 29180
rect 6549 29155 6607 29161
rect 5736 29124 6224 29152
rect 5902 29084 5908 29096
rect 5863 29056 5908 29084
rect 5902 29044 5908 29056
rect 5960 29044 5966 29096
rect 6196 29093 6224 29124
rect 6549 29121 6561 29155
rect 6595 29152 6607 29155
rect 7396 29152 7424 29260
rect 10318 29248 10324 29260
rect 10376 29248 10382 29300
rect 10502 29288 10508 29300
rect 10463 29260 10508 29288
rect 10502 29248 10508 29260
rect 10560 29248 10566 29300
rect 11422 29248 11428 29300
rect 11480 29288 11486 29300
rect 11698 29288 11704 29300
rect 11480 29260 11560 29288
rect 11659 29260 11704 29288
rect 11480 29248 11486 29260
rect 10520 29192 11284 29220
rect 8386 29152 8392 29164
rect 6595 29124 7424 29152
rect 8347 29124 8392 29152
rect 6595 29121 6607 29124
rect 6549 29115 6607 29121
rect 8386 29112 8392 29124
rect 8444 29112 8450 29164
rect 6089 29087 6147 29093
rect 6089 29084 6101 29087
rect 6012 29056 6101 29084
rect 6012 29028 6040 29056
rect 6089 29053 6101 29056
rect 6135 29053 6147 29087
rect 6089 29047 6147 29053
rect 6181 29087 6239 29093
rect 6181 29053 6193 29087
rect 6227 29053 6239 29087
rect 6181 29047 6239 29053
rect 6307 29087 6365 29093
rect 6307 29053 6319 29087
rect 6353 29084 6365 29087
rect 8846 29084 8852 29096
rect 6353 29056 8852 29084
rect 6353 29053 6365 29056
rect 6307 29047 6365 29053
rect 8846 29044 8852 29056
rect 8904 29044 8910 29096
rect 5810 29016 5816 29028
rect 5644 28988 5816 29016
rect 5169 28979 5227 28985
rect 5810 28976 5816 28988
rect 5868 28976 5874 29028
rect 5994 28976 6000 29028
rect 6052 28976 6058 29028
rect 6546 28976 6552 29028
rect 6604 29016 6610 29028
rect 6914 29016 6920 29028
rect 6604 28988 6920 29016
rect 6604 28976 6610 28988
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 7190 28976 7196 29028
rect 7248 29016 7254 29028
rect 8122 29019 8180 29025
rect 8122 29016 8134 29019
rect 7248 28988 8134 29016
rect 7248 28976 7254 28988
rect 8122 28985 8134 28988
rect 8168 28985 8180 29019
rect 8122 28979 8180 28985
rect 9674 28976 9680 29028
rect 9732 29016 9738 29028
rect 9861 29019 9919 29025
rect 9861 29016 9873 29019
rect 9732 28988 9873 29016
rect 9732 28976 9738 28988
rect 9861 28985 9873 28988
rect 9907 28985 9919 29019
rect 9861 28979 9919 28985
rect 2682 28948 2688 28960
rect 2643 28920 2688 28948
rect 2682 28908 2688 28920
rect 2740 28908 2746 28960
rect 3145 28951 3203 28957
rect 3145 28917 3157 28951
rect 3191 28948 3203 28951
rect 3786 28948 3792 28960
rect 3191 28920 3792 28948
rect 3191 28917 3203 28920
rect 3145 28911 3203 28917
rect 3786 28908 3792 28920
rect 3844 28908 3850 28960
rect 4154 28908 4160 28960
rect 4212 28948 4218 28960
rect 7834 28948 7840 28960
rect 4212 28920 7840 28948
rect 4212 28908 4218 28920
rect 7834 28908 7840 28920
rect 7892 28908 7898 28960
rect 9033 28951 9091 28957
rect 9033 28917 9045 28951
rect 9079 28948 9091 28951
rect 9490 28948 9496 28960
rect 9079 28920 9496 28948
rect 9079 28917 9091 28920
rect 9033 28911 9091 28917
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 10520 28948 10548 29192
rect 10594 29112 10600 29164
rect 10652 29152 10658 29164
rect 10965 29155 11023 29161
rect 10965 29152 10977 29155
rect 10652 29124 10977 29152
rect 10652 29112 10658 29124
rect 10965 29121 10977 29124
rect 11011 29121 11023 29155
rect 10965 29115 11023 29121
rect 10689 29087 10747 29093
rect 10689 29053 10701 29087
rect 10735 29053 10747 29087
rect 10870 29084 10876 29096
rect 10831 29056 10876 29084
rect 10689 29047 10747 29053
rect 10704 29016 10732 29047
rect 10870 29044 10876 29056
rect 10928 29044 10934 29096
rect 11054 29084 11060 29096
rect 11015 29056 11060 29084
rect 11054 29044 11060 29056
rect 11112 29044 11118 29096
rect 11256 29093 11284 29192
rect 11532 29152 11560 29260
rect 11698 29248 11704 29260
rect 11756 29248 11762 29300
rect 12526 29288 12532 29300
rect 12487 29260 12532 29288
rect 12526 29248 12532 29260
rect 12584 29248 12590 29300
rect 16298 29248 16304 29300
rect 16356 29288 16362 29300
rect 19334 29288 19340 29300
rect 16356 29260 19196 29288
rect 19295 29260 19340 29288
rect 16356 29248 16362 29260
rect 11793 29223 11851 29229
rect 11793 29189 11805 29223
rect 11839 29220 11851 29223
rect 11882 29220 11888 29232
rect 11839 29192 11888 29220
rect 11839 29189 11851 29192
rect 11793 29183 11851 29189
rect 11882 29180 11888 29192
rect 11940 29220 11946 29232
rect 12066 29220 12072 29232
rect 11940 29192 12072 29220
rect 11940 29180 11946 29192
rect 12066 29180 12072 29192
rect 12124 29180 12130 29232
rect 18414 29220 18420 29232
rect 12268 29192 17264 29220
rect 18375 29192 18420 29220
rect 12268 29152 12296 29192
rect 11532 29124 12296 29152
rect 12342 29112 12348 29164
rect 12400 29152 12406 29164
rect 12897 29155 12955 29161
rect 12897 29152 12909 29155
rect 12400 29124 12909 29152
rect 12400 29112 12406 29124
rect 12897 29121 12909 29124
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 12989 29155 13047 29161
rect 12989 29121 13001 29155
rect 13035 29152 13047 29155
rect 13354 29152 13360 29164
rect 13035 29124 13360 29152
rect 13035 29121 13047 29124
rect 12989 29115 13047 29121
rect 13354 29112 13360 29124
rect 13412 29152 13418 29164
rect 14553 29155 14611 29161
rect 14553 29152 14565 29155
rect 13412 29124 14565 29152
rect 13412 29112 13418 29124
rect 14553 29121 14565 29124
rect 14599 29121 14611 29155
rect 14553 29115 14611 29121
rect 14645 29155 14703 29161
rect 14645 29121 14657 29155
rect 14691 29152 14703 29155
rect 15102 29152 15108 29164
rect 14691 29124 15108 29152
rect 14691 29121 14703 29124
rect 14645 29115 14703 29121
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 16114 29112 16120 29164
rect 16172 29152 16178 29164
rect 16850 29152 16856 29164
rect 16172 29124 16856 29152
rect 16172 29112 16178 29124
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 17236 29152 17264 29192
rect 18414 29180 18420 29192
rect 18472 29180 18478 29232
rect 19168 29220 19196 29260
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 19794 29288 19800 29300
rect 19755 29260 19800 29288
rect 19794 29248 19800 29260
rect 19852 29248 19858 29300
rect 21174 29288 21180 29300
rect 20272 29260 21180 29288
rect 20272 29220 20300 29260
rect 21174 29248 21180 29260
rect 21232 29248 21238 29300
rect 22094 29248 22100 29300
rect 22152 29288 22158 29300
rect 23290 29288 23296 29300
rect 22152 29260 23296 29288
rect 22152 29248 22158 29260
rect 23290 29248 23296 29260
rect 23348 29248 23354 29300
rect 26234 29248 26240 29300
rect 26292 29288 26298 29300
rect 27617 29291 27675 29297
rect 27617 29288 27629 29291
rect 26292 29260 27629 29288
rect 26292 29248 26298 29260
rect 27617 29257 27629 29260
rect 27663 29257 27675 29291
rect 27617 29251 27675 29257
rect 30650 29248 30656 29300
rect 30708 29288 30714 29300
rect 30708 29260 30972 29288
rect 30708 29248 30714 29260
rect 19168 29192 20300 29220
rect 17678 29152 17684 29164
rect 17236 29124 17356 29152
rect 17639 29124 17684 29152
rect 11241 29087 11299 29093
rect 11241 29053 11253 29087
rect 11287 29053 11299 29087
rect 11241 29047 11299 29053
rect 11330 29044 11336 29096
rect 11388 29084 11394 29096
rect 11701 29087 11759 29093
rect 11701 29084 11713 29087
rect 11388 29056 11713 29084
rect 11388 29044 11394 29056
rect 11701 29053 11713 29056
rect 11747 29084 11759 29087
rect 12710 29084 12716 29096
rect 11747 29056 12572 29084
rect 12671 29056 12716 29084
rect 11747 29053 11759 29056
rect 11701 29047 11759 29053
rect 11146 29016 11152 29028
rect 10704 28988 11152 29016
rect 11146 28976 11152 28988
rect 11204 28976 11210 29028
rect 11977 29019 12035 29025
rect 11977 28985 11989 29019
rect 12023 28985 12035 29019
rect 12544 29016 12572 29056
rect 12710 29044 12716 29056
rect 12768 29044 12774 29096
rect 13081 29087 13139 29093
rect 13081 29053 13093 29087
rect 13127 29053 13139 29087
rect 13081 29047 13139 29053
rect 13096 29016 13124 29047
rect 13170 29044 13176 29096
rect 13228 29084 13234 29096
rect 13265 29087 13323 29093
rect 13265 29084 13277 29087
rect 13228 29056 13277 29084
rect 13228 29044 13234 29056
rect 13265 29053 13277 29056
rect 13311 29053 13323 29087
rect 14274 29084 14280 29096
rect 14235 29056 14280 29084
rect 13265 29047 13323 29053
rect 14274 29044 14280 29056
rect 14332 29044 14338 29096
rect 14458 29084 14464 29096
rect 14419 29056 14464 29084
rect 14458 29044 14464 29056
rect 14516 29044 14522 29096
rect 14826 29084 14832 29096
rect 14787 29056 14832 29084
rect 14826 29044 14832 29056
rect 14884 29044 14890 29096
rect 15010 29084 15016 29096
rect 14971 29056 15016 29084
rect 15010 29044 15016 29056
rect 15068 29044 15074 29096
rect 15562 29084 15568 29096
rect 15523 29056 15568 29084
rect 15562 29044 15568 29056
rect 15620 29044 15626 29096
rect 16666 29044 16672 29096
rect 16724 29084 16730 29096
rect 17034 29084 17040 29096
rect 16724 29056 17040 29084
rect 16724 29044 16730 29056
rect 17034 29044 17040 29056
rect 17092 29044 17098 29096
rect 14090 29016 14096 29028
rect 12544 28988 13032 29016
rect 13096 28988 14096 29016
rect 11977 28979 12035 28985
rect 10962 28948 10968 28960
rect 10520 28920 10968 28948
rect 10962 28908 10968 28920
rect 11020 28908 11026 28960
rect 11054 28908 11060 28960
rect 11112 28948 11118 28960
rect 11992 28948 12020 28979
rect 12250 28948 12256 28960
rect 11112 28920 12256 28948
rect 11112 28908 11118 28920
rect 12250 28908 12256 28920
rect 12308 28908 12314 28960
rect 13004 28948 13032 28988
rect 14090 28976 14096 28988
rect 14148 29016 14154 29028
rect 14844 29016 14872 29044
rect 15838 29016 15844 29028
rect 14148 28988 14872 29016
rect 14936 28988 15844 29016
rect 14148 28976 14154 28988
rect 14936 28948 14964 28988
rect 15838 28976 15844 28988
rect 15896 28976 15902 29028
rect 16298 28948 16304 28960
rect 13004 28920 14964 28948
rect 16259 28920 16304 28948
rect 16298 28908 16304 28920
rect 16356 28908 16362 28960
rect 17328 28948 17356 29124
rect 17678 29112 17684 29124
rect 17736 29112 17742 29164
rect 17957 29155 18015 29161
rect 17957 29121 17969 29155
rect 18003 29152 18015 29155
rect 18966 29152 18972 29164
rect 18003 29124 18972 29152
rect 18003 29121 18015 29124
rect 17957 29115 18015 29121
rect 18966 29112 18972 29124
rect 19024 29112 19030 29164
rect 26142 29112 26148 29164
rect 26200 29152 26206 29164
rect 26237 29155 26295 29161
rect 26237 29152 26249 29155
rect 26200 29124 26249 29152
rect 26200 29112 26206 29124
rect 26237 29121 26249 29124
rect 26283 29121 26295 29155
rect 28166 29152 28172 29164
rect 28127 29124 28172 29152
rect 26237 29115 26295 29121
rect 28166 29112 28172 29124
rect 28224 29112 28230 29164
rect 28994 29152 29000 29164
rect 28276 29124 29000 29152
rect 18601 29087 18659 29093
rect 18601 29053 18613 29087
rect 18647 29084 18659 29087
rect 20162 29084 20168 29096
rect 18647 29056 20168 29084
rect 18647 29053 18659 29056
rect 18601 29047 18659 29053
rect 17494 28976 17500 29028
rect 17552 29016 17558 29028
rect 18616 29016 18644 29047
rect 20162 29044 20168 29056
rect 20220 29044 20226 29096
rect 21177 29087 21235 29093
rect 21177 29053 21189 29087
rect 21223 29084 21235 29087
rect 22002 29084 22008 29096
rect 21223 29056 22008 29084
rect 21223 29053 21235 29056
rect 21177 29047 21235 29053
rect 22002 29044 22008 29056
rect 22060 29084 22066 29096
rect 22186 29084 22192 29096
rect 22060 29056 22192 29084
rect 22060 29044 22066 29056
rect 22186 29044 22192 29056
rect 22244 29044 22250 29096
rect 23198 29044 23204 29096
rect 23256 29093 23262 29096
rect 23256 29084 23268 29093
rect 23256 29056 23301 29084
rect 23256 29047 23268 29056
rect 23256 29044 23262 29047
rect 23382 29044 23388 29096
rect 23440 29084 23446 29096
rect 23477 29087 23535 29093
rect 23477 29084 23489 29087
rect 23440 29056 23489 29084
rect 23440 29044 23446 29056
rect 23477 29053 23489 29056
rect 23523 29084 23535 29087
rect 24397 29087 24455 29093
rect 24397 29084 24409 29087
rect 23523 29056 24409 29084
rect 23523 29053 23535 29056
rect 23477 29047 23535 29053
rect 24397 29053 24409 29056
rect 24443 29084 24455 29087
rect 28276 29084 28304 29124
rect 28994 29112 29000 29124
rect 29052 29112 29058 29164
rect 30944 29161 30972 29260
rect 30929 29155 30987 29161
rect 30929 29121 30941 29155
rect 30975 29152 30987 29155
rect 31202 29152 31208 29164
rect 30975 29124 31208 29152
rect 30975 29121 30987 29124
rect 30929 29115 30987 29121
rect 31202 29112 31208 29124
rect 31260 29112 31266 29164
rect 24443 29056 24900 29084
rect 24443 29053 24455 29056
rect 24397 29047 24455 29053
rect 24872 29028 24900 29056
rect 26344 29056 28304 29084
rect 28445 29087 28503 29093
rect 17552 28988 18644 29016
rect 17552 28976 17558 28988
rect 19978 28976 19984 29028
rect 20036 29016 20042 29028
rect 20910 29019 20968 29025
rect 20910 29016 20922 29019
rect 20036 28988 20922 29016
rect 20036 28976 20042 28988
rect 20910 28985 20922 28988
rect 20956 28985 20968 29019
rect 20910 28979 20968 28985
rect 24578 28976 24584 29028
rect 24636 29025 24642 29028
rect 24636 29019 24700 29025
rect 24636 28985 24654 29019
rect 24688 28985 24700 29019
rect 24636 28979 24700 28985
rect 24636 28976 24642 28979
rect 24854 28976 24860 29028
rect 24912 28976 24918 29028
rect 25314 28976 25320 29028
rect 25372 29016 25378 29028
rect 26344 29016 26372 29056
rect 28445 29053 28457 29087
rect 28491 29084 28503 29087
rect 28626 29084 28632 29096
rect 28491 29056 28632 29084
rect 28491 29053 28503 29056
rect 28445 29047 28503 29053
rect 28626 29044 28632 29056
rect 28684 29044 28690 29096
rect 26510 29025 26516 29028
rect 25372 28988 26372 29016
rect 25372 28976 25378 28988
rect 26504 28979 26516 29025
rect 26568 29016 26574 29028
rect 26568 28988 26604 29016
rect 26510 28976 26516 28979
rect 26568 28976 26574 28988
rect 30282 28976 30288 29028
rect 30340 29016 30346 29028
rect 30662 29019 30720 29025
rect 30662 29016 30674 29019
rect 30340 28988 30674 29016
rect 30340 28976 30346 28988
rect 30662 28985 30674 28988
rect 30708 28985 30720 29019
rect 30662 28979 30720 28985
rect 18506 28948 18512 28960
rect 17328 28920 18512 28948
rect 18506 28908 18512 28920
rect 18564 28948 18570 28960
rect 19886 28948 19892 28960
rect 18564 28920 19892 28948
rect 18564 28908 18570 28920
rect 19886 28908 19892 28920
rect 19944 28908 19950 28960
rect 23198 28908 23204 28960
rect 23256 28948 23262 28960
rect 23382 28948 23388 28960
rect 23256 28920 23388 28948
rect 23256 28908 23262 28920
rect 23382 28908 23388 28920
rect 23440 28908 23446 28960
rect 25038 28908 25044 28960
rect 25096 28948 25102 28960
rect 25777 28951 25835 28957
rect 25777 28948 25789 28951
rect 25096 28920 25789 28948
rect 25096 28908 25102 28920
rect 25777 28917 25789 28920
rect 25823 28917 25835 28951
rect 25777 28911 25835 28917
rect 29086 28908 29092 28960
rect 29144 28948 29150 28960
rect 29549 28951 29607 28957
rect 29549 28948 29561 28951
rect 29144 28920 29561 28948
rect 29144 28908 29150 28920
rect 29549 28917 29561 28920
rect 29595 28917 29607 28951
rect 29549 28911 29607 28917
rect 1104 28858 32016 28880
rect 1104 28806 11253 28858
rect 11305 28806 11317 28858
rect 11369 28806 11381 28858
rect 11433 28806 11445 28858
rect 11497 28806 11509 28858
rect 11561 28806 21557 28858
rect 21609 28806 21621 28858
rect 21673 28806 21685 28858
rect 21737 28806 21749 28858
rect 21801 28806 21813 28858
rect 21865 28806 32016 28858
rect 1104 28784 32016 28806
rect 3878 28704 3884 28756
rect 3936 28744 3942 28756
rect 4062 28744 4068 28756
rect 3936 28716 4068 28744
rect 3936 28704 3942 28716
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 4338 28704 4344 28756
rect 4396 28744 4402 28756
rect 4433 28747 4491 28753
rect 4433 28744 4445 28747
rect 4396 28716 4445 28744
rect 4396 28704 4402 28716
rect 4433 28713 4445 28716
rect 4479 28713 4491 28747
rect 4433 28707 4491 28713
rect 5721 28747 5779 28753
rect 5721 28713 5733 28747
rect 5767 28744 5779 28747
rect 5902 28744 5908 28756
rect 5767 28716 5908 28744
rect 5767 28713 5779 28716
rect 5721 28707 5779 28713
rect 5902 28704 5908 28716
rect 5960 28704 5966 28756
rect 8846 28704 8852 28756
rect 8904 28744 8910 28756
rect 9214 28744 9220 28756
rect 8904 28716 9220 28744
rect 8904 28704 8910 28716
rect 9214 28704 9220 28716
rect 9272 28704 9278 28756
rect 11054 28744 11060 28756
rect 10428 28716 11060 28744
rect 1673 28679 1731 28685
rect 1673 28645 1685 28679
rect 1719 28676 1731 28679
rect 4154 28676 4160 28688
rect 1719 28648 2268 28676
rect 1719 28645 1731 28648
rect 1673 28639 1731 28645
rect 1946 28608 1952 28620
rect 1907 28580 1952 28608
rect 1946 28568 1952 28580
rect 2004 28568 2010 28620
rect 2240 28608 2268 28648
rect 3160 28648 4160 28676
rect 2685 28611 2743 28617
rect 2240 28606 2636 28608
rect 2685 28606 2697 28611
rect 2240 28580 2697 28606
rect 2608 28578 2697 28580
rect 2685 28577 2697 28578
rect 2731 28577 2743 28611
rect 3050 28608 3056 28620
rect 3011 28580 3056 28608
rect 2685 28571 2743 28577
rect 3050 28568 3056 28580
rect 3108 28568 3114 28620
rect 1670 28540 1676 28552
rect 1631 28512 1676 28540
rect 1670 28500 1676 28512
rect 1728 28500 1734 28552
rect 2314 28432 2320 28484
rect 2372 28472 2378 28484
rect 3160 28481 3188 28648
rect 4154 28636 4160 28648
rect 4212 28636 4218 28688
rect 4982 28636 4988 28688
rect 5040 28676 5046 28688
rect 5040 28648 6776 28676
rect 5040 28636 5046 28648
rect 3326 28608 3332 28620
rect 3287 28580 3332 28608
rect 3326 28568 3332 28580
rect 3384 28568 3390 28620
rect 4341 28611 4399 28617
rect 4341 28608 4353 28611
rect 3436 28580 4353 28608
rect 3145 28475 3203 28481
rect 2372 28444 3112 28472
rect 2372 28432 2378 28444
rect 1857 28407 1915 28413
rect 1857 28373 1869 28407
rect 1903 28404 1915 28407
rect 2406 28404 2412 28416
rect 1903 28376 2412 28404
rect 1903 28373 1915 28376
rect 1857 28367 1915 28373
rect 2406 28364 2412 28376
rect 2464 28364 2470 28416
rect 3084 28404 3112 28444
rect 3145 28441 3157 28475
rect 3191 28441 3203 28475
rect 3145 28435 3203 28441
rect 3436 28404 3464 28580
rect 4341 28577 4353 28580
rect 4387 28577 4399 28611
rect 4341 28571 4399 28577
rect 5445 28611 5503 28617
rect 5445 28577 5457 28611
rect 5491 28608 5503 28611
rect 6181 28611 6239 28617
rect 6181 28608 6193 28611
rect 5491 28580 6193 28608
rect 5491 28577 5503 28580
rect 5445 28571 5503 28577
rect 6181 28577 6193 28580
rect 6227 28577 6239 28611
rect 6181 28571 6239 28577
rect 6454 28568 6460 28620
rect 6512 28608 6518 28620
rect 6748 28617 6776 28648
rect 6641 28611 6699 28617
rect 6641 28608 6653 28611
rect 6512 28580 6653 28608
rect 6512 28568 6518 28580
rect 6641 28577 6653 28580
rect 6687 28577 6699 28611
rect 6641 28571 6699 28577
rect 6733 28611 6791 28617
rect 6733 28577 6745 28611
rect 6779 28577 6791 28611
rect 6733 28571 6791 28577
rect 6822 28568 6828 28620
rect 6880 28608 6886 28620
rect 7009 28611 7067 28617
rect 6880 28580 6925 28608
rect 6880 28568 6886 28580
rect 7009 28577 7021 28611
rect 7055 28577 7067 28611
rect 7009 28571 7067 28577
rect 7745 28611 7803 28617
rect 7745 28577 7757 28611
rect 7791 28608 7803 28611
rect 7926 28608 7932 28620
rect 7791 28580 7932 28608
rect 7791 28577 7803 28580
rect 7745 28571 7803 28577
rect 3697 28543 3755 28549
rect 3697 28509 3709 28543
rect 3743 28540 3755 28543
rect 3878 28540 3884 28552
rect 3743 28512 3884 28540
rect 3743 28509 3755 28512
rect 3697 28503 3755 28509
rect 3878 28500 3884 28512
rect 3936 28500 3942 28552
rect 4706 28500 4712 28552
rect 4764 28540 4770 28552
rect 5537 28543 5595 28549
rect 5537 28540 5549 28543
rect 4764 28512 5549 28540
rect 4764 28500 4770 28512
rect 5537 28509 5549 28512
rect 5583 28509 5595 28543
rect 5537 28503 5595 28509
rect 5721 28543 5779 28549
rect 5721 28509 5733 28543
rect 5767 28540 5779 28543
rect 6365 28543 6423 28549
rect 6365 28540 6377 28543
rect 5767 28512 6377 28540
rect 5767 28509 5779 28512
rect 5721 28503 5779 28509
rect 6365 28509 6377 28512
rect 6411 28509 6423 28543
rect 6365 28503 6423 28509
rect 6914 28500 6920 28552
rect 6972 28540 6978 28552
rect 7024 28540 7052 28571
rect 7926 28568 7932 28580
rect 7984 28568 7990 28620
rect 8570 28568 8576 28620
rect 8628 28608 8634 28620
rect 9217 28611 9275 28617
rect 9217 28608 9229 28611
rect 8628 28580 9229 28608
rect 8628 28568 8634 28580
rect 9217 28577 9229 28580
rect 9263 28577 9275 28611
rect 9217 28571 9275 28577
rect 9585 28611 9643 28617
rect 9585 28577 9597 28611
rect 9631 28608 9643 28611
rect 9674 28608 9680 28620
rect 9631 28580 9680 28608
rect 9631 28577 9643 28580
rect 9585 28571 9643 28577
rect 9674 28568 9680 28580
rect 9732 28568 9738 28620
rect 10428 28617 10456 28716
rect 11054 28704 11060 28716
rect 11112 28704 11118 28756
rect 11517 28747 11575 28753
rect 11517 28713 11529 28747
rect 11563 28744 11575 28747
rect 11882 28744 11888 28756
rect 11563 28716 11888 28744
rect 11563 28713 11575 28716
rect 11517 28707 11575 28713
rect 11882 28704 11888 28716
rect 11940 28704 11946 28756
rect 12986 28704 12992 28756
rect 13044 28744 13050 28756
rect 13170 28744 13176 28756
rect 13044 28716 13176 28744
rect 13044 28704 13050 28716
rect 13170 28704 13176 28716
rect 13228 28704 13234 28756
rect 14274 28704 14280 28756
rect 14332 28744 14338 28756
rect 14369 28747 14427 28753
rect 14369 28744 14381 28747
rect 14332 28716 14381 28744
rect 14332 28704 14338 28716
rect 14369 28713 14381 28716
rect 14415 28744 14427 28747
rect 14458 28744 14464 28756
rect 14415 28716 14464 28744
rect 14415 28713 14427 28716
rect 14369 28707 14427 28713
rect 14458 28704 14464 28716
rect 14516 28744 14522 28756
rect 16669 28747 16727 28753
rect 14516 28716 16068 28744
rect 14516 28704 14522 28716
rect 10594 28636 10600 28688
rect 10652 28636 10658 28688
rect 11146 28676 11152 28688
rect 10796 28648 11152 28676
rect 9769 28611 9827 28617
rect 9769 28577 9781 28611
rect 9815 28577 9827 28611
rect 9769 28571 9827 28577
rect 10413 28611 10471 28617
rect 10413 28577 10425 28611
rect 10459 28577 10471 28611
rect 10612 28608 10640 28636
rect 10796 28617 10824 28648
rect 11146 28636 11152 28648
rect 11204 28636 11210 28688
rect 13262 28685 13268 28688
rect 13256 28676 13268 28685
rect 13223 28648 13268 28676
rect 13256 28639 13268 28648
rect 13262 28636 13268 28639
rect 13320 28636 13326 28688
rect 15289 28679 15347 28685
rect 15289 28645 15301 28679
rect 15335 28676 15347 28679
rect 15930 28676 15936 28688
rect 15335 28648 15936 28676
rect 15335 28645 15347 28648
rect 15289 28639 15347 28645
rect 15930 28636 15936 28648
rect 15988 28636 15994 28688
rect 10689 28611 10747 28617
rect 10689 28608 10701 28611
rect 10612 28580 10701 28608
rect 10413 28571 10471 28577
rect 10689 28577 10701 28580
rect 10735 28577 10747 28611
rect 10689 28571 10747 28577
rect 10781 28611 10839 28617
rect 10781 28577 10793 28611
rect 10827 28577 10839 28611
rect 10962 28608 10968 28620
rect 10923 28580 10968 28608
rect 10781 28571 10839 28577
rect 6972 28512 7052 28540
rect 6972 28500 6978 28512
rect 7190 28500 7196 28552
rect 7248 28540 7254 28552
rect 8021 28543 8079 28549
rect 8021 28540 8033 28543
rect 7248 28512 8033 28540
rect 7248 28500 7254 28512
rect 8021 28509 8033 28512
rect 8067 28540 8079 28543
rect 9401 28543 9459 28549
rect 9401 28540 9413 28543
rect 8067 28512 9413 28540
rect 8067 28509 8079 28512
rect 8021 28503 8079 28509
rect 9401 28509 9413 28512
rect 9447 28509 9459 28543
rect 9401 28503 9459 28509
rect 9490 28500 9496 28552
rect 9548 28540 9554 28552
rect 9548 28512 9593 28540
rect 9548 28500 9554 28512
rect 6086 28472 6092 28484
rect 5847 28444 6092 28472
rect 3084 28376 3464 28404
rect 4154 28364 4160 28416
rect 4212 28404 4218 28416
rect 4798 28404 4804 28416
rect 4212 28376 4804 28404
rect 4212 28364 4218 28376
rect 4798 28364 4804 28376
rect 4856 28364 4862 28416
rect 5626 28364 5632 28416
rect 5684 28404 5690 28416
rect 5847 28404 5875 28444
rect 6086 28432 6092 28444
rect 6144 28432 6150 28484
rect 6181 28475 6239 28481
rect 6181 28441 6193 28475
rect 6227 28472 6239 28475
rect 7282 28472 7288 28484
rect 6227 28444 7288 28472
rect 6227 28441 6239 28444
rect 6181 28435 6239 28441
rect 7282 28432 7288 28444
rect 7340 28432 7346 28484
rect 7834 28432 7840 28484
rect 7892 28472 7898 28484
rect 9784 28472 9812 28571
rect 10962 28568 10968 28580
rect 11020 28568 11026 28620
rect 11164 28608 11192 28636
rect 11701 28611 11759 28617
rect 11701 28608 11713 28611
rect 11164 28580 11713 28608
rect 11701 28577 11713 28580
rect 11747 28577 11759 28611
rect 12066 28608 12072 28620
rect 12027 28580 12072 28608
rect 11701 28571 11759 28577
rect 12066 28568 12072 28580
rect 12124 28568 12130 28620
rect 12250 28608 12256 28620
rect 12211 28580 12256 28608
rect 12250 28568 12256 28580
rect 12308 28568 12314 28620
rect 15010 28608 15016 28620
rect 14971 28580 15016 28608
rect 15010 28568 15016 28580
rect 15068 28568 15074 28620
rect 15381 28611 15439 28617
rect 15381 28577 15393 28611
rect 15427 28577 15439 28611
rect 15381 28571 15439 28577
rect 15841 28611 15899 28617
rect 15841 28577 15853 28611
rect 15887 28608 15899 28611
rect 16040 28608 16068 28716
rect 16669 28713 16681 28747
rect 16715 28744 16727 28747
rect 16850 28744 16856 28756
rect 16715 28716 16856 28744
rect 16715 28713 16727 28716
rect 16669 28707 16727 28713
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 18138 28744 18144 28756
rect 16960 28716 18144 28744
rect 16960 28676 16988 28716
rect 18138 28704 18144 28716
rect 18196 28704 18202 28756
rect 19978 28744 19984 28756
rect 19939 28716 19984 28744
rect 19978 28704 19984 28716
rect 20036 28704 20042 28756
rect 21269 28747 21327 28753
rect 21269 28713 21281 28747
rect 21315 28744 21327 28747
rect 23937 28747 23995 28753
rect 21315 28716 23888 28744
rect 21315 28713 21327 28716
rect 21269 28707 21327 28713
rect 17678 28676 17684 28688
rect 16868 28648 16988 28676
rect 17052 28648 17684 28676
rect 16868 28617 16896 28648
rect 17052 28617 17080 28648
rect 17678 28636 17684 28648
rect 17736 28636 17742 28688
rect 18230 28676 18236 28688
rect 17880 28648 18236 28676
rect 15887 28580 16068 28608
rect 16853 28611 16911 28617
rect 15887 28577 15899 28580
rect 15841 28571 15899 28577
rect 16853 28577 16865 28611
rect 16899 28577 16911 28611
rect 16853 28571 16911 28577
rect 17037 28611 17095 28617
rect 17037 28577 17049 28611
rect 17083 28577 17095 28611
rect 17037 28571 17095 28577
rect 17221 28611 17279 28617
rect 17221 28577 17233 28611
rect 17267 28577 17279 28611
rect 17221 28571 17279 28577
rect 10597 28543 10655 28549
rect 10597 28509 10609 28543
rect 10643 28509 10655 28543
rect 10597 28503 10655 28509
rect 7892 28444 9812 28472
rect 7892 28432 7898 28444
rect 9858 28432 9864 28484
rect 9916 28472 9922 28484
rect 10612 28472 10640 28503
rect 11790 28500 11796 28552
rect 11848 28540 11854 28552
rect 11885 28543 11943 28549
rect 11885 28540 11897 28543
rect 11848 28512 11897 28540
rect 11848 28500 11854 28512
rect 11885 28509 11897 28512
rect 11931 28509 11943 28543
rect 11885 28503 11943 28509
rect 11977 28543 12035 28549
rect 11977 28509 11989 28543
rect 12023 28509 12035 28543
rect 11977 28503 12035 28509
rect 10870 28472 10876 28484
rect 9916 28444 10548 28472
rect 10612 28444 10876 28472
rect 9916 28432 9922 28444
rect 5684 28376 5875 28404
rect 9033 28407 9091 28413
rect 5684 28364 5690 28376
rect 9033 28373 9045 28407
rect 9079 28404 9091 28407
rect 9214 28404 9220 28416
rect 9079 28376 9220 28404
rect 9079 28373 9091 28376
rect 9033 28367 9091 28373
rect 9214 28364 9220 28376
rect 9272 28364 9278 28416
rect 10226 28404 10232 28416
rect 10187 28376 10232 28404
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 10520 28404 10548 28444
rect 10870 28432 10876 28444
rect 10928 28472 10934 28484
rect 11992 28472 12020 28503
rect 12158 28500 12164 28552
rect 12216 28540 12222 28552
rect 12986 28540 12992 28552
rect 12216 28512 12992 28540
rect 12216 28500 12222 28512
rect 12986 28500 12992 28512
rect 13044 28500 13050 28552
rect 14826 28540 14832 28552
rect 14787 28512 14832 28540
rect 14826 28500 14832 28512
rect 14884 28500 14890 28552
rect 15396 28540 15424 28571
rect 15930 28540 15936 28552
rect 15396 28512 15936 28540
rect 15930 28500 15936 28512
rect 15988 28500 15994 28552
rect 17126 28540 17132 28552
rect 17087 28512 17132 28540
rect 17126 28500 17132 28512
rect 17184 28500 17190 28552
rect 17236 28540 17264 28571
rect 17310 28568 17316 28620
rect 17368 28608 17374 28620
rect 17405 28611 17463 28617
rect 17405 28608 17417 28611
rect 17368 28580 17417 28608
rect 17368 28568 17374 28580
rect 17405 28577 17417 28580
rect 17451 28608 17463 28611
rect 17880 28608 17908 28648
rect 18230 28636 18236 28648
rect 18288 28636 18294 28688
rect 20622 28676 20628 28688
rect 20535 28648 20628 28676
rect 17451 28580 17908 28608
rect 17451 28577 17463 28580
rect 17405 28571 17463 28577
rect 17954 28568 17960 28620
rect 18012 28608 18018 28620
rect 18121 28611 18179 28617
rect 18121 28608 18133 28611
rect 18012 28580 18133 28608
rect 18012 28568 18018 28580
rect 18121 28577 18133 28580
rect 18167 28577 18179 28611
rect 18121 28571 18179 28577
rect 19794 28568 19800 28620
rect 19852 28608 19858 28620
rect 20162 28608 20168 28620
rect 19852 28580 20168 28608
rect 19852 28568 19858 28580
rect 20162 28568 20168 28580
rect 20220 28568 20226 28620
rect 20438 28608 20444 28620
rect 20399 28580 20444 28608
rect 20438 28568 20444 28580
rect 20496 28568 20502 28620
rect 20548 28617 20576 28648
rect 20622 28636 20628 28648
rect 20680 28676 20686 28688
rect 22094 28676 22100 28688
rect 20680 28648 22100 28676
rect 20680 28636 20686 28648
rect 22094 28636 22100 28648
rect 22152 28636 22158 28688
rect 22186 28636 22192 28688
rect 22244 28676 22250 28688
rect 23198 28676 23204 28688
rect 22244 28648 23204 28676
rect 22244 28636 22250 28648
rect 23198 28636 23204 28648
rect 23256 28636 23262 28688
rect 23860 28676 23888 28716
rect 23937 28713 23949 28747
rect 23983 28744 23995 28747
rect 24302 28744 24308 28756
rect 23983 28716 24308 28744
rect 23983 28713 23995 28716
rect 23937 28707 23995 28713
rect 24302 28704 24308 28716
rect 24360 28704 24366 28756
rect 26142 28744 26148 28756
rect 24964 28716 26148 28744
rect 24964 28688 24992 28716
rect 26142 28704 26148 28716
rect 26200 28704 26206 28756
rect 26421 28747 26479 28753
rect 26421 28713 26433 28747
rect 26467 28744 26479 28747
rect 26510 28744 26516 28756
rect 26467 28716 26516 28744
rect 26467 28713 26479 28716
rect 26421 28707 26479 28713
rect 26510 28704 26516 28716
rect 26568 28704 26574 28756
rect 28169 28747 28227 28753
rect 28169 28713 28181 28747
rect 28215 28744 28227 28747
rect 30374 28744 30380 28756
rect 28215 28716 30380 28744
rect 28215 28713 28227 28716
rect 28169 28707 28227 28713
rect 30374 28704 30380 28716
rect 30432 28704 30438 28756
rect 24762 28676 24768 28688
rect 23860 28648 24768 28676
rect 24762 28636 24768 28648
rect 24820 28636 24826 28688
rect 24946 28676 24952 28688
rect 24872 28648 24952 28676
rect 20533 28611 20591 28617
rect 20533 28577 20545 28611
rect 20579 28577 20591 28611
rect 20533 28571 20591 28577
rect 20717 28611 20775 28617
rect 20717 28577 20729 28611
rect 20763 28608 20775 28611
rect 21266 28608 21272 28620
rect 20763 28580 21272 28608
rect 20763 28577 20775 28580
rect 20717 28571 20775 28577
rect 21266 28568 21272 28580
rect 21324 28568 21330 28620
rect 22554 28568 22560 28620
rect 22612 28608 22618 28620
rect 23118 28611 23176 28617
rect 23118 28608 23130 28611
rect 22612 28580 23130 28608
rect 22612 28568 22618 28580
rect 23118 28577 23130 28580
rect 23164 28577 23176 28611
rect 23216 28608 23244 28636
rect 23360 28611 23418 28617
rect 23360 28608 23372 28611
rect 23216 28580 23372 28608
rect 23118 28571 23176 28577
rect 23360 28577 23372 28580
rect 23406 28577 23418 28611
rect 23360 28571 23418 28577
rect 23750 28568 23756 28620
rect 23808 28608 23814 28620
rect 24872 28617 24900 28648
rect 24946 28636 24952 28648
rect 25004 28636 25010 28688
rect 25792 28648 27476 28676
rect 24029 28611 24087 28617
rect 24029 28608 24041 28611
rect 23808 28580 24041 28608
rect 23808 28568 23814 28580
rect 24029 28577 24041 28580
rect 24075 28577 24087 28611
rect 24029 28571 24087 28577
rect 24673 28611 24731 28617
rect 24673 28577 24685 28611
rect 24719 28577 24731 28611
rect 24673 28571 24731 28577
rect 24857 28611 24915 28617
rect 24857 28577 24869 28611
rect 24903 28577 24915 28611
rect 25038 28608 25044 28620
rect 24999 28580 25044 28608
rect 24857 28571 24915 28577
rect 17770 28540 17776 28552
rect 17236 28512 17776 28540
rect 12342 28472 12348 28484
rect 10928 28444 11928 28472
rect 11992 28444 12348 28472
rect 10928 28432 10934 28444
rect 11900 28416 11928 28444
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 16666 28432 16672 28484
rect 16724 28472 16730 28484
rect 17034 28472 17040 28484
rect 16724 28444 17040 28472
rect 16724 28432 16730 28444
rect 17034 28432 17040 28444
rect 17092 28432 17098 28484
rect 11790 28404 11796 28416
rect 10520 28376 11796 28404
rect 11790 28364 11796 28376
rect 11848 28364 11854 28416
rect 11882 28364 11888 28416
rect 11940 28364 11946 28416
rect 14642 28364 14648 28416
rect 14700 28404 14706 28416
rect 15933 28407 15991 28413
rect 15933 28404 15945 28407
rect 14700 28376 15945 28404
rect 14700 28364 14706 28376
rect 15933 28373 15945 28376
rect 15979 28373 15991 28407
rect 15933 28367 15991 28373
rect 16850 28364 16856 28416
rect 16908 28404 16914 28416
rect 17236 28404 17264 28512
rect 17770 28500 17776 28512
rect 17828 28500 17834 28552
rect 17865 28543 17923 28549
rect 17865 28509 17877 28543
rect 17911 28509 17923 28543
rect 20346 28540 20352 28552
rect 20307 28512 20352 28540
rect 17865 28503 17923 28509
rect 17880 28472 17908 28503
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 24688 28472 24716 28571
rect 25038 28568 25044 28580
rect 25096 28568 25102 28620
rect 25225 28611 25283 28617
rect 25225 28577 25237 28611
rect 25271 28608 25283 28611
rect 25682 28608 25688 28620
rect 25271 28580 25688 28608
rect 25271 28577 25283 28580
rect 25225 28571 25283 28577
rect 25682 28568 25688 28580
rect 25740 28608 25746 28620
rect 25792 28608 25820 28648
rect 25740 28580 25820 28608
rect 25740 28578 25748 28580
rect 25740 28568 25746 28578
rect 25866 28568 25872 28620
rect 25924 28608 25930 28620
rect 26234 28608 26240 28620
rect 25924 28580 25969 28608
rect 26195 28580 26240 28608
rect 25924 28568 25930 28580
rect 26234 28568 26240 28580
rect 26292 28568 26298 28620
rect 27448 28617 27476 28648
rect 27433 28611 27491 28617
rect 27433 28577 27445 28611
rect 27479 28577 27491 28611
rect 27614 28608 27620 28620
rect 27575 28580 27620 28608
rect 27433 28571 27491 28577
rect 27614 28568 27620 28580
rect 27672 28568 27678 28620
rect 27985 28611 28043 28617
rect 27985 28577 27997 28611
rect 28031 28577 28043 28611
rect 28626 28608 28632 28620
rect 28587 28580 28632 28608
rect 27985 28571 28043 28577
rect 24949 28543 25007 28549
rect 24949 28509 24961 28543
rect 24995 28540 25007 28543
rect 25961 28543 26019 28549
rect 25961 28540 25973 28543
rect 24995 28512 25973 28540
rect 24995 28509 25007 28512
rect 24949 28503 25007 28509
rect 25961 28509 25973 28512
rect 26007 28509 26019 28543
rect 25961 28503 26019 28509
rect 26053 28543 26111 28549
rect 26053 28509 26065 28543
rect 26099 28540 26111 28543
rect 26142 28540 26148 28552
rect 26099 28512 26148 28540
rect 26099 28509 26111 28512
rect 26053 28503 26111 28509
rect 25866 28472 25872 28484
rect 17788 28444 17908 28472
rect 23391 28444 24624 28472
rect 24688 28444 25872 28472
rect 17788 28416 17816 28444
rect 16908 28376 17264 28404
rect 16908 28364 16914 28376
rect 17770 28364 17776 28416
rect 17828 28364 17834 28416
rect 18046 28364 18052 28416
rect 18104 28404 18110 28416
rect 19150 28404 19156 28416
rect 18104 28376 19156 28404
rect 18104 28364 18110 28376
rect 19150 28364 19156 28376
rect 19208 28404 19214 28416
rect 19245 28407 19303 28413
rect 19245 28404 19257 28407
rect 19208 28376 19257 28404
rect 19208 28364 19214 28376
rect 19245 28373 19257 28376
rect 19291 28373 19303 28407
rect 19245 28367 19303 28373
rect 22005 28407 22063 28413
rect 22005 28373 22017 28407
rect 22051 28404 22063 28407
rect 22278 28404 22284 28416
rect 22051 28376 22284 28404
rect 22051 28373 22063 28376
rect 22005 28367 22063 28373
rect 22278 28364 22284 28376
rect 22336 28404 22342 28416
rect 22462 28404 22468 28416
rect 22336 28376 22468 28404
rect 22336 28364 22342 28376
rect 22462 28364 22468 28376
rect 22520 28364 22526 28416
rect 22738 28364 22744 28416
rect 22796 28404 22802 28416
rect 23391 28404 23419 28444
rect 24486 28404 24492 28416
rect 22796 28376 23419 28404
rect 24447 28376 24492 28404
rect 22796 28364 22802 28376
rect 24486 28364 24492 28376
rect 24544 28364 24550 28416
rect 24596 28404 24624 28444
rect 25866 28432 25872 28444
rect 25924 28432 25930 28484
rect 25976 28472 26004 28503
rect 26142 28500 26148 28512
rect 26200 28500 26206 28552
rect 27709 28543 27767 28549
rect 27709 28509 27721 28543
rect 27755 28509 27767 28543
rect 27709 28503 27767 28509
rect 27801 28543 27859 28549
rect 27801 28509 27813 28543
rect 27847 28509 27859 28543
rect 28000 28540 28028 28571
rect 28626 28568 28632 28580
rect 28684 28568 28690 28620
rect 28813 28611 28871 28617
rect 28813 28577 28825 28611
rect 28859 28608 28871 28611
rect 29086 28608 29092 28620
rect 28859 28580 29092 28608
rect 28859 28577 28871 28580
rect 28813 28571 28871 28577
rect 29086 28568 29092 28580
rect 29144 28568 29150 28620
rect 29181 28611 29239 28617
rect 29181 28577 29193 28611
rect 29227 28577 29239 28611
rect 29181 28571 29239 28577
rect 29365 28611 29423 28617
rect 29365 28577 29377 28611
rect 29411 28608 29423 28611
rect 30938 28611 30996 28617
rect 30938 28608 30950 28611
rect 29411 28580 30950 28608
rect 29411 28577 29423 28580
rect 29365 28571 29423 28577
rect 30938 28577 30950 28580
rect 30984 28577 30996 28611
rect 31202 28608 31208 28620
rect 31163 28580 31208 28608
rect 30938 28571 30996 28577
rect 28718 28540 28724 28552
rect 28000 28512 28724 28540
rect 27801 28503 27859 28509
rect 27522 28472 27528 28484
rect 25976 28444 27528 28472
rect 27522 28432 27528 28444
rect 27580 28472 27586 28484
rect 27724 28472 27752 28503
rect 27580 28444 27752 28472
rect 27816 28472 27844 28503
rect 28718 28500 28724 28512
rect 28776 28500 28782 28552
rect 28902 28540 28908 28552
rect 28863 28512 28908 28540
rect 28902 28500 28908 28512
rect 28960 28500 28966 28552
rect 28994 28500 29000 28552
rect 29052 28540 29058 28552
rect 29196 28540 29224 28571
rect 31202 28568 31208 28580
rect 31260 28568 31266 28620
rect 29052 28512 29097 28540
rect 29196 28512 29776 28540
rect 29052 28500 29058 28512
rect 29012 28472 29040 28500
rect 27816 28444 29040 28472
rect 27580 28432 27586 28444
rect 29748 28416 29776 28512
rect 24946 28404 24952 28416
rect 24596 28376 24952 28404
rect 24946 28364 24952 28376
rect 25004 28404 25010 28416
rect 28534 28404 28540 28416
rect 25004 28376 28540 28404
rect 25004 28364 25010 28376
rect 28534 28364 28540 28376
rect 28592 28364 28598 28416
rect 29730 28364 29736 28416
rect 29788 28404 29794 28416
rect 29825 28407 29883 28413
rect 29825 28404 29837 28407
rect 29788 28376 29837 28404
rect 29788 28364 29794 28376
rect 29825 28373 29837 28376
rect 29871 28373 29883 28407
rect 29825 28367 29883 28373
rect 1104 28314 32016 28336
rect 1104 28262 6102 28314
rect 6154 28262 6166 28314
rect 6218 28262 6230 28314
rect 6282 28262 6294 28314
rect 6346 28262 6358 28314
rect 6410 28262 16405 28314
rect 16457 28262 16469 28314
rect 16521 28262 16533 28314
rect 16585 28262 16597 28314
rect 16649 28262 16661 28314
rect 16713 28262 26709 28314
rect 26761 28262 26773 28314
rect 26825 28262 26837 28314
rect 26889 28262 26901 28314
rect 26953 28262 26965 28314
rect 27017 28262 32016 28314
rect 1104 28240 32016 28262
rect 1302 28160 1308 28212
rect 1360 28200 1366 28212
rect 1581 28203 1639 28209
rect 1581 28200 1593 28203
rect 1360 28172 1593 28200
rect 1360 28160 1366 28172
rect 1581 28169 1593 28172
rect 1627 28169 1639 28203
rect 1581 28163 1639 28169
rect 2406 28160 2412 28212
rect 2464 28200 2470 28212
rect 3878 28200 3884 28212
rect 2464 28172 3464 28200
rect 3839 28172 3884 28200
rect 2464 28160 2470 28172
rect 1210 28092 1216 28144
rect 1268 28132 1274 28144
rect 3053 28135 3111 28141
rect 1268 28104 3004 28132
rect 1268 28092 1274 28104
rect 2409 28067 2467 28073
rect 2409 28033 2421 28067
rect 2455 28064 2467 28067
rect 2682 28064 2688 28076
rect 2455 28036 2688 28064
rect 2455 28033 2467 28036
rect 2409 28027 2467 28033
rect 2682 28024 2688 28036
rect 2740 28024 2746 28076
rect 2976 28064 3004 28104
rect 3053 28101 3065 28135
rect 3099 28132 3111 28135
rect 3326 28132 3332 28144
rect 3099 28104 3332 28132
rect 3099 28101 3111 28104
rect 3053 28095 3111 28101
rect 3326 28092 3332 28104
rect 3384 28092 3390 28144
rect 3436 28132 3464 28172
rect 3878 28160 3884 28172
rect 3936 28160 3942 28212
rect 4890 28200 4896 28212
rect 4851 28172 4896 28200
rect 4890 28160 4896 28172
rect 4948 28160 4954 28212
rect 4982 28160 4988 28212
rect 5040 28200 5046 28212
rect 7098 28200 7104 28212
rect 5040 28172 6316 28200
rect 7059 28172 7104 28200
rect 5040 28160 5046 28172
rect 4154 28132 4160 28144
rect 3436 28104 4160 28132
rect 4154 28092 4160 28104
rect 4212 28092 4218 28144
rect 4430 28064 4436 28076
rect 2976 28036 4436 28064
rect 4430 28024 4436 28036
rect 4488 28064 4494 28076
rect 4798 28064 4804 28076
rect 4488 28036 4804 28064
rect 4488 28024 4494 28036
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 4908 28036 5580 28064
rect 4908 28008 4936 28036
rect 1486 27996 1492 28008
rect 1447 27968 1492 27996
rect 1486 27956 1492 27968
rect 1544 27956 1550 28008
rect 2593 27999 2651 28005
rect 2593 27965 2605 27999
rect 2639 27965 2651 27999
rect 2774 27996 2780 28008
rect 2735 27968 2780 27996
rect 2593 27959 2651 27965
rect 2608 27928 2636 27959
rect 2774 27956 2780 27968
rect 2832 27956 2838 28008
rect 2958 27956 2964 28008
rect 3016 27996 3022 28008
rect 3053 27999 3111 28005
rect 3053 27996 3065 27999
rect 3016 27968 3065 27996
rect 3016 27956 3022 27968
rect 3053 27965 3065 27968
rect 3099 27965 3111 27999
rect 3786 27996 3792 28008
rect 3747 27968 3792 27996
rect 3053 27959 3111 27965
rect 3786 27956 3792 27968
rect 3844 27956 3850 28008
rect 4890 27996 4896 28008
rect 4803 27968 4896 27996
rect 4890 27956 4896 27968
rect 4948 27956 4954 28008
rect 5552 28005 5580 28036
rect 5847 28005 5875 28172
rect 6178 28132 6184 28144
rect 6139 28104 6184 28132
rect 6178 28092 6184 28104
rect 6236 28092 6242 28144
rect 6288 28132 6316 28172
rect 7098 28160 7104 28172
rect 7156 28160 7162 28212
rect 10781 28203 10839 28209
rect 10781 28169 10793 28203
rect 10827 28200 10839 28203
rect 11054 28200 11060 28212
rect 10827 28172 11060 28200
rect 10827 28169 10839 28172
rect 10781 28163 10839 28169
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 14826 28200 14832 28212
rect 14787 28172 14832 28200
rect 14826 28160 14832 28172
rect 14884 28160 14890 28212
rect 16758 28160 16764 28212
rect 16816 28200 16822 28212
rect 17770 28200 17776 28212
rect 16816 28172 17776 28200
rect 16816 28160 16822 28172
rect 17770 28160 17776 28172
rect 17828 28160 17834 28212
rect 17954 28160 17960 28212
rect 18012 28200 18018 28212
rect 18230 28200 18236 28212
rect 18012 28172 18236 28200
rect 18012 28160 18018 28172
rect 18230 28160 18236 28172
rect 18288 28160 18294 28212
rect 18506 28160 18512 28212
rect 18564 28200 18570 28212
rect 20530 28200 20536 28212
rect 18564 28172 20536 28200
rect 18564 28160 18570 28172
rect 20530 28160 20536 28172
rect 20588 28160 20594 28212
rect 23753 28203 23811 28209
rect 23753 28169 23765 28203
rect 23799 28200 23811 28203
rect 24670 28200 24676 28212
rect 23799 28172 24676 28200
rect 23799 28169 23811 28172
rect 23753 28163 23811 28169
rect 24670 28160 24676 28172
rect 24728 28160 24734 28212
rect 28994 28160 29000 28212
rect 29052 28200 29058 28212
rect 29914 28200 29920 28212
rect 29052 28172 29920 28200
rect 29052 28160 29058 28172
rect 29914 28160 29920 28172
rect 29972 28160 29978 28212
rect 30282 28200 30288 28212
rect 30243 28172 30288 28200
rect 30282 28160 30288 28172
rect 30340 28160 30346 28212
rect 8294 28132 8300 28144
rect 6288 28104 8300 28132
rect 8294 28092 8300 28104
rect 8352 28092 8358 28144
rect 19426 28132 19432 28144
rect 14384 28104 19432 28132
rect 6454 28064 6460 28076
rect 5920 28036 6460 28064
rect 5920 28005 5948 28036
rect 6454 28024 6460 28036
rect 6512 28024 6518 28076
rect 7190 28024 7196 28076
rect 7248 28064 7254 28076
rect 7469 28067 7527 28073
rect 7469 28064 7481 28067
rect 7248 28036 7481 28064
rect 7248 28024 7254 28036
rect 7469 28033 7481 28036
rect 7515 28033 7527 28067
rect 7469 28027 7527 28033
rect 7558 28024 7564 28076
rect 7616 28064 7622 28076
rect 8202 28064 8208 28076
rect 7616 28036 8208 28064
rect 7616 28024 7622 28036
rect 8202 28024 8208 28036
rect 8260 28024 8266 28076
rect 13446 28024 13452 28076
rect 13504 28064 13510 28076
rect 14384 28073 14412 28104
rect 19426 28092 19432 28104
rect 19484 28132 19490 28144
rect 20070 28132 20076 28144
rect 19484 28104 20076 28132
rect 19484 28092 19490 28104
rect 20070 28092 20076 28104
rect 20128 28092 20134 28144
rect 20349 28135 20407 28141
rect 20349 28101 20361 28135
rect 20395 28132 20407 28135
rect 24394 28132 24400 28144
rect 20395 28104 24400 28132
rect 20395 28101 20407 28104
rect 20349 28095 20407 28101
rect 24394 28092 24400 28104
rect 24452 28092 24458 28144
rect 13541 28067 13599 28073
rect 13541 28064 13553 28067
rect 13504 28036 13553 28064
rect 13504 28024 13510 28036
rect 13541 28033 13553 28036
rect 13587 28064 13599 28067
rect 14369 28067 14427 28073
rect 14369 28064 14381 28067
rect 13587 28036 14381 28064
rect 13587 28033 13599 28036
rect 13541 28027 13599 28033
rect 14369 28033 14381 28036
rect 14415 28033 14427 28067
rect 14369 28027 14427 28033
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28064 15991 28067
rect 17037 28067 17095 28073
rect 17037 28064 17049 28067
rect 15979 28036 17049 28064
rect 15979 28033 15991 28036
rect 15933 28027 15991 28033
rect 17037 28033 17049 28036
rect 17083 28064 17095 28067
rect 17494 28064 17500 28076
rect 17083 28036 17500 28064
rect 17083 28033 17095 28036
rect 17037 28027 17095 28033
rect 17494 28024 17500 28036
rect 17552 28024 17558 28076
rect 17770 28024 17776 28076
rect 17828 28064 17834 28076
rect 17954 28064 17960 28076
rect 17828 28036 17960 28064
rect 17828 28024 17834 28036
rect 17954 28024 17960 28036
rect 18012 28024 18018 28076
rect 18046 28024 18052 28076
rect 18104 28064 18110 28076
rect 22281 28067 22339 28073
rect 18104 28036 18552 28064
rect 18104 28024 18110 28036
rect 5077 27999 5135 28005
rect 5077 27990 5089 27999
rect 5000 27965 5089 27990
rect 5123 27965 5135 27999
rect 5000 27962 5135 27965
rect 4246 27928 4252 27940
rect 2608 27900 4252 27928
rect 4246 27888 4252 27900
rect 4304 27888 4310 27940
rect 5000 27928 5028 27962
rect 5077 27959 5135 27962
rect 5537 27999 5595 28005
rect 5537 27965 5549 27999
rect 5583 27965 5595 27999
rect 5537 27959 5595 27965
rect 5721 27999 5779 28005
rect 5721 27965 5733 27999
rect 5767 27965 5779 27999
rect 5721 27959 5779 27965
rect 5816 27999 5875 28005
rect 5816 27965 5828 27999
rect 5862 27968 5875 27999
rect 5905 27999 5963 28005
rect 5862 27965 5874 27968
rect 5816 27959 5874 27965
rect 5905 27965 5917 27999
rect 5951 27965 5963 27999
rect 5905 27959 5963 27965
rect 5000 27900 5212 27928
rect 2774 27820 2780 27872
rect 2832 27860 2838 27872
rect 3234 27860 3240 27872
rect 2832 27832 3240 27860
rect 2832 27820 2838 27832
rect 3234 27820 3240 27832
rect 3292 27820 3298 27872
rect 4522 27820 4528 27872
rect 4580 27860 4586 27872
rect 4798 27860 4804 27872
rect 4580 27832 4804 27860
rect 4580 27820 4586 27832
rect 4798 27820 4804 27832
rect 4856 27820 4862 27872
rect 5184 27860 5212 27900
rect 5422 27888 5428 27940
rect 5480 27888 5486 27940
rect 5736 27928 5764 27959
rect 7098 27956 7104 28008
rect 7156 27996 7162 28008
rect 7282 27996 7288 28008
rect 7156 27968 7288 27996
rect 7156 27956 7162 27968
rect 7282 27956 7288 27968
rect 7340 27956 7346 28008
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27965 7711 27999
rect 7834 27996 7840 28008
rect 7795 27968 7840 27996
rect 7653 27959 7711 27965
rect 6454 27928 6460 27940
rect 5736 27900 6460 27928
rect 6454 27888 6460 27900
rect 6512 27928 6518 27940
rect 7668 27928 7696 27959
rect 7834 27956 7840 27968
rect 7892 27956 7898 28008
rect 9030 27956 9036 28008
rect 9088 27996 9094 28008
rect 9398 27996 9404 28008
rect 9088 27968 9404 27996
rect 9088 27956 9094 27968
rect 9398 27956 9404 27968
rect 9456 27956 9462 28008
rect 9668 27999 9726 28005
rect 9668 27965 9680 27999
rect 9714 27996 9726 27999
rect 10226 27996 10232 28008
rect 9714 27968 10232 27996
rect 9714 27965 9726 27968
rect 9668 27959 9726 27965
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 12342 27956 12348 28008
rect 12400 27996 12406 28008
rect 12618 27996 12624 28008
rect 12400 27968 12624 27996
rect 12400 27956 12406 27968
rect 12618 27956 12624 27968
rect 12676 27956 12682 28008
rect 14090 27996 14096 28008
rect 14051 27968 14096 27996
rect 14090 27956 14096 27968
rect 14148 27956 14154 28008
rect 14274 27996 14280 28008
rect 14235 27968 14280 27996
rect 14274 27956 14280 27968
rect 14332 27956 14338 28008
rect 14461 27999 14519 28005
rect 14461 27965 14473 27999
rect 14507 27965 14519 27999
rect 14642 27996 14648 28008
rect 14603 27968 14648 27996
rect 14461 27959 14519 27965
rect 6512 27900 7696 27928
rect 6512 27888 6518 27900
rect 11146 27888 11152 27940
rect 11204 27928 11210 27940
rect 11241 27931 11299 27937
rect 11241 27928 11253 27931
rect 11204 27900 11253 27928
rect 11204 27888 11210 27900
rect 11241 27897 11253 27900
rect 11287 27928 11299 27931
rect 12802 27928 12808 27940
rect 11287 27900 12808 27928
rect 11287 27897 11299 27900
rect 11241 27891 11299 27897
rect 12802 27888 12808 27900
rect 12860 27888 12866 27940
rect 12986 27928 12992 27940
rect 12947 27900 12992 27928
rect 12986 27888 12992 27900
rect 13044 27888 13050 27940
rect 13906 27888 13912 27940
rect 13964 27928 13970 27940
rect 14182 27928 14188 27940
rect 13964 27900 14188 27928
rect 13964 27888 13970 27900
rect 14182 27888 14188 27900
rect 14240 27928 14246 27940
rect 14476 27928 14504 27959
rect 14642 27956 14648 27968
rect 14700 27956 14706 28008
rect 15286 27956 15292 28008
rect 15344 27996 15350 28008
rect 16209 27999 16267 28005
rect 16209 27996 16221 27999
rect 15344 27968 16221 27996
rect 15344 27956 15350 27968
rect 16209 27965 16221 27968
rect 16255 27996 16267 27999
rect 16298 27996 16304 28008
rect 16255 27968 16304 27996
rect 16255 27965 16267 27968
rect 16209 27959 16267 27965
rect 16298 27956 16304 27968
rect 16356 27956 16362 28008
rect 17126 27956 17132 28008
rect 17184 27996 17190 28008
rect 17313 27999 17371 28005
rect 17313 27996 17325 27999
rect 17184 27968 17325 27996
rect 17184 27956 17190 27968
rect 17313 27965 17325 27968
rect 17359 27996 17371 27999
rect 18138 27996 18144 28008
rect 17359 27968 18144 27996
rect 17359 27965 17371 27968
rect 17313 27959 17371 27965
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 18524 28005 18552 28036
rect 22281 28033 22293 28067
rect 22327 28064 22339 28067
rect 22922 28064 22928 28076
rect 22327 28036 22928 28064
rect 22327 28033 22339 28036
rect 22281 28027 22339 28033
rect 22922 28024 22928 28036
rect 22980 28024 22986 28076
rect 23842 28064 23848 28076
rect 23492 28036 23848 28064
rect 18509 27999 18567 28005
rect 18509 27965 18521 27999
rect 18555 27965 18567 27999
rect 19610 27996 19616 28008
rect 19571 27968 19616 27996
rect 18509 27959 18567 27965
rect 19610 27956 19616 27968
rect 19668 27956 19674 28008
rect 19794 27996 19800 28008
rect 19755 27968 19800 27996
rect 19794 27956 19800 27968
rect 19852 27956 19858 28008
rect 20257 27999 20315 28005
rect 20257 27965 20269 27999
rect 20303 27965 20315 27999
rect 21174 27996 21180 28008
rect 21135 27968 21180 27996
rect 20257 27959 20315 27965
rect 17954 27928 17960 27940
rect 14240 27900 17960 27928
rect 14240 27888 14246 27900
rect 17954 27888 17960 27900
rect 18012 27888 18018 27940
rect 20272 27928 20300 27959
rect 21174 27956 21180 27968
rect 21232 27956 21238 28008
rect 21266 27956 21272 28008
rect 21324 27996 21330 28008
rect 21545 27999 21603 28005
rect 21545 27996 21557 27999
rect 21324 27968 21557 27996
rect 21324 27956 21330 27968
rect 21545 27965 21557 27968
rect 21591 27965 21603 27999
rect 22002 27996 22008 28008
rect 21963 27968 22008 27996
rect 21545 27959 21603 27965
rect 22002 27956 22008 27968
rect 22060 27996 22066 28008
rect 23492 27996 23520 28036
rect 23842 28024 23848 28036
rect 23900 28024 23906 28076
rect 24854 28064 24860 28076
rect 24815 28036 24860 28064
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 27522 28064 27528 28076
rect 27483 28036 27528 28064
rect 27522 28024 27528 28036
rect 27580 28024 27586 28076
rect 29086 28024 29092 28076
rect 29144 28064 29150 28076
rect 29144 28036 30144 28064
rect 29144 28024 29150 28036
rect 22060 27968 23520 27996
rect 23569 27999 23627 28005
rect 22060 27956 22066 27968
rect 23569 27965 23581 27999
rect 23615 27996 23627 27999
rect 23615 27968 24348 27996
rect 23615 27965 23627 27968
rect 23569 27959 23627 27965
rect 18064 27900 20300 27928
rect 22925 27931 22983 27937
rect 5440 27860 5468 27888
rect 5184 27832 5468 27860
rect 8202 27820 8208 27872
rect 8260 27860 8266 27872
rect 8389 27863 8447 27869
rect 8389 27860 8401 27863
rect 8260 27832 8401 27860
rect 8260 27820 8266 27832
rect 8389 27829 8401 27832
rect 8435 27860 8447 27863
rect 9490 27860 9496 27872
rect 8435 27832 9496 27860
rect 8435 27829 8447 27832
rect 8389 27823 8447 27829
rect 9490 27820 9496 27832
rect 9548 27820 9554 27872
rect 11790 27820 11796 27872
rect 11848 27860 11854 27872
rect 14734 27860 14740 27872
rect 11848 27832 14740 27860
rect 11848 27820 11854 27832
rect 14734 27820 14740 27832
rect 14792 27820 14798 27872
rect 15930 27820 15936 27872
rect 15988 27860 15994 27872
rect 18064 27860 18092 27900
rect 22925 27897 22937 27931
rect 22971 27928 22983 27931
rect 23658 27928 23664 27940
rect 22971 27900 23664 27928
rect 22971 27897 22983 27900
rect 22925 27891 22983 27897
rect 23658 27888 23664 27900
rect 23716 27888 23722 27940
rect 24320 27928 24348 27968
rect 24486 27956 24492 28008
rect 24544 27996 24550 28008
rect 25113 27999 25171 28005
rect 25113 27996 25125 27999
rect 24544 27968 25125 27996
rect 24544 27956 24550 27968
rect 25113 27965 25125 27968
rect 25159 27965 25171 27999
rect 25113 27959 25171 27965
rect 27249 27999 27307 28005
rect 27249 27965 27261 27999
rect 27295 27965 27307 27999
rect 27249 27959 27307 27965
rect 27264 27928 27292 27959
rect 27614 27956 27620 28008
rect 27672 27996 27678 28008
rect 28537 27999 28595 28005
rect 28537 27996 28549 27999
rect 27672 27968 28549 27996
rect 27672 27956 27678 27968
rect 28537 27965 28549 27968
rect 28583 27965 28595 27999
rect 28537 27959 28595 27965
rect 28626 27956 28632 28008
rect 28684 27996 28690 28008
rect 29546 27996 29552 28008
rect 28684 27968 29552 27996
rect 28684 27956 28690 27968
rect 29546 27956 29552 27968
rect 29604 27956 29610 28008
rect 29733 27999 29791 28005
rect 29733 27965 29745 27999
rect 29779 27965 29791 27999
rect 29733 27959 29791 27965
rect 29825 27999 29883 28005
rect 29825 27965 29837 27999
rect 29871 27965 29883 27999
rect 29825 27959 29883 27965
rect 24320 27900 26464 27928
rect 27264 27900 27660 27928
rect 26436 27872 26464 27900
rect 27632 27872 27660 27900
rect 15988 27832 18092 27860
rect 18601 27863 18659 27869
rect 15988 27820 15994 27832
rect 18601 27829 18613 27863
rect 18647 27860 18659 27863
rect 19242 27860 19248 27872
rect 18647 27832 19248 27860
rect 18647 27829 18659 27832
rect 18601 27823 18659 27829
rect 19242 27820 19248 27832
rect 19300 27820 19306 27872
rect 23017 27863 23075 27869
rect 23017 27829 23029 27863
rect 23063 27860 23075 27863
rect 25682 27860 25688 27872
rect 23063 27832 25688 27860
rect 23063 27829 23075 27832
rect 23017 27823 23075 27829
rect 25682 27820 25688 27832
rect 25740 27820 25746 27872
rect 25774 27820 25780 27872
rect 25832 27860 25838 27872
rect 26237 27863 26295 27869
rect 26237 27860 26249 27863
rect 25832 27832 26249 27860
rect 25832 27820 25838 27832
rect 26237 27829 26249 27832
rect 26283 27829 26295 27863
rect 26237 27823 26295 27829
rect 26418 27820 26424 27872
rect 26476 27860 26482 27872
rect 26602 27860 26608 27872
rect 26476 27832 26608 27860
rect 26476 27820 26482 27832
rect 26602 27820 26608 27832
rect 26660 27860 26666 27872
rect 26697 27863 26755 27869
rect 26697 27860 26709 27863
rect 26660 27832 26709 27860
rect 26660 27820 26666 27832
rect 26697 27829 26709 27832
rect 26743 27829 26755 27863
rect 26697 27823 26755 27829
rect 27614 27820 27620 27872
rect 27672 27820 27678 27872
rect 28258 27820 28264 27872
rect 28316 27860 28322 27872
rect 28629 27863 28687 27869
rect 28629 27860 28641 27863
rect 28316 27832 28641 27860
rect 28316 27820 28322 27832
rect 28629 27829 28641 27832
rect 28675 27829 28687 27863
rect 28629 27823 28687 27829
rect 28810 27820 28816 27872
rect 28868 27860 28874 27872
rect 29748 27860 29776 27959
rect 29840 27928 29868 27959
rect 29914 27956 29920 28008
rect 29972 27996 29978 28008
rect 30116 28005 30144 28036
rect 30101 27999 30159 28005
rect 29972 27968 30017 27996
rect 29972 27956 29978 27968
rect 30101 27965 30113 27999
rect 30147 27965 30159 27999
rect 31110 27996 31116 28008
rect 31071 27968 31116 27996
rect 30101 27959 30159 27965
rect 31110 27956 31116 27968
rect 31168 27956 31174 28008
rect 30006 27928 30012 27940
rect 29840 27900 30012 27928
rect 30006 27888 30012 27900
rect 30064 27888 30070 27940
rect 28868 27832 29776 27860
rect 31297 27863 31355 27869
rect 28868 27820 28874 27832
rect 31297 27829 31309 27863
rect 31343 27860 31355 27863
rect 31343 27832 32076 27860
rect 31343 27829 31355 27832
rect 31297 27823 31355 27829
rect 1104 27770 32016 27792
rect 1104 27718 11253 27770
rect 11305 27718 11317 27770
rect 11369 27718 11381 27770
rect 11433 27718 11445 27770
rect 11497 27718 11509 27770
rect 11561 27718 21557 27770
rect 21609 27718 21621 27770
rect 21673 27718 21685 27770
rect 21737 27718 21749 27770
rect 21801 27718 21813 27770
rect 21865 27718 32016 27770
rect 1104 27696 32016 27718
rect 1486 27616 1492 27668
rect 1544 27616 1550 27668
rect 2225 27659 2283 27665
rect 2225 27625 2237 27659
rect 2271 27656 2283 27659
rect 2682 27656 2688 27668
rect 2271 27628 2688 27656
rect 2271 27625 2283 27628
rect 2225 27619 2283 27625
rect 2682 27616 2688 27628
rect 2740 27616 2746 27668
rect 7098 27656 7104 27668
rect 6288 27628 7104 27656
rect 0 27588 800 27602
rect 1504 27588 1532 27616
rect 0 27560 1532 27588
rect 0 27546 800 27560
rect 1578 27548 1584 27600
rect 1636 27588 1642 27600
rect 1636 27560 1681 27588
rect 1636 27548 1642 27560
rect 1946 27548 1952 27600
rect 2004 27588 2010 27600
rect 2774 27588 2780 27600
rect 2004 27560 2780 27588
rect 2004 27548 2010 27560
rect 2774 27548 2780 27560
rect 2832 27548 2838 27600
rect 3602 27548 3608 27600
rect 3660 27588 3666 27600
rect 5537 27591 5595 27597
rect 3660 27560 3924 27588
rect 3660 27548 3666 27560
rect 3896 27532 3924 27560
rect 5537 27557 5549 27591
rect 5583 27588 5595 27591
rect 5994 27588 6000 27600
rect 5583 27560 6000 27588
rect 5583 27557 5595 27560
rect 5537 27551 5595 27557
rect 5994 27548 6000 27560
rect 6052 27548 6058 27600
rect 1489 27523 1547 27529
rect 1489 27489 1501 27523
rect 1535 27489 1547 27523
rect 1489 27483 1547 27489
rect 1394 27412 1400 27464
rect 1452 27452 1458 27464
rect 1504 27452 1532 27483
rect 2038 27480 2044 27532
rect 2096 27520 2102 27532
rect 2133 27523 2191 27529
rect 2133 27520 2145 27523
rect 2096 27492 2145 27520
rect 2096 27480 2102 27492
rect 2133 27489 2145 27492
rect 2179 27489 2191 27523
rect 2133 27483 2191 27489
rect 2222 27480 2228 27532
rect 2280 27520 2286 27532
rect 2317 27523 2375 27529
rect 2317 27520 2329 27523
rect 2280 27492 2329 27520
rect 2280 27480 2286 27492
rect 2317 27489 2329 27492
rect 2363 27489 2375 27523
rect 3326 27520 3332 27532
rect 3287 27492 3332 27520
rect 2317 27483 2375 27489
rect 3326 27480 3332 27492
rect 3384 27480 3390 27532
rect 3510 27520 3516 27532
rect 3471 27492 3516 27520
rect 3510 27480 3516 27492
rect 3568 27480 3574 27532
rect 3878 27520 3884 27532
rect 3791 27492 3884 27520
rect 3878 27480 3884 27492
rect 3936 27480 3942 27532
rect 4890 27480 4896 27532
rect 4948 27520 4954 27532
rect 4985 27523 5043 27529
rect 4985 27520 4997 27523
rect 4948 27492 4997 27520
rect 4948 27480 4954 27492
rect 4985 27489 4997 27492
rect 5031 27489 5043 27523
rect 4985 27483 5043 27489
rect 5077 27523 5135 27529
rect 5077 27489 5089 27523
rect 5123 27520 5135 27523
rect 5813 27523 5871 27529
rect 5123 27492 5488 27520
rect 5123 27489 5135 27492
rect 5077 27483 5135 27489
rect 2498 27452 2504 27464
rect 1452 27424 2504 27452
rect 1452 27412 1458 27424
rect 2498 27412 2504 27424
rect 2556 27412 2562 27464
rect 2869 27455 2927 27461
rect 2869 27421 2881 27455
rect 2915 27452 2927 27455
rect 3234 27452 3240 27464
rect 2915 27424 3240 27452
rect 2915 27421 2927 27424
rect 2869 27415 2927 27421
rect 3234 27412 3240 27424
rect 3292 27452 3298 27464
rect 3605 27455 3663 27461
rect 3605 27452 3617 27455
rect 3292 27424 3617 27452
rect 3292 27412 3298 27424
rect 3605 27421 3617 27424
rect 3651 27421 3663 27455
rect 3605 27415 3663 27421
rect 3697 27455 3755 27461
rect 3697 27421 3709 27455
rect 3743 27452 3755 27455
rect 4154 27452 4160 27464
rect 3743 27424 4160 27452
rect 3743 27421 3755 27424
rect 3697 27415 3755 27421
rect 4154 27412 4160 27424
rect 4212 27412 4218 27464
rect 4338 27412 4344 27464
rect 4396 27452 4402 27464
rect 4396 27424 4936 27452
rect 4396 27412 4402 27424
rect 1670 27344 1676 27396
rect 1728 27384 1734 27396
rect 4706 27384 4712 27396
rect 1728 27356 4712 27384
rect 1728 27344 1734 27356
rect 4706 27344 4712 27356
rect 4764 27344 4770 27396
rect 4908 27328 4936 27424
rect 5460 27384 5488 27492
rect 5813 27489 5825 27523
rect 5859 27520 5871 27523
rect 6288 27520 6316 27628
rect 7098 27616 7104 27628
rect 7156 27656 7162 27668
rect 7156 27628 9628 27656
rect 7156 27616 7162 27628
rect 6457 27591 6515 27597
rect 6457 27557 6469 27591
rect 6503 27588 6515 27591
rect 6638 27588 6644 27600
rect 6503 27560 6644 27588
rect 6503 27557 6515 27560
rect 6457 27551 6515 27557
rect 6638 27548 6644 27560
rect 6696 27548 6702 27600
rect 7742 27588 7748 27600
rect 7300 27560 7748 27588
rect 5859 27492 6316 27520
rect 6365 27523 6423 27529
rect 5859 27489 5871 27492
rect 5813 27483 5871 27489
rect 6365 27489 6377 27523
rect 6411 27520 6423 27523
rect 6549 27523 6607 27529
rect 6411 27492 6500 27520
rect 6411 27489 6423 27492
rect 6365 27483 6423 27489
rect 6472 27464 6500 27492
rect 6549 27489 6561 27523
rect 6595 27520 6607 27523
rect 6914 27520 6920 27532
rect 6595 27492 6920 27520
rect 6595 27489 6607 27492
rect 6549 27483 6607 27489
rect 5537 27455 5595 27461
rect 5537 27421 5549 27455
rect 5583 27452 5595 27455
rect 6270 27452 6276 27464
rect 5583 27424 6276 27452
rect 5583 27421 5595 27424
rect 5537 27415 5595 27421
rect 6270 27412 6276 27424
rect 6328 27412 6334 27464
rect 6454 27412 6460 27464
rect 6512 27412 6518 27464
rect 6564 27384 6592 27483
rect 6914 27480 6920 27492
rect 6972 27480 6978 27532
rect 7300 27529 7328 27560
rect 7742 27548 7748 27560
rect 7800 27548 7806 27600
rect 8021 27591 8079 27597
rect 8021 27557 8033 27591
rect 8067 27588 8079 27591
rect 8726 27591 8784 27597
rect 8726 27588 8738 27591
rect 8067 27560 8738 27588
rect 8067 27557 8079 27560
rect 8021 27551 8079 27557
rect 8726 27557 8738 27560
rect 8772 27557 8784 27591
rect 9600 27588 9628 27628
rect 9674 27616 9680 27668
rect 9732 27656 9738 27668
rect 14737 27659 14795 27665
rect 9732 27628 14688 27656
rect 9732 27616 9738 27628
rect 10321 27591 10379 27597
rect 10321 27588 10333 27591
rect 9600 27560 10333 27588
rect 8726 27551 8784 27557
rect 10321 27557 10333 27560
rect 10367 27557 10379 27591
rect 10321 27551 10379 27557
rect 10962 27548 10968 27600
rect 11020 27588 11026 27600
rect 11238 27588 11244 27600
rect 11020 27560 11244 27588
rect 11020 27548 11026 27560
rect 11238 27548 11244 27560
rect 11296 27548 11302 27600
rect 14553 27591 14611 27597
rect 11900 27560 12434 27588
rect 7285 27523 7343 27529
rect 7285 27489 7297 27523
rect 7331 27489 7343 27523
rect 7285 27483 7343 27489
rect 7469 27523 7527 27529
rect 7469 27489 7481 27523
rect 7515 27520 7527 27523
rect 7515 27492 7788 27520
rect 7515 27489 7527 27492
rect 7469 27483 7527 27489
rect 7558 27452 7564 27464
rect 7519 27424 7564 27452
rect 7558 27412 7564 27424
rect 7616 27412 7622 27464
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27421 7711 27455
rect 7653 27415 7711 27421
rect 5460 27356 6592 27384
rect 7190 27344 7196 27396
rect 7248 27384 7254 27396
rect 7668 27384 7696 27415
rect 7248 27356 7696 27384
rect 7760 27384 7788 27492
rect 7834 27480 7840 27532
rect 7892 27520 7898 27532
rect 7892 27492 7937 27520
rect 7892 27480 7898 27492
rect 8386 27480 8392 27532
rect 8444 27520 8450 27532
rect 8481 27523 8539 27529
rect 8481 27520 8493 27523
rect 8444 27492 8493 27520
rect 8444 27480 8450 27492
rect 8481 27489 8493 27492
rect 8527 27489 8539 27523
rect 8481 27483 8539 27489
rect 8570 27480 8576 27532
rect 8628 27520 8634 27532
rect 10226 27520 10232 27532
rect 8628 27492 10232 27520
rect 8628 27480 8634 27492
rect 10226 27480 10232 27492
rect 10284 27480 10290 27532
rect 11900 27529 11928 27560
rect 11885 27523 11943 27529
rect 11885 27489 11897 27523
rect 11931 27489 11943 27523
rect 11885 27483 11943 27489
rect 11974 27480 11980 27532
rect 12032 27520 12038 27532
rect 12141 27523 12199 27529
rect 12141 27520 12153 27523
rect 12032 27492 12153 27520
rect 12032 27480 12038 27492
rect 12141 27489 12153 27492
rect 12187 27489 12199 27523
rect 12406 27520 12434 27560
rect 14553 27557 14565 27591
rect 14599 27557 14611 27591
rect 14660 27588 14688 27628
rect 14737 27625 14749 27659
rect 14783 27656 14795 27659
rect 15010 27656 15016 27668
rect 14783 27628 15016 27656
rect 14783 27625 14795 27628
rect 14737 27619 14795 27625
rect 15010 27616 15016 27628
rect 15068 27616 15074 27668
rect 15120 27628 18736 27656
rect 15120 27588 15148 27628
rect 14660 27560 15148 27588
rect 15764 27560 16574 27588
rect 14553 27551 14611 27557
rect 12986 27520 12992 27532
rect 12406 27492 12992 27520
rect 12141 27483 12199 27489
rect 12986 27480 12992 27492
rect 13044 27480 13050 27532
rect 14090 27480 14096 27532
rect 14148 27520 14154 27532
rect 14185 27523 14243 27529
rect 14185 27520 14197 27523
rect 14148 27492 14197 27520
rect 14148 27480 14154 27492
rect 14185 27489 14197 27492
rect 14231 27489 14243 27523
rect 14568 27520 14596 27551
rect 14642 27520 14648 27532
rect 14568 27492 14648 27520
rect 14185 27483 14243 27489
rect 14642 27480 14648 27492
rect 14700 27480 14706 27532
rect 15654 27520 15660 27532
rect 15615 27492 15660 27520
rect 15654 27480 15660 27492
rect 15712 27480 15718 27532
rect 8588 27452 8616 27480
rect 8496 27424 8616 27452
rect 8496 27384 8524 27424
rect 7760 27356 8524 27384
rect 7248 27344 7254 27356
rect 9490 27344 9496 27396
rect 9548 27384 9554 27396
rect 15764 27384 15792 27560
rect 15930 27452 15936 27464
rect 15891 27424 15936 27452
rect 15930 27412 15936 27424
rect 15988 27412 15994 27464
rect 16546 27452 16574 27560
rect 17678 27548 17684 27600
rect 17736 27588 17742 27600
rect 18598 27588 18604 27600
rect 17736 27560 18276 27588
rect 18559 27560 18604 27588
rect 17736 27548 17742 27560
rect 16850 27520 16856 27532
rect 16811 27492 16856 27520
rect 16850 27480 16856 27492
rect 16908 27480 16914 27532
rect 17126 27520 17132 27532
rect 17087 27492 17132 27520
rect 17126 27480 17132 27492
rect 17184 27480 17190 27532
rect 17221 27530 17279 27535
rect 17310 27530 17316 27532
rect 17221 27529 17316 27530
rect 17221 27495 17233 27529
rect 17267 27502 17316 27529
rect 17267 27495 17279 27502
rect 17221 27489 17279 27495
rect 17310 27480 17316 27502
rect 17368 27480 17374 27532
rect 17405 27523 17463 27529
rect 17405 27489 17417 27523
rect 17451 27518 17463 27523
rect 17770 27520 17776 27532
rect 17595 27518 17776 27520
rect 17451 27492 17776 27518
rect 17451 27490 17623 27492
rect 17451 27489 17463 27490
rect 17405 27483 17463 27489
rect 17770 27480 17776 27492
rect 17828 27520 17834 27532
rect 17865 27523 17923 27529
rect 17865 27520 17877 27523
rect 17828 27492 17877 27520
rect 17828 27480 17834 27492
rect 17865 27489 17877 27492
rect 17911 27489 17923 27523
rect 18046 27520 18052 27532
rect 18007 27492 18052 27520
rect 17865 27483 17923 27489
rect 18046 27480 18052 27492
rect 18104 27480 18110 27532
rect 18248 27529 18276 27560
rect 18598 27548 18604 27560
rect 18656 27548 18662 27600
rect 18708 27588 18736 27628
rect 18782 27616 18788 27668
rect 18840 27656 18846 27668
rect 19518 27656 19524 27668
rect 18840 27628 19524 27656
rect 18840 27616 18846 27628
rect 19518 27616 19524 27628
rect 19576 27616 19582 27668
rect 19610 27616 19616 27668
rect 19668 27656 19674 27668
rect 19797 27659 19855 27665
rect 19797 27656 19809 27659
rect 19668 27628 19809 27656
rect 19668 27616 19674 27628
rect 19797 27625 19809 27628
rect 19843 27625 19855 27659
rect 21174 27656 21180 27668
rect 21135 27628 21180 27656
rect 19797 27619 19855 27625
rect 21174 27616 21180 27628
rect 21232 27616 21238 27668
rect 24213 27659 24271 27665
rect 21284 27628 23244 27656
rect 18966 27588 18972 27600
rect 18708 27560 18972 27588
rect 18966 27548 18972 27560
rect 19024 27548 19030 27600
rect 19150 27548 19156 27600
rect 19208 27588 19214 27600
rect 19208 27560 19656 27588
rect 19208 27548 19214 27560
rect 18233 27523 18291 27529
rect 18233 27489 18245 27523
rect 18279 27489 18291 27523
rect 18233 27483 18291 27489
rect 18417 27523 18475 27529
rect 18417 27489 18429 27523
rect 18463 27520 18475 27523
rect 19058 27520 19064 27532
rect 18463 27492 19064 27520
rect 18463 27489 18475 27492
rect 18417 27483 18475 27489
rect 19058 27480 19064 27492
rect 19116 27480 19122 27532
rect 19242 27520 19248 27532
rect 19203 27492 19248 27520
rect 19242 27480 19248 27492
rect 19300 27480 19306 27532
rect 19628 27529 19656 27560
rect 19978 27548 19984 27600
rect 20036 27588 20042 27600
rect 21284 27588 21312 27628
rect 20036 27560 21312 27588
rect 23017 27591 23075 27597
rect 20036 27548 20042 27560
rect 23017 27557 23029 27591
rect 23063 27588 23075 27591
rect 23106 27588 23112 27600
rect 23063 27560 23112 27588
rect 23063 27557 23075 27560
rect 23017 27551 23075 27557
rect 19337 27523 19395 27529
rect 19337 27489 19349 27523
rect 19383 27520 19395 27523
rect 19613 27523 19671 27529
rect 19383 27492 19564 27520
rect 19383 27489 19395 27492
rect 19337 27483 19395 27489
rect 17037 27455 17095 27461
rect 16546 27424 16896 27452
rect 9548 27356 11008 27384
rect 9548 27344 9554 27356
rect 1302 27276 1308 27328
rect 1360 27316 1366 27328
rect 3786 27316 3792 27328
rect 1360 27288 3792 27316
rect 1360 27276 1366 27288
rect 3786 27276 3792 27288
rect 3844 27276 3850 27328
rect 4065 27319 4123 27325
rect 4065 27285 4077 27319
rect 4111 27316 4123 27319
rect 4522 27316 4528 27328
rect 4111 27288 4528 27316
rect 4111 27285 4123 27288
rect 4065 27279 4123 27285
rect 4522 27276 4528 27288
rect 4580 27276 4586 27328
rect 4890 27276 4896 27328
rect 4948 27316 4954 27328
rect 5721 27319 5779 27325
rect 5721 27316 5733 27319
rect 4948 27288 5733 27316
rect 4948 27276 4954 27288
rect 5721 27285 5733 27288
rect 5767 27285 5779 27319
rect 5721 27279 5779 27285
rect 8754 27276 8760 27328
rect 8812 27316 8818 27328
rect 10980 27325 11008 27356
rect 12820 27356 15792 27384
rect 9861 27319 9919 27325
rect 9861 27316 9873 27319
rect 8812 27288 9873 27316
rect 8812 27276 8818 27288
rect 9861 27285 9873 27288
rect 9907 27285 9919 27319
rect 9861 27279 9919 27285
rect 10965 27319 11023 27325
rect 10965 27285 10977 27319
rect 11011 27316 11023 27319
rect 12820 27316 12848 27356
rect 16206 27344 16212 27396
rect 16264 27384 16270 27396
rect 16868 27384 16896 27424
rect 17037 27421 17049 27455
rect 17083 27452 17095 27455
rect 17678 27452 17684 27464
rect 17083 27424 17684 27452
rect 17083 27421 17095 27424
rect 17037 27415 17095 27421
rect 17678 27412 17684 27424
rect 17736 27412 17742 27464
rect 18138 27452 18144 27464
rect 18099 27424 18144 27452
rect 18138 27412 18144 27424
rect 18196 27412 18202 27464
rect 19426 27452 19432 27464
rect 19387 27424 19432 27452
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 19536 27452 19564 27492
rect 19613 27489 19625 27523
rect 19659 27489 19671 27523
rect 19613 27483 19671 27489
rect 20162 27480 20168 27532
rect 20220 27520 20226 27532
rect 20441 27523 20499 27529
rect 20441 27520 20453 27523
rect 20220 27492 20453 27520
rect 20220 27480 20226 27492
rect 20441 27489 20453 27492
rect 20487 27489 20499 27523
rect 20622 27520 20628 27532
rect 20583 27492 20628 27520
rect 20441 27483 20499 27489
rect 20622 27480 20628 27492
rect 20680 27480 20686 27532
rect 20993 27523 21051 27529
rect 20993 27489 21005 27523
rect 21039 27520 21051 27523
rect 22094 27520 22100 27532
rect 21039 27492 22100 27520
rect 21039 27489 21051 27492
rect 20993 27483 21051 27489
rect 22094 27480 22100 27492
rect 22152 27480 22158 27532
rect 22281 27523 22339 27529
rect 22281 27489 22293 27523
rect 22327 27520 22339 27523
rect 23032 27520 23060 27551
rect 23106 27548 23112 27560
rect 23164 27548 23170 27600
rect 23216 27588 23244 27628
rect 24213 27625 24225 27659
rect 24259 27656 24271 27659
rect 24394 27656 24400 27668
rect 24259 27628 24400 27656
rect 24259 27625 24271 27628
rect 24213 27619 24271 27625
rect 24394 27616 24400 27628
rect 24452 27616 24458 27668
rect 27522 27656 27528 27668
rect 24504 27628 27528 27656
rect 24302 27588 24308 27600
rect 23216 27560 23879 27588
rect 24263 27560 24308 27588
rect 22327 27492 23060 27520
rect 23385 27523 23443 27529
rect 22327 27489 22339 27492
rect 22281 27483 22339 27489
rect 23385 27489 23397 27523
rect 23431 27520 23443 27523
rect 23750 27520 23756 27532
rect 23431 27492 23756 27520
rect 23431 27489 23443 27492
rect 23385 27483 23443 27489
rect 19978 27452 19984 27464
rect 19536 27424 19984 27452
rect 19978 27412 19984 27424
rect 20036 27412 20042 27464
rect 20070 27412 20076 27464
rect 20128 27452 20134 27464
rect 20717 27455 20775 27461
rect 20717 27452 20729 27455
rect 20128 27424 20729 27452
rect 20128 27412 20134 27424
rect 20717 27421 20729 27424
rect 20763 27421 20775 27455
rect 20717 27415 20775 27421
rect 20806 27412 20812 27464
rect 20864 27452 20870 27464
rect 22738 27452 22744 27464
rect 20864 27424 22744 27452
rect 20864 27412 20870 27424
rect 22738 27412 22744 27424
rect 22796 27412 22802 27464
rect 22922 27412 22928 27464
rect 22980 27452 22986 27464
rect 23400 27452 23428 27483
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 23851 27520 23879 27560
rect 24302 27548 24308 27560
rect 24360 27548 24366 27600
rect 24504 27520 24532 27628
rect 27522 27616 27528 27628
rect 27580 27616 27586 27668
rect 31110 27616 31116 27668
rect 31168 27656 31174 27668
rect 31297 27659 31355 27665
rect 31297 27656 31309 27659
rect 31168 27628 31309 27656
rect 31168 27616 31174 27628
rect 31297 27625 31309 27628
rect 31343 27625 31355 27659
rect 31297 27619 31355 27625
rect 24762 27548 24768 27600
rect 24820 27588 24826 27600
rect 25222 27588 25228 27600
rect 24820 27560 25228 27588
rect 24820 27548 24826 27560
rect 25222 27548 25228 27560
rect 25280 27588 25286 27600
rect 25406 27588 25412 27600
rect 25280 27560 25412 27588
rect 25280 27548 25286 27560
rect 25406 27548 25412 27560
rect 25464 27548 25470 27600
rect 26142 27548 26148 27600
rect 26200 27548 26206 27600
rect 27801 27591 27859 27597
rect 27801 27557 27813 27591
rect 27847 27588 27859 27591
rect 28994 27588 29000 27600
rect 27847 27560 29000 27588
rect 27847 27557 27859 27560
rect 27801 27551 27859 27557
rect 28994 27548 29000 27560
rect 29052 27548 29058 27600
rect 32048 27588 32076 27832
rect 32320 27588 33120 27602
rect 32048 27560 33120 27588
rect 23851 27492 24532 27520
rect 25869 27523 25927 27529
rect 25869 27489 25881 27523
rect 25915 27520 25927 27523
rect 26160 27520 26188 27548
rect 32320 27546 33120 27560
rect 25915 27492 26188 27520
rect 27617 27523 27675 27529
rect 25915 27489 25927 27492
rect 25869 27483 25927 27489
rect 27617 27489 27629 27523
rect 27663 27489 27675 27523
rect 27617 27483 27675 27489
rect 28813 27523 28871 27529
rect 28813 27489 28825 27523
rect 28859 27520 28871 27523
rect 28902 27520 28908 27532
rect 28859 27492 28908 27520
rect 28859 27489 28871 27492
rect 28813 27483 28871 27489
rect 22980 27424 23428 27452
rect 22980 27412 22986 27424
rect 25682 27412 25688 27464
rect 25740 27452 25746 27464
rect 26145 27455 26203 27461
rect 26145 27452 26157 27455
rect 25740 27424 26157 27452
rect 25740 27412 25746 27424
rect 26145 27421 26157 27424
rect 26191 27452 26203 27455
rect 27632 27452 27660 27483
rect 28902 27480 28908 27492
rect 28960 27520 28966 27532
rect 29546 27520 29552 27532
rect 28960 27492 29224 27520
rect 29507 27492 29552 27520
rect 28960 27480 28966 27492
rect 27982 27452 27988 27464
rect 26191 27424 27988 27452
rect 26191 27421 26203 27424
rect 26145 27415 26203 27421
rect 27982 27412 27988 27424
rect 28040 27412 28046 27464
rect 28718 27412 28724 27464
rect 28776 27452 28782 27464
rect 29089 27455 29147 27461
rect 29089 27452 29101 27455
rect 28776 27424 29101 27452
rect 28776 27412 28782 27424
rect 29089 27421 29101 27424
rect 29135 27421 29147 27455
rect 29196 27452 29224 27492
rect 29546 27480 29552 27492
rect 29604 27480 29610 27532
rect 29730 27520 29736 27532
rect 29691 27492 29736 27520
rect 29730 27480 29736 27492
rect 29788 27480 29794 27532
rect 30006 27520 30012 27532
rect 29840 27492 30012 27520
rect 29638 27452 29644 27464
rect 29196 27424 29644 27452
rect 29089 27415 29147 27421
rect 29638 27412 29644 27424
rect 29696 27452 29702 27464
rect 29840 27461 29868 27492
rect 30006 27480 30012 27492
rect 30064 27480 30070 27532
rect 30101 27523 30159 27529
rect 30101 27489 30113 27523
rect 30147 27520 30159 27523
rect 30466 27520 30472 27532
rect 30147 27492 30472 27520
rect 30147 27489 30159 27492
rect 30101 27483 30159 27489
rect 30466 27480 30472 27492
rect 30524 27480 30530 27532
rect 31113 27523 31171 27529
rect 31113 27489 31125 27523
rect 31159 27520 31171 27523
rect 31294 27520 31300 27532
rect 31159 27492 31300 27520
rect 31159 27489 31171 27492
rect 31113 27483 31171 27489
rect 31294 27480 31300 27492
rect 31352 27480 31358 27532
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 29696 27424 29837 27452
rect 29696 27412 29702 27424
rect 29825 27421 29837 27424
rect 29871 27421 29883 27455
rect 29825 27415 29883 27421
rect 29914 27412 29920 27464
rect 29972 27452 29978 27464
rect 29972 27424 30017 27452
rect 29972 27412 29978 27424
rect 23566 27384 23572 27396
rect 16264 27356 16804 27384
rect 16868 27356 23572 27384
rect 16264 27344 16270 27356
rect 11011 27288 12848 27316
rect 11011 27285 11023 27288
rect 10965 27279 11023 27285
rect 13262 27276 13268 27328
rect 13320 27316 13326 27328
rect 13320 27288 13365 27316
rect 13320 27276 13326 27288
rect 14274 27276 14280 27328
rect 14332 27316 14338 27328
rect 14553 27319 14611 27325
rect 14553 27316 14565 27319
rect 14332 27288 14565 27316
rect 14332 27276 14338 27288
rect 14553 27285 14565 27288
rect 14599 27285 14611 27319
rect 14553 27279 14611 27285
rect 16298 27276 16304 27328
rect 16356 27316 16362 27328
rect 16669 27319 16727 27325
rect 16669 27316 16681 27319
rect 16356 27288 16681 27316
rect 16356 27276 16362 27288
rect 16669 27285 16681 27288
rect 16715 27285 16727 27319
rect 16776 27316 16804 27356
rect 23566 27344 23572 27356
rect 23624 27344 23630 27396
rect 24302 27344 24308 27396
rect 24360 27384 24366 27396
rect 26973 27387 27031 27393
rect 26973 27384 26985 27387
rect 24360 27356 26985 27384
rect 24360 27344 24366 27356
rect 26973 27353 26985 27356
rect 27019 27353 27031 27387
rect 26973 27347 27031 27353
rect 27246 27344 27252 27396
rect 27304 27384 27310 27396
rect 30834 27384 30840 27396
rect 27304 27356 30840 27384
rect 27304 27344 27310 27356
rect 30834 27344 30840 27356
rect 30892 27344 30898 27396
rect 17310 27316 17316 27328
rect 16776 27288 17316 27316
rect 16669 27279 16727 27285
rect 17310 27276 17316 27288
rect 17368 27316 17374 27328
rect 18598 27316 18604 27328
rect 17368 27288 18604 27316
rect 17368 27276 17374 27288
rect 18598 27276 18604 27288
rect 18656 27276 18662 27328
rect 22465 27319 22523 27325
rect 22465 27285 22477 27319
rect 22511 27316 22523 27319
rect 27614 27316 27620 27328
rect 22511 27288 27620 27316
rect 22511 27285 22523 27288
rect 22465 27279 22523 27285
rect 27614 27276 27620 27288
rect 27672 27316 27678 27328
rect 28166 27316 28172 27328
rect 27672 27288 28172 27316
rect 27672 27276 27678 27288
rect 28166 27276 28172 27288
rect 28224 27316 28230 27328
rect 28718 27316 28724 27328
rect 28224 27288 28724 27316
rect 28224 27276 28230 27288
rect 28718 27276 28724 27288
rect 28776 27276 28782 27328
rect 30285 27319 30343 27325
rect 30285 27285 30297 27319
rect 30331 27316 30343 27319
rect 30926 27316 30932 27328
rect 30331 27288 30932 27316
rect 30331 27285 30343 27288
rect 30285 27279 30343 27285
rect 30926 27276 30932 27288
rect 30984 27276 30990 27328
rect 1104 27226 32016 27248
rect 1104 27174 6102 27226
rect 6154 27174 6166 27226
rect 6218 27174 6230 27226
rect 6282 27174 6294 27226
rect 6346 27174 6358 27226
rect 6410 27174 16405 27226
rect 16457 27174 16469 27226
rect 16521 27174 16533 27226
rect 16585 27174 16597 27226
rect 16649 27174 16661 27226
rect 16713 27174 26709 27226
rect 26761 27174 26773 27226
rect 26825 27174 26837 27226
rect 26889 27174 26901 27226
rect 26953 27174 26965 27226
rect 27017 27174 32016 27226
rect 1104 27152 32016 27174
rect 1762 27112 1768 27124
rect 1723 27084 1768 27112
rect 1762 27072 1768 27084
rect 1820 27072 1826 27124
rect 4246 27072 4252 27124
rect 4304 27112 4310 27124
rect 6273 27115 6331 27121
rect 4304 27084 4844 27112
rect 4304 27072 4310 27084
rect 4062 27004 4068 27056
rect 4120 27044 4126 27056
rect 4706 27044 4712 27056
rect 4120 27016 4712 27044
rect 4120 27004 4126 27016
rect 4706 27004 4712 27016
rect 4764 27004 4770 27056
rect 4816 26976 4844 27084
rect 6273 27081 6285 27115
rect 6319 27112 6331 27115
rect 6730 27112 6736 27124
rect 6319 27084 6736 27112
rect 6319 27081 6331 27084
rect 6273 27075 6331 27081
rect 6730 27072 6736 27084
rect 6788 27112 6794 27124
rect 8386 27112 8392 27124
rect 6788 27084 8392 27112
rect 6788 27072 6794 27084
rect 8386 27072 8392 27084
rect 8444 27072 8450 27124
rect 10226 27072 10232 27124
rect 10284 27112 10290 27124
rect 10321 27115 10379 27121
rect 10321 27112 10333 27115
rect 10284 27084 10333 27112
rect 10284 27072 10290 27084
rect 10321 27081 10333 27084
rect 10367 27081 10379 27115
rect 11974 27112 11980 27124
rect 11935 27084 11980 27112
rect 10321 27075 10379 27081
rect 11974 27072 11980 27084
rect 12032 27072 12038 27124
rect 15289 27115 15347 27121
rect 15289 27081 15301 27115
rect 15335 27112 15347 27115
rect 16850 27112 16856 27124
rect 15335 27084 16856 27112
rect 15335 27081 15347 27084
rect 15289 27075 15347 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 17129 27115 17187 27121
rect 17129 27081 17141 27115
rect 17175 27112 17187 27115
rect 17175 27084 18828 27112
rect 17175 27081 17187 27084
rect 17129 27075 17187 27081
rect 5258 27004 5264 27056
rect 5316 27044 5322 27056
rect 7558 27044 7564 27056
rect 5316 27016 7564 27044
rect 5316 27004 5322 27016
rect 7558 27004 7564 27016
rect 7616 27004 7622 27056
rect 10594 27004 10600 27056
rect 10652 27044 10658 27056
rect 10652 27016 11560 27044
rect 10652 27004 10658 27016
rect 7006 26976 7012 26988
rect 4816 26948 7012 26976
rect 7006 26936 7012 26948
rect 7064 26936 7070 26988
rect 11054 26936 11060 26988
rect 11112 26976 11118 26988
rect 11532 26985 11560 27016
rect 12894 27004 12900 27056
rect 12952 27044 12958 27056
rect 12952 27016 13216 27044
rect 12952 27004 12958 27016
rect 13188 26985 13216 27016
rect 16684 27016 18736 27044
rect 11517 26979 11575 26985
rect 11112 26948 11468 26976
rect 11112 26936 11118 26948
rect 2409 26911 2467 26917
rect 2409 26877 2421 26911
rect 2455 26908 2467 26911
rect 2498 26908 2504 26920
rect 2455 26880 2504 26908
rect 2455 26877 2467 26880
rect 2409 26871 2467 26877
rect 2498 26868 2504 26880
rect 2556 26868 2562 26920
rect 3326 26908 3332 26920
rect 2976 26880 3332 26908
rect 1946 26800 1952 26852
rect 2004 26840 2010 26852
rect 2976 26840 3004 26880
rect 3326 26868 3332 26880
rect 3384 26908 3390 26920
rect 3789 26911 3847 26917
rect 3789 26908 3801 26911
rect 3384 26880 3801 26908
rect 3384 26868 3390 26880
rect 3789 26877 3801 26880
rect 3835 26877 3847 26911
rect 3789 26871 3847 26877
rect 3878 26868 3884 26920
rect 3936 26908 3942 26920
rect 3973 26911 4031 26917
rect 3973 26908 3985 26911
rect 3936 26880 3985 26908
rect 3936 26868 3942 26880
rect 3973 26877 3985 26880
rect 4019 26877 4031 26911
rect 3973 26871 4031 26877
rect 4065 26911 4123 26917
rect 4065 26877 4077 26911
rect 4111 26877 4123 26911
rect 4065 26871 4123 26877
rect 4080 26840 4108 26871
rect 4154 26868 4160 26920
rect 4212 26908 4218 26920
rect 4212 26880 4257 26908
rect 4212 26868 4218 26880
rect 4338 26868 4344 26920
rect 4396 26908 4402 26920
rect 4396 26880 4476 26908
rect 4396 26868 4402 26880
rect 2004 26812 3004 26840
rect 3712 26812 4108 26840
rect 4448 26840 4476 26880
rect 4798 26868 4804 26920
rect 4856 26908 4862 26920
rect 5166 26908 5172 26920
rect 4856 26880 5172 26908
rect 4856 26868 4862 26880
rect 5166 26868 5172 26880
rect 5224 26868 5230 26920
rect 8202 26868 8208 26920
rect 8260 26908 8266 26920
rect 8297 26911 8355 26917
rect 8297 26908 8309 26911
rect 8260 26880 8309 26908
rect 8260 26868 8266 26880
rect 8297 26877 8309 26880
rect 8343 26877 8355 26911
rect 8297 26871 8355 26877
rect 8941 26911 8999 26917
rect 8941 26877 8953 26911
rect 8987 26908 8999 26911
rect 9030 26908 9036 26920
rect 8987 26880 9036 26908
rect 8987 26877 8999 26880
rect 8941 26871 8999 26877
rect 9030 26868 9036 26880
rect 9088 26868 9094 26920
rect 11146 26908 11152 26920
rect 9140 26880 11152 26908
rect 4982 26840 4988 26852
rect 4448 26812 4988 26840
rect 2004 26800 2010 26812
rect 3712 26784 3740 26812
rect 4982 26800 4988 26812
rect 5040 26800 5046 26852
rect 7561 26843 7619 26849
rect 7561 26809 7573 26843
rect 7607 26840 7619 26843
rect 9140 26840 9168 26880
rect 11146 26868 11152 26880
rect 11204 26868 11210 26920
rect 11238 26868 11244 26920
rect 11296 26908 11302 26920
rect 11440 26917 11468 26948
rect 11517 26945 11529 26979
rect 11563 26945 11575 26979
rect 11517 26939 11575 26945
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26976 13231 26979
rect 14918 26976 14924 26988
rect 13219 26948 14924 26976
rect 13219 26945 13231 26948
rect 13173 26939 13231 26945
rect 14918 26936 14924 26948
rect 14976 26936 14982 26988
rect 16684 26976 16712 27016
rect 17589 26979 17647 26985
rect 16592 26948 16712 26976
rect 16868 26948 17448 26976
rect 11425 26911 11483 26917
rect 11296 26880 11341 26908
rect 11296 26868 11302 26880
rect 11425 26877 11437 26911
rect 11471 26877 11483 26911
rect 11425 26871 11483 26877
rect 11609 26911 11667 26917
rect 11609 26877 11621 26911
rect 11655 26877 11667 26911
rect 11790 26908 11796 26920
rect 11751 26880 11796 26908
rect 11609 26871 11667 26877
rect 9214 26849 9220 26852
rect 7607 26812 9168 26840
rect 7607 26809 7619 26812
rect 7561 26803 7619 26809
rect 9208 26803 9220 26849
rect 9272 26840 9278 26852
rect 9272 26812 9308 26840
rect 9214 26800 9220 26803
rect 9272 26800 9278 26812
rect 11054 26800 11060 26852
rect 11112 26840 11118 26852
rect 11624 26840 11652 26871
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 11974 26868 11980 26920
rect 12032 26908 12038 26920
rect 12805 26911 12863 26917
rect 12805 26908 12817 26911
rect 12032 26880 12817 26908
rect 12032 26868 12038 26880
rect 12805 26877 12817 26880
rect 12851 26877 12863 26911
rect 12805 26871 12863 26877
rect 12989 26911 13047 26917
rect 12989 26877 13001 26911
rect 13035 26877 13047 26911
rect 12989 26871 13047 26877
rect 13081 26911 13139 26917
rect 13081 26877 13093 26911
rect 13127 26877 13139 26911
rect 13081 26871 13139 26877
rect 11882 26840 11888 26852
rect 11112 26812 11888 26840
rect 11112 26800 11118 26812
rect 11882 26800 11888 26812
rect 11940 26800 11946 26852
rect 12342 26800 12348 26852
rect 12400 26840 12406 26852
rect 13004 26840 13032 26871
rect 12400 26812 13032 26840
rect 13096 26840 13124 26871
rect 13262 26868 13268 26920
rect 13320 26908 13326 26920
rect 13357 26911 13415 26917
rect 13357 26908 13369 26911
rect 13320 26880 13369 26908
rect 13320 26868 13326 26880
rect 13357 26877 13369 26880
rect 13403 26877 13415 26911
rect 13538 26908 13544 26920
rect 13499 26880 13544 26908
rect 13357 26871 13415 26877
rect 13538 26868 13544 26880
rect 13596 26868 13602 26920
rect 13630 26868 13636 26920
rect 13688 26908 13694 26920
rect 14274 26908 14280 26920
rect 13688 26880 14280 26908
rect 13688 26868 13694 26880
rect 14274 26868 14280 26880
rect 14332 26908 14338 26920
rect 14737 26911 14795 26917
rect 14737 26908 14749 26911
rect 14332 26880 14749 26908
rect 14332 26868 14338 26880
rect 14737 26877 14749 26880
rect 14783 26908 14795 26911
rect 16592 26908 16620 26948
rect 14783 26880 16620 26908
rect 16669 26911 16727 26917
rect 14783 26877 14795 26880
rect 14737 26871 14795 26877
rect 16669 26877 16681 26911
rect 16715 26908 16727 26911
rect 16758 26908 16764 26920
rect 16715 26880 16764 26908
rect 16715 26877 16727 26880
rect 16669 26871 16727 26877
rect 16758 26868 16764 26880
rect 16816 26868 16822 26920
rect 14458 26840 14464 26852
rect 13096 26812 14464 26840
rect 12400 26800 12406 26812
rect 14458 26800 14464 26812
rect 14516 26800 14522 26852
rect 14642 26800 14648 26852
rect 14700 26840 14706 26852
rect 15010 26840 15016 26852
rect 14700 26812 15016 26840
rect 14700 26800 14706 26812
rect 15010 26800 15016 26812
rect 15068 26840 15074 26852
rect 15068 26812 16160 26840
rect 15068 26800 15074 26812
rect 2501 26775 2559 26781
rect 2501 26741 2513 26775
rect 2547 26772 2559 26775
rect 2590 26772 2596 26784
rect 2547 26744 2596 26772
rect 2547 26741 2559 26744
rect 2501 26735 2559 26741
rect 2590 26732 2596 26744
rect 2648 26772 2654 26784
rect 2774 26772 2780 26784
rect 2648 26744 2780 26772
rect 2648 26732 2654 26744
rect 2774 26732 2780 26744
rect 2832 26732 2838 26784
rect 3234 26772 3240 26784
rect 3147 26744 3240 26772
rect 3234 26732 3240 26744
rect 3292 26772 3298 26784
rect 3694 26772 3700 26784
rect 3292 26744 3700 26772
rect 3292 26732 3298 26744
rect 3694 26732 3700 26744
rect 3752 26732 3758 26784
rect 4062 26732 4068 26784
rect 4120 26772 4126 26784
rect 4525 26775 4583 26781
rect 4525 26772 4537 26775
rect 4120 26744 4537 26772
rect 4120 26732 4126 26744
rect 4525 26741 4537 26744
rect 4571 26741 4583 26775
rect 4525 26735 4583 26741
rect 14553 26775 14611 26781
rect 14553 26741 14565 26775
rect 14599 26772 14611 26775
rect 16022 26772 16028 26784
rect 14599 26744 16028 26772
rect 14599 26741 14611 26744
rect 14553 26735 14611 26741
rect 16022 26732 16028 26744
rect 16080 26732 16086 26784
rect 16132 26772 16160 26812
rect 16298 26800 16304 26852
rect 16356 26840 16362 26852
rect 16402 26843 16460 26849
rect 16402 26840 16414 26843
rect 16356 26812 16414 26840
rect 16356 26800 16362 26812
rect 16402 26809 16414 26812
rect 16448 26809 16460 26843
rect 16402 26803 16460 26809
rect 16574 26800 16580 26852
rect 16632 26840 16638 26852
rect 16868 26840 16896 26948
rect 17420 26917 17448 26948
rect 17589 26945 17601 26979
rect 17635 26976 17647 26979
rect 17678 26976 17684 26988
rect 17635 26948 17684 26976
rect 17635 26945 17647 26948
rect 17589 26939 17647 26945
rect 17678 26936 17684 26948
rect 17736 26936 17742 26988
rect 17221 26911 17279 26917
rect 17221 26877 17233 26911
rect 17267 26877 17279 26911
rect 17221 26871 17279 26877
rect 17405 26911 17463 26917
rect 17405 26877 17417 26911
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 17497 26911 17555 26917
rect 17497 26877 17509 26911
rect 17543 26908 17555 26911
rect 17773 26911 17831 26917
rect 17543 26880 17724 26908
rect 17543 26877 17555 26880
rect 17497 26871 17555 26877
rect 16632 26812 16896 26840
rect 17236 26840 17264 26871
rect 17696 26840 17724 26880
rect 17773 26877 17785 26911
rect 17819 26908 17831 26911
rect 18138 26908 18144 26920
rect 17819 26880 18144 26908
rect 17819 26877 17831 26880
rect 17773 26871 17831 26877
rect 18138 26868 18144 26880
rect 18196 26908 18202 26920
rect 18601 26911 18659 26917
rect 18601 26908 18613 26911
rect 18196 26880 18613 26908
rect 18196 26868 18202 26880
rect 18601 26877 18613 26880
rect 18647 26877 18659 26911
rect 18708 26908 18736 27016
rect 18800 26976 18828 27084
rect 19150 27072 19156 27124
rect 19208 27112 19214 27124
rect 19613 27115 19671 27121
rect 19613 27112 19625 27115
rect 19208 27084 19625 27112
rect 19208 27072 19214 27084
rect 19613 27081 19625 27084
rect 19659 27081 19671 27115
rect 19794 27112 19800 27124
rect 19755 27084 19800 27112
rect 19613 27075 19671 27081
rect 19794 27072 19800 27084
rect 19852 27072 19858 27124
rect 20070 27072 20076 27124
rect 20128 27112 20134 27124
rect 20128 27084 20576 27112
rect 20128 27072 20134 27084
rect 19058 27004 19064 27056
rect 19116 27044 19122 27056
rect 19245 27047 19303 27053
rect 19245 27044 19257 27047
rect 19116 27016 19257 27044
rect 19116 27004 19122 27016
rect 19245 27013 19257 27016
rect 19291 27013 19303 27047
rect 19245 27007 19303 27013
rect 20162 27004 20168 27056
rect 20220 27044 20226 27056
rect 20349 27047 20407 27053
rect 20349 27044 20361 27047
rect 20220 27016 20361 27044
rect 20220 27004 20226 27016
rect 20349 27013 20361 27016
rect 20395 27013 20407 27047
rect 20548 27044 20576 27084
rect 20622 27072 20628 27124
rect 20680 27112 20686 27124
rect 20717 27115 20775 27121
rect 20717 27112 20729 27115
rect 20680 27084 20729 27112
rect 20680 27072 20686 27084
rect 20717 27081 20729 27084
rect 20763 27081 20775 27115
rect 20717 27075 20775 27081
rect 20901 27115 20959 27121
rect 20901 27081 20913 27115
rect 20947 27112 20959 27115
rect 21266 27112 21272 27124
rect 20947 27084 21272 27112
rect 20947 27081 20959 27084
rect 20901 27075 20959 27081
rect 21266 27072 21272 27084
rect 21324 27072 21330 27124
rect 24581 27115 24639 27121
rect 22949 27084 24532 27112
rect 22949 27044 22977 27084
rect 20548 27016 22977 27044
rect 20349 27007 20407 27013
rect 23014 27004 23020 27056
rect 23072 27044 23078 27056
rect 23201 27047 23259 27053
rect 23201 27044 23213 27047
rect 23072 27016 23213 27044
rect 23072 27004 23078 27016
rect 23201 27013 23213 27016
rect 23247 27013 23259 27047
rect 23201 27007 23259 27013
rect 23658 27004 23664 27056
rect 23716 27044 23722 27056
rect 24394 27044 24400 27056
rect 23716 27016 24400 27044
rect 23716 27004 23722 27016
rect 24394 27004 24400 27016
rect 24452 27004 24458 27056
rect 24504 27044 24532 27084
rect 24581 27081 24593 27115
rect 24627 27112 24639 27115
rect 24762 27112 24768 27124
rect 24627 27084 24768 27112
rect 24627 27081 24639 27084
rect 24581 27075 24639 27081
rect 24762 27072 24768 27084
rect 24820 27072 24826 27124
rect 25130 27072 25136 27124
rect 25188 27112 25194 27124
rect 25593 27115 25651 27121
rect 25593 27112 25605 27115
rect 25188 27084 25605 27112
rect 25188 27072 25194 27084
rect 25593 27081 25605 27084
rect 25639 27081 25651 27115
rect 27614 27112 27620 27124
rect 27575 27084 27620 27112
rect 25593 27075 25651 27081
rect 27614 27072 27620 27084
rect 27672 27072 27678 27124
rect 28442 27044 28448 27056
rect 24504 27016 28448 27044
rect 28442 27004 28448 27016
rect 28500 27004 28506 27056
rect 20714 26976 20720 26988
rect 18800 26948 20720 26976
rect 20714 26936 20720 26948
rect 20772 26936 20778 26988
rect 21729 26979 21787 26985
rect 21729 26945 21741 26979
rect 21775 26976 21787 26979
rect 22002 26976 22008 26988
rect 21775 26948 22008 26976
rect 21775 26945 21787 26948
rect 21729 26939 21787 26945
rect 22002 26936 22008 26948
rect 22060 26976 22066 26988
rect 25130 26976 25136 26988
rect 22060 26948 23244 26976
rect 22060 26936 22066 26948
rect 23216 26920 23244 26948
rect 24228 26948 25136 26976
rect 22554 26908 22560 26920
rect 18708 26880 22094 26908
rect 22515 26880 22560 26908
rect 18601 26871 18659 26877
rect 18230 26840 18236 26852
rect 17236 26812 17623 26840
rect 17696 26812 18236 26840
rect 16632 26800 16638 26812
rect 17129 26775 17187 26781
rect 17129 26772 17141 26775
rect 16132 26744 17141 26772
rect 17129 26741 17141 26744
rect 17175 26741 17187 26775
rect 17595 26772 17623 26812
rect 18230 26800 18236 26812
rect 18288 26800 18294 26852
rect 18340 26812 18828 26840
rect 17678 26772 17684 26784
rect 17595 26744 17684 26772
rect 17129 26735 17187 26741
rect 17678 26732 17684 26744
rect 17736 26732 17742 26784
rect 17770 26732 17776 26784
rect 17828 26772 17834 26784
rect 17957 26775 18015 26781
rect 17957 26772 17969 26775
rect 17828 26744 17969 26772
rect 17828 26732 17834 26744
rect 17957 26741 17969 26744
rect 18003 26741 18015 26775
rect 17957 26735 18015 26741
rect 18046 26732 18052 26784
rect 18104 26772 18110 26784
rect 18340 26772 18368 26812
rect 18104 26744 18368 26772
rect 18104 26732 18110 26744
rect 18414 26732 18420 26784
rect 18472 26772 18478 26784
rect 18509 26775 18567 26781
rect 18509 26772 18521 26775
rect 18472 26744 18521 26772
rect 18472 26732 18478 26744
rect 18509 26741 18521 26744
rect 18555 26741 18567 26775
rect 18800 26772 18828 26812
rect 18874 26800 18880 26852
rect 18932 26840 18938 26852
rect 19058 26840 19064 26852
rect 18932 26812 19064 26840
rect 18932 26800 18938 26812
rect 19058 26800 19064 26812
rect 19116 26800 19122 26852
rect 19518 26800 19524 26852
rect 19576 26840 19582 26852
rect 19613 26843 19671 26849
rect 19613 26840 19625 26843
rect 19576 26812 19625 26840
rect 19576 26800 19582 26812
rect 19613 26809 19625 26812
rect 19659 26809 19671 26843
rect 20714 26840 20720 26852
rect 20627 26812 20720 26840
rect 19613 26803 19671 26809
rect 20714 26800 20720 26812
rect 20772 26840 20778 26852
rect 20898 26840 20904 26852
rect 20772 26812 20904 26840
rect 20772 26800 20778 26812
rect 20898 26800 20904 26812
rect 20956 26800 20962 26852
rect 21450 26840 21456 26852
rect 21411 26812 21456 26840
rect 21450 26800 21456 26812
rect 21508 26800 21514 26852
rect 22066 26840 22094 26880
rect 22554 26868 22560 26880
rect 22612 26868 22618 26920
rect 22738 26908 22744 26920
rect 22699 26880 22744 26908
rect 22738 26868 22744 26880
rect 22796 26868 22802 26920
rect 23198 26908 23204 26920
rect 23159 26880 23204 26908
rect 23198 26868 23204 26880
rect 23256 26868 23262 26920
rect 24228 26908 24256 26948
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 29730 26976 29736 26988
rect 28368 26948 29736 26976
rect 23308 26880 24256 26908
rect 24949 26911 25007 26917
rect 23308 26840 23336 26880
rect 24949 26877 24961 26911
rect 24995 26908 25007 26911
rect 25222 26908 25228 26920
rect 24995 26880 25228 26908
rect 24995 26877 25007 26880
rect 24949 26871 25007 26877
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 26513 26911 26571 26917
rect 26513 26877 26525 26911
rect 26559 26908 26571 26911
rect 26602 26908 26608 26920
rect 26559 26880 26608 26908
rect 26559 26877 26571 26880
rect 26513 26871 26571 26877
rect 26602 26868 26608 26880
rect 26660 26868 26666 26920
rect 26970 26908 26976 26920
rect 26931 26880 26976 26908
rect 26970 26868 26976 26880
rect 27028 26868 27034 26920
rect 27157 26911 27215 26917
rect 27157 26877 27169 26911
rect 27203 26908 27215 26911
rect 27430 26908 27436 26920
rect 27203 26880 27436 26908
rect 27203 26877 27215 26880
rect 27157 26871 27215 26877
rect 27430 26868 27436 26880
rect 27488 26868 27494 26920
rect 28368 26917 28396 26948
rect 29730 26936 29736 26948
rect 29788 26936 29794 26988
rect 31202 26976 31208 26988
rect 31163 26948 31208 26976
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 28353 26911 28411 26917
rect 28353 26877 28365 26911
rect 28399 26877 28411 26911
rect 28353 26871 28411 26877
rect 28997 26911 29055 26917
rect 28997 26877 29009 26911
rect 29043 26908 29055 26911
rect 29086 26908 29092 26920
rect 29043 26880 29092 26908
rect 29043 26877 29055 26880
rect 28997 26871 29055 26877
rect 29086 26868 29092 26880
rect 29144 26868 29150 26920
rect 30926 26868 30932 26920
rect 30984 26917 30990 26920
rect 30984 26908 30996 26917
rect 30984 26880 31029 26908
rect 30984 26871 30996 26880
rect 30984 26868 30990 26871
rect 22066 26812 23336 26840
rect 23750 26800 23756 26852
rect 23808 26840 23814 26852
rect 25501 26843 25559 26849
rect 25501 26840 25513 26843
rect 23808 26812 25513 26840
rect 23808 26800 23814 26812
rect 25501 26809 25513 26812
rect 25547 26809 25559 26843
rect 25501 26803 25559 26809
rect 25682 26800 25688 26852
rect 25740 26840 25746 26852
rect 27065 26843 27123 26849
rect 27065 26840 27077 26843
rect 25740 26812 27077 26840
rect 25740 26800 25746 26812
rect 27065 26809 27077 26812
rect 27111 26809 27123 26843
rect 27065 26803 27123 26809
rect 27522 26800 27528 26852
rect 27580 26840 27586 26852
rect 31018 26840 31024 26852
rect 27580 26812 31024 26840
rect 27580 26800 27586 26812
rect 31018 26800 31024 26812
rect 31076 26800 31082 26852
rect 21082 26772 21088 26784
rect 18800 26744 21088 26772
rect 18509 26735 18567 26741
rect 21082 26732 21088 26744
rect 21140 26732 21146 26784
rect 24394 26772 24400 26784
rect 24355 26744 24400 26772
rect 24394 26732 24400 26744
rect 24452 26732 24458 26784
rect 24486 26732 24492 26784
rect 24544 26772 24550 26784
rect 24581 26775 24639 26781
rect 24581 26772 24593 26775
rect 24544 26744 24593 26772
rect 24544 26732 24550 26744
rect 24581 26741 24593 26744
rect 24627 26741 24639 26775
rect 24581 26735 24639 26741
rect 26326 26732 26332 26784
rect 26384 26772 26390 26784
rect 26421 26775 26479 26781
rect 26421 26772 26433 26775
rect 26384 26744 26433 26772
rect 26384 26732 26390 26744
rect 26421 26741 26433 26744
rect 26467 26741 26479 26775
rect 26421 26735 26479 26741
rect 27890 26732 27896 26784
rect 27948 26772 27954 26784
rect 28261 26775 28319 26781
rect 28261 26772 28273 26775
rect 27948 26744 28273 26772
rect 27948 26732 27954 26744
rect 28261 26741 28273 26744
rect 28307 26741 28319 26775
rect 28902 26772 28908 26784
rect 28863 26744 28908 26772
rect 28261 26735 28319 26741
rect 28902 26732 28908 26744
rect 28960 26732 28966 26784
rect 29825 26775 29883 26781
rect 29825 26741 29837 26775
rect 29871 26772 29883 26775
rect 30466 26772 30472 26784
rect 29871 26744 30472 26772
rect 29871 26741 29883 26744
rect 29825 26735 29883 26741
rect 30466 26732 30472 26744
rect 30524 26732 30530 26784
rect 1104 26682 32016 26704
rect 1104 26630 11253 26682
rect 11305 26630 11317 26682
rect 11369 26630 11381 26682
rect 11433 26630 11445 26682
rect 11497 26630 11509 26682
rect 11561 26630 21557 26682
rect 21609 26630 21621 26682
rect 21673 26630 21685 26682
rect 21737 26630 21749 26682
rect 21801 26630 21813 26682
rect 21865 26630 32016 26682
rect 1104 26608 32016 26630
rect 2038 26528 2044 26580
rect 2096 26528 2102 26580
rect 3421 26571 3479 26577
rect 3421 26537 3433 26571
rect 3467 26568 3479 26571
rect 3878 26568 3884 26580
rect 3467 26540 3884 26568
rect 3467 26537 3479 26540
rect 3421 26531 3479 26537
rect 3878 26528 3884 26540
rect 3936 26528 3942 26580
rect 5534 26528 5540 26580
rect 5592 26568 5598 26580
rect 5721 26571 5779 26577
rect 5721 26568 5733 26571
rect 5592 26540 5733 26568
rect 5592 26528 5598 26540
rect 5721 26537 5733 26540
rect 5767 26568 5779 26571
rect 6822 26568 6828 26580
rect 5767 26540 6828 26568
rect 5767 26537 5779 26540
rect 5721 26531 5779 26537
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 7834 26528 7840 26580
rect 7892 26568 7898 26580
rect 8754 26568 8760 26580
rect 7892 26540 8760 26568
rect 7892 26528 7898 26540
rect 8754 26528 8760 26540
rect 8812 26528 8818 26580
rect 10965 26571 11023 26577
rect 10965 26537 10977 26571
rect 11011 26568 11023 26571
rect 15654 26568 15660 26580
rect 11011 26540 15660 26568
rect 11011 26537 11023 26540
rect 10965 26531 11023 26537
rect 15654 26528 15660 26540
rect 15712 26528 15718 26580
rect 15841 26571 15899 26577
rect 15841 26537 15853 26571
rect 15887 26568 15899 26571
rect 17126 26568 17132 26580
rect 15887 26540 17132 26568
rect 15887 26537 15899 26540
rect 15841 26531 15899 26537
rect 17126 26528 17132 26540
rect 17184 26528 17190 26580
rect 17402 26528 17408 26580
rect 17460 26568 17466 26580
rect 17678 26568 17684 26580
rect 17460 26540 17684 26568
rect 17460 26528 17466 26540
rect 17678 26528 17684 26540
rect 17736 26528 17742 26580
rect 18693 26571 18751 26577
rect 18693 26537 18705 26571
rect 18739 26568 18751 26571
rect 20806 26568 20812 26580
rect 18739 26540 20812 26568
rect 18739 26537 18751 26540
rect 18693 26531 18751 26537
rect 20806 26528 20812 26540
rect 20864 26528 20870 26580
rect 22554 26528 22560 26580
rect 22612 26568 22618 26580
rect 22925 26571 22983 26577
rect 22925 26568 22937 26571
rect 22612 26540 22937 26568
rect 22612 26528 22618 26540
rect 22925 26537 22937 26540
rect 22971 26537 22983 26571
rect 22925 26531 22983 26537
rect 28718 26528 28724 26580
rect 28776 26568 28782 26580
rect 28905 26571 28963 26577
rect 28905 26568 28917 26571
rect 28776 26540 28917 26568
rect 28776 26528 28782 26540
rect 28905 26537 28917 26540
rect 28951 26537 28963 26571
rect 28905 26531 28963 26537
rect 2056 26500 2084 26528
rect 4154 26500 4160 26512
rect 2056 26472 2268 26500
rect 1946 26392 1952 26444
rect 2004 26432 2010 26444
rect 2240 26441 2268 26472
rect 2424 26472 4160 26500
rect 2424 26441 2452 26472
rect 4154 26460 4160 26472
rect 4212 26460 4218 26512
rect 4522 26460 4528 26512
rect 4580 26509 4586 26512
rect 4580 26500 4592 26509
rect 4580 26472 4625 26500
rect 4580 26463 4592 26472
rect 4580 26460 4586 26463
rect 7190 26460 7196 26512
rect 7248 26500 7254 26512
rect 11790 26500 11796 26512
rect 7248 26472 8984 26500
rect 11703 26472 11796 26500
rect 7248 26460 7254 26472
rect 2041 26435 2099 26441
rect 2041 26432 2053 26435
rect 2004 26404 2053 26432
rect 2004 26392 2010 26404
rect 2041 26401 2053 26404
rect 2087 26401 2099 26435
rect 2041 26395 2099 26401
rect 2225 26435 2283 26441
rect 2225 26401 2237 26435
rect 2271 26401 2283 26435
rect 2225 26395 2283 26401
rect 2409 26435 2467 26441
rect 2409 26401 2421 26435
rect 2455 26401 2467 26435
rect 2590 26432 2596 26444
rect 2551 26404 2596 26432
rect 2409 26395 2467 26401
rect 2590 26392 2596 26404
rect 2648 26392 2654 26444
rect 5813 26435 5871 26441
rect 5813 26401 5825 26435
rect 5859 26432 5871 26435
rect 5902 26432 5908 26444
rect 5859 26404 5908 26432
rect 5859 26401 5871 26404
rect 5813 26395 5871 26401
rect 5902 26392 5908 26404
rect 5960 26392 5966 26444
rect 6730 26432 6736 26444
rect 6691 26404 6736 26432
rect 6730 26392 6736 26404
rect 6788 26392 6794 26444
rect 6822 26392 6828 26444
rect 6880 26432 6886 26444
rect 6989 26435 7047 26441
rect 6989 26432 7001 26435
rect 6880 26404 7001 26432
rect 6880 26392 6886 26404
rect 6989 26401 7001 26404
rect 7035 26401 7047 26435
rect 6989 26395 7047 26401
rect 7742 26392 7748 26444
rect 7800 26432 7806 26444
rect 8573 26435 8631 26441
rect 8573 26432 8585 26435
rect 7800 26404 8585 26432
rect 7800 26392 7806 26404
rect 8573 26401 8585 26404
rect 8619 26401 8631 26435
rect 8754 26432 8760 26444
rect 8715 26404 8760 26432
rect 8573 26395 8631 26401
rect 8754 26392 8760 26404
rect 8812 26392 8818 26444
rect 8956 26441 8984 26472
rect 8941 26435 8999 26441
rect 8941 26401 8953 26435
rect 8987 26401 8999 26435
rect 8941 26395 8999 26401
rect 9125 26435 9183 26441
rect 9125 26401 9137 26435
rect 9171 26432 9183 26435
rect 9490 26432 9496 26444
rect 9171 26404 9496 26432
rect 9171 26401 9183 26404
rect 9125 26395 9183 26401
rect 9490 26392 9496 26404
rect 9548 26392 9554 26444
rect 11146 26392 11152 26444
rect 11204 26432 11210 26444
rect 11514 26432 11520 26444
rect 11204 26404 11520 26432
rect 11204 26392 11210 26404
rect 11514 26392 11520 26404
rect 11572 26392 11578 26444
rect 11716 26441 11744 26472
rect 11790 26460 11796 26472
rect 11848 26500 11854 26512
rect 11848 26472 12434 26500
rect 11848 26460 11854 26472
rect 11701 26435 11759 26441
rect 11701 26401 11713 26435
rect 11747 26401 11759 26435
rect 11882 26432 11888 26444
rect 11843 26404 11888 26432
rect 11701 26395 11759 26401
rect 11882 26392 11888 26404
rect 11940 26392 11946 26444
rect 11974 26392 11980 26444
rect 12032 26432 12038 26444
rect 12069 26435 12127 26441
rect 12069 26432 12081 26435
rect 12032 26404 12081 26432
rect 12032 26392 12038 26404
rect 12069 26401 12081 26404
rect 12115 26401 12127 26435
rect 12406 26432 12434 26472
rect 12526 26460 12532 26512
rect 12584 26500 12590 26512
rect 16117 26503 16175 26509
rect 12584 26472 12940 26500
rect 12584 26460 12590 26472
rect 12912 26444 12940 26472
rect 16117 26469 16129 26503
rect 16163 26500 16175 26503
rect 16206 26500 16212 26512
rect 16163 26472 16212 26500
rect 16163 26469 16175 26472
rect 16117 26463 16175 26469
rect 16206 26460 16212 26472
rect 16264 26460 16270 26512
rect 16574 26460 16580 26512
rect 16632 26500 16638 26512
rect 19613 26503 19671 26509
rect 16632 26472 19288 26500
rect 16632 26460 16638 26472
rect 12710 26432 12716 26444
rect 12406 26404 12716 26432
rect 12069 26395 12127 26401
rect 12710 26392 12716 26404
rect 12768 26392 12774 26444
rect 12894 26392 12900 26444
rect 12952 26392 12958 26444
rect 13538 26432 13544 26444
rect 13499 26404 13544 26432
rect 13538 26392 13544 26404
rect 13596 26392 13602 26444
rect 13630 26392 13636 26444
rect 13688 26432 13694 26444
rect 13725 26435 13783 26441
rect 13725 26432 13737 26435
rect 13688 26404 13737 26432
rect 13688 26392 13694 26404
rect 13725 26401 13737 26404
rect 13771 26401 13783 26435
rect 13725 26395 13783 26401
rect 14277 26435 14335 26441
rect 14277 26401 14289 26435
rect 14323 26432 14335 26435
rect 15013 26435 15071 26441
rect 15013 26432 15025 26435
rect 14323 26404 15025 26432
rect 14323 26401 14335 26404
rect 14277 26395 14335 26401
rect 15013 26401 15025 26404
rect 15059 26432 15071 26435
rect 15562 26432 15568 26444
rect 15059 26404 15568 26432
rect 15059 26401 15071 26404
rect 15013 26395 15071 26401
rect 15562 26392 15568 26404
rect 15620 26392 15626 26444
rect 15838 26432 15844 26444
rect 15799 26404 15844 26432
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 16850 26392 16856 26444
rect 16908 26432 16914 26444
rect 16908 26404 17080 26432
rect 16908 26392 16914 26404
rect 1581 26367 1639 26373
rect 1581 26333 1593 26367
rect 1627 26364 1639 26367
rect 2317 26367 2375 26373
rect 2317 26364 2329 26367
rect 1627 26336 2329 26364
rect 1627 26333 1639 26336
rect 1581 26327 1639 26333
rect 2317 26333 2329 26336
rect 2363 26364 2375 26367
rect 3234 26364 3240 26376
rect 2363 26336 3240 26364
rect 2363 26333 2375 26336
rect 2317 26327 2375 26333
rect 3234 26324 3240 26336
rect 3292 26324 3298 26376
rect 4798 26324 4804 26376
rect 4856 26364 4862 26376
rect 6748 26364 6776 26392
rect 4856 26336 6776 26364
rect 4856 26324 4862 26336
rect 8202 26324 8208 26376
rect 8260 26364 8266 26376
rect 8849 26367 8907 26373
rect 8849 26364 8861 26367
rect 8260 26336 8861 26364
rect 8260 26324 8266 26336
rect 8849 26333 8861 26336
rect 8895 26333 8907 26367
rect 8849 26327 8907 26333
rect 10594 26324 10600 26376
rect 10652 26364 10658 26376
rect 11793 26367 11851 26373
rect 11793 26364 11805 26367
rect 10652 26336 11805 26364
rect 10652 26324 10658 26336
rect 11793 26333 11805 26336
rect 11839 26333 11851 26367
rect 11793 26327 11851 26333
rect 12342 26324 12348 26376
rect 12400 26364 12406 26376
rect 12728 26364 12756 26392
rect 13262 26364 13268 26376
rect 12400 26336 12664 26364
rect 12728 26336 13268 26364
rect 12400 26324 12406 26336
rect 2498 26256 2504 26308
rect 2556 26296 2562 26308
rect 2777 26299 2835 26305
rect 2777 26296 2789 26299
rect 2556 26268 2789 26296
rect 2556 26256 2562 26268
rect 2777 26265 2789 26268
rect 2823 26265 2835 26299
rect 2777 26259 2835 26265
rect 8294 26256 8300 26308
rect 8352 26296 8358 26308
rect 9769 26299 9827 26305
rect 9769 26296 9781 26299
rect 8352 26268 9781 26296
rect 8352 26256 8358 26268
rect 9769 26265 9781 26268
rect 9815 26265 9827 26299
rect 9769 26259 9827 26265
rect 10413 26299 10471 26305
rect 10413 26265 10425 26299
rect 10459 26296 10471 26299
rect 12253 26299 12311 26305
rect 10459 26268 12204 26296
rect 10459 26265 10471 26268
rect 10413 26259 10471 26265
rect 1854 26188 1860 26240
rect 1912 26228 1918 26240
rect 2314 26228 2320 26240
rect 1912 26200 2320 26228
rect 1912 26188 1918 26200
rect 2314 26188 2320 26200
rect 2372 26188 2378 26240
rect 5902 26188 5908 26240
rect 5960 26228 5966 26240
rect 6454 26228 6460 26240
rect 5960 26200 6460 26228
rect 5960 26188 5966 26200
rect 6454 26188 6460 26200
rect 6512 26228 6518 26240
rect 7006 26228 7012 26240
rect 6512 26200 7012 26228
rect 6512 26188 6518 26200
rect 7006 26188 7012 26200
rect 7064 26228 7070 26240
rect 8113 26231 8171 26237
rect 8113 26228 8125 26231
rect 7064 26200 8125 26228
rect 7064 26188 7070 26200
rect 8113 26197 8125 26200
rect 8159 26197 8171 26231
rect 9306 26228 9312 26240
rect 9267 26200 9312 26228
rect 8113 26191 8171 26197
rect 9306 26188 9312 26200
rect 9364 26188 9370 26240
rect 11514 26188 11520 26240
rect 11572 26228 11578 26240
rect 12066 26228 12072 26240
rect 11572 26200 12072 26228
rect 11572 26188 11578 26200
rect 12066 26188 12072 26200
rect 12124 26188 12130 26240
rect 12176 26228 12204 26268
rect 12253 26265 12265 26299
rect 12299 26296 12311 26299
rect 12434 26296 12440 26308
rect 12299 26268 12440 26296
rect 12299 26265 12311 26268
rect 12253 26259 12311 26265
rect 12434 26256 12440 26268
rect 12492 26256 12498 26308
rect 12526 26256 12532 26308
rect 12584 26256 12590 26308
rect 12636 26296 12664 26336
rect 13262 26324 13268 26336
rect 13320 26324 13326 26376
rect 14458 26324 14464 26376
rect 14516 26364 14522 26376
rect 16298 26364 16304 26376
rect 14516 26336 16304 26364
rect 14516 26324 14522 26336
rect 16298 26324 16304 26336
rect 16356 26324 16362 26376
rect 16942 26364 16948 26376
rect 16903 26336 16948 26364
rect 16942 26324 16948 26336
rect 17000 26324 17006 26376
rect 17052 26364 17080 26404
rect 17126 26392 17132 26444
rect 17184 26432 17190 26444
rect 17589 26435 17647 26441
rect 17589 26432 17601 26435
rect 17184 26404 17229 26432
rect 17328 26404 17601 26432
rect 17184 26392 17190 26404
rect 17328 26364 17356 26404
rect 17589 26401 17601 26404
rect 17635 26401 17647 26435
rect 17862 26432 17868 26444
rect 17823 26404 17868 26432
rect 17589 26395 17647 26401
rect 17862 26392 17868 26404
rect 17920 26392 17926 26444
rect 17954 26392 17960 26444
rect 18012 26432 18018 26444
rect 19260 26441 19288 26472
rect 19613 26469 19625 26503
rect 19659 26500 19671 26503
rect 20714 26500 20720 26512
rect 19659 26472 20720 26500
rect 19659 26469 19671 26472
rect 19613 26463 19671 26469
rect 20714 26460 20720 26472
rect 20772 26460 20778 26512
rect 22646 26460 22652 26512
rect 22704 26500 22710 26512
rect 22704 26472 22784 26500
rect 22704 26460 22710 26472
rect 18509 26435 18567 26441
rect 18509 26432 18521 26435
rect 18012 26404 18521 26432
rect 18012 26392 18018 26404
rect 18509 26401 18521 26404
rect 18555 26401 18567 26435
rect 18509 26395 18567 26401
rect 19245 26435 19303 26441
rect 19245 26401 19257 26435
rect 19291 26432 19303 26435
rect 19702 26432 19708 26444
rect 19291 26404 19708 26432
rect 19291 26401 19303 26404
rect 19245 26395 19303 26401
rect 19702 26392 19708 26404
rect 19760 26432 19766 26444
rect 20257 26435 20315 26441
rect 20257 26432 20269 26435
rect 19760 26404 20269 26432
rect 19760 26392 19766 26404
rect 20257 26401 20269 26404
rect 20303 26401 20315 26435
rect 20438 26432 20444 26444
rect 20399 26404 20444 26432
rect 20257 26395 20315 26401
rect 20438 26392 20444 26404
rect 20496 26392 20502 26444
rect 20530 26392 20536 26444
rect 20588 26432 20594 26444
rect 20809 26435 20867 26441
rect 20588 26404 20633 26432
rect 20588 26392 20594 26404
rect 20809 26401 20821 26435
rect 20855 26432 20867 26435
rect 22189 26435 22247 26441
rect 20855 26404 20944 26432
rect 20855 26401 20867 26404
rect 20809 26395 20867 26401
rect 18414 26364 18420 26376
rect 17052 26336 17356 26364
rect 17420 26336 18420 26364
rect 12805 26299 12863 26305
rect 12805 26296 12817 26299
rect 12636 26268 12817 26296
rect 12805 26265 12817 26268
rect 12851 26265 12863 26299
rect 12805 26259 12863 26265
rect 13078 26256 13084 26308
rect 13136 26296 13142 26308
rect 14185 26299 14243 26305
rect 14185 26296 14197 26299
rect 13136 26268 14197 26296
rect 13136 26256 13142 26268
rect 14185 26265 14197 26268
rect 14231 26265 14243 26299
rect 14185 26259 14243 26265
rect 15933 26299 15991 26305
rect 15933 26265 15945 26299
rect 15979 26296 15991 26299
rect 17420 26296 17448 26336
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 19978 26364 19984 26376
rect 19306 26336 19984 26364
rect 19306 26308 19334 26336
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 20162 26324 20168 26376
rect 20220 26364 20226 26376
rect 20625 26367 20683 26373
rect 20625 26364 20637 26367
rect 20220 26336 20637 26364
rect 20220 26324 20226 26336
rect 20625 26333 20637 26336
rect 20671 26333 20683 26367
rect 20625 26327 20683 26333
rect 19306 26296 19340 26308
rect 15979 26268 17448 26296
rect 17926 26268 19340 26296
rect 15979 26265 15991 26268
rect 15933 26259 15991 26265
rect 12544 26228 12572 26256
rect 12176 26200 12572 26228
rect 13814 26188 13820 26240
rect 13872 26228 13878 26240
rect 15105 26231 15163 26237
rect 15105 26228 15117 26231
rect 13872 26200 15117 26228
rect 13872 26188 13878 26200
rect 15105 26197 15117 26200
rect 15151 26228 15163 26231
rect 15378 26228 15384 26240
rect 15151 26200 15384 26228
rect 15151 26197 15163 26200
rect 15105 26191 15163 26197
rect 15378 26188 15384 26200
rect 15436 26228 15442 26240
rect 16206 26228 16212 26240
rect 15436 26200 16212 26228
rect 15436 26188 15442 26200
rect 16206 26188 16212 26200
rect 16264 26188 16270 26240
rect 16298 26188 16304 26240
rect 16356 26228 16362 26240
rect 17926 26228 17954 26268
rect 19334 26256 19340 26268
rect 19392 26256 19398 26308
rect 19797 26299 19855 26305
rect 19797 26265 19809 26299
rect 19843 26296 19855 26299
rect 20714 26296 20720 26308
rect 19843 26268 20720 26296
rect 19843 26265 19855 26268
rect 19797 26259 19855 26265
rect 20714 26256 20720 26268
rect 20772 26256 20778 26308
rect 20916 26296 20944 26404
rect 22189 26401 22201 26435
rect 22235 26432 22247 26435
rect 22278 26432 22284 26444
rect 22235 26404 22284 26432
rect 22235 26401 22247 26404
rect 22189 26395 22247 26401
rect 22278 26392 22284 26404
rect 22336 26392 22342 26444
rect 22756 26441 22784 26472
rect 23198 26460 23204 26512
rect 23256 26500 23262 26512
rect 23753 26503 23811 26509
rect 23256 26472 23336 26500
rect 23256 26460 23262 26472
rect 22373 26435 22431 26441
rect 22373 26401 22385 26435
rect 22419 26432 22431 26435
rect 22741 26435 22799 26441
rect 22419 26404 22701 26432
rect 22419 26401 22431 26404
rect 22373 26395 22431 26401
rect 22465 26367 22523 26373
rect 22465 26364 22477 26367
rect 22204 26336 22477 26364
rect 20835 26268 20944 26296
rect 20835 26240 20863 26268
rect 22002 26256 22008 26308
rect 22060 26296 22066 26308
rect 22204 26296 22232 26336
rect 22465 26333 22477 26336
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 22557 26367 22615 26373
rect 22557 26333 22569 26367
rect 22603 26333 22615 26367
rect 22673 26364 22701 26404
rect 22741 26401 22753 26435
rect 22787 26432 22799 26435
rect 23106 26432 23112 26444
rect 22787 26404 23112 26432
rect 22787 26401 22799 26404
rect 22741 26395 22799 26401
rect 23106 26392 23112 26404
rect 23164 26392 23170 26444
rect 23198 26364 23204 26376
rect 22673 26336 23204 26364
rect 22557 26327 22615 26333
rect 22060 26268 22232 26296
rect 22060 26256 22066 26268
rect 16356 26200 17954 26228
rect 19613 26231 19671 26237
rect 16356 26188 16362 26200
rect 19613 26197 19625 26231
rect 19659 26228 19671 26231
rect 20806 26228 20812 26240
rect 19659 26200 20812 26228
rect 19659 26197 19671 26200
rect 19613 26191 19671 26197
rect 20806 26188 20812 26200
rect 20864 26188 20870 26240
rect 20990 26228 20996 26240
rect 20951 26200 20996 26228
rect 20990 26188 20996 26200
rect 21048 26188 21054 26240
rect 21082 26188 21088 26240
rect 21140 26228 21146 26240
rect 22572 26228 22600 26327
rect 23198 26324 23204 26336
rect 23256 26324 23262 26376
rect 22646 26256 22652 26308
rect 22704 26296 22710 26308
rect 23308 26296 23336 26472
rect 23753 26469 23765 26503
rect 23799 26500 23811 26503
rect 24026 26500 24032 26512
rect 23799 26472 24032 26500
rect 23799 26469 23811 26472
rect 23753 26463 23811 26469
rect 24026 26460 24032 26472
rect 24084 26460 24090 26512
rect 24394 26460 24400 26512
rect 24452 26500 24458 26512
rect 24452 26472 24900 26500
rect 24452 26460 24458 26472
rect 23385 26435 23443 26441
rect 23385 26401 23397 26435
rect 23431 26401 23443 26435
rect 23566 26432 23572 26444
rect 23527 26404 23572 26432
rect 23385 26395 23443 26401
rect 23400 26364 23428 26395
rect 23566 26392 23572 26404
rect 23624 26392 23630 26444
rect 23842 26392 23848 26444
rect 23900 26432 23906 26444
rect 24581 26435 24639 26441
rect 24581 26432 24593 26435
rect 23900 26404 24593 26432
rect 23900 26392 23906 26404
rect 24581 26401 24593 26404
rect 24627 26432 24639 26435
rect 24670 26432 24676 26444
rect 24627 26404 24676 26432
rect 24627 26401 24639 26404
rect 24581 26395 24639 26401
rect 24670 26392 24676 26404
rect 24728 26392 24734 26444
rect 24872 26441 24900 26472
rect 26234 26460 26240 26512
rect 26292 26500 26298 26512
rect 28445 26503 28503 26509
rect 28445 26500 28457 26503
rect 26292 26472 28457 26500
rect 26292 26460 26298 26472
rect 28445 26469 28457 26472
rect 28491 26469 28503 26503
rect 28445 26463 28503 26469
rect 24857 26435 24915 26441
rect 24857 26401 24869 26435
rect 24903 26401 24915 26435
rect 24857 26395 24915 26401
rect 25130 26392 25136 26444
rect 25188 26432 25194 26444
rect 25869 26435 25927 26441
rect 25869 26432 25881 26435
rect 25188 26404 25881 26432
rect 25188 26392 25194 26404
rect 25869 26401 25881 26404
rect 25915 26401 25927 26435
rect 25869 26395 25927 26401
rect 26142 26392 26148 26444
rect 26200 26432 26206 26444
rect 26973 26435 27031 26441
rect 26973 26432 26985 26435
rect 26200 26404 26985 26432
rect 26200 26392 26206 26404
rect 26973 26401 26985 26404
rect 27019 26401 27031 26435
rect 27706 26432 27712 26444
rect 27667 26404 27712 26432
rect 26973 26395 27031 26401
rect 27706 26392 27712 26404
rect 27764 26392 27770 26444
rect 27890 26432 27896 26444
rect 27851 26404 27896 26432
rect 27890 26392 27896 26404
rect 27948 26392 27954 26444
rect 28261 26435 28319 26441
rect 28261 26401 28273 26435
rect 28307 26432 28319 26435
rect 28902 26432 28908 26444
rect 28307 26404 28908 26432
rect 28307 26401 28319 26404
rect 28261 26395 28319 26401
rect 28902 26392 28908 26404
rect 28960 26392 28966 26444
rect 29270 26392 29276 26444
rect 29328 26432 29334 26444
rect 29457 26435 29515 26441
rect 29457 26432 29469 26435
rect 29328 26404 29469 26432
rect 29328 26392 29334 26404
rect 29457 26401 29469 26404
rect 29503 26432 29515 26435
rect 29546 26432 29552 26444
rect 29503 26404 29552 26432
rect 29503 26401 29515 26404
rect 29457 26395 29515 26401
rect 29546 26392 29552 26404
rect 29604 26392 29610 26444
rect 29641 26435 29699 26441
rect 29641 26401 29653 26435
rect 29687 26432 29699 26435
rect 29687 26404 29969 26432
rect 29687 26401 29699 26404
rect 29641 26395 29699 26401
rect 24026 26364 24032 26376
rect 23400 26336 24032 26364
rect 24026 26324 24032 26336
rect 24084 26324 24090 26376
rect 24946 26324 24952 26376
rect 25004 26364 25010 26376
rect 25225 26367 25283 26373
rect 25225 26364 25237 26367
rect 25004 26336 25237 26364
rect 25004 26324 25010 26336
rect 25225 26333 25237 26336
rect 25271 26333 25283 26367
rect 27246 26364 27252 26376
rect 25225 26327 25283 26333
rect 25332 26336 27252 26364
rect 22704 26268 23336 26296
rect 22704 26256 22710 26268
rect 24302 26256 24308 26308
rect 24360 26296 24366 26308
rect 24578 26296 24584 26308
rect 24360 26268 24584 26296
rect 24360 26256 24366 26268
rect 24578 26256 24584 26268
rect 24636 26256 24642 26308
rect 23014 26228 23020 26240
rect 21140 26200 23020 26228
rect 21140 26188 21146 26200
rect 23014 26188 23020 26200
rect 23072 26228 23078 26240
rect 25332 26228 25360 26336
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 27522 26324 27528 26376
rect 27580 26364 27586 26376
rect 27985 26367 28043 26373
rect 27985 26364 27997 26367
rect 27580 26336 27997 26364
rect 27580 26324 27586 26336
rect 27985 26333 27997 26336
rect 28031 26333 28043 26367
rect 27985 26327 28043 26333
rect 28074 26324 28080 26376
rect 28132 26364 28138 26376
rect 29733 26367 29791 26373
rect 29733 26364 29745 26367
rect 28132 26336 28177 26364
rect 29564 26336 29745 26364
rect 28132 26324 28138 26336
rect 27065 26299 27123 26305
rect 27065 26265 27077 26299
rect 27111 26296 27123 26299
rect 27154 26296 27160 26308
rect 27111 26268 27160 26296
rect 27111 26265 27123 26268
rect 27065 26259 27123 26265
rect 27154 26256 27160 26268
rect 27212 26256 27218 26308
rect 28092 26296 28120 26324
rect 29564 26308 29592 26336
rect 29733 26333 29745 26336
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 29825 26367 29883 26373
rect 29825 26333 29837 26367
rect 29871 26333 29883 26367
rect 29941 26364 29969 26404
rect 30006 26392 30012 26444
rect 30064 26432 30070 26444
rect 30064 26404 30109 26432
rect 30064 26392 30070 26404
rect 30558 26392 30564 26444
rect 30616 26432 30622 26444
rect 30837 26435 30895 26441
rect 30837 26432 30849 26435
rect 30616 26404 30849 26432
rect 30616 26392 30622 26404
rect 30837 26401 30849 26404
rect 30883 26401 30895 26435
rect 30837 26395 30895 26401
rect 31018 26392 31024 26444
rect 31076 26392 31082 26444
rect 30466 26364 30472 26376
rect 29941 26336 30472 26364
rect 29825 26327 29883 26333
rect 27264 26268 28120 26296
rect 25866 26228 25872 26240
rect 23072 26200 25360 26228
rect 25827 26200 25872 26228
rect 23072 26188 23078 26200
rect 25866 26188 25872 26200
rect 25924 26188 25930 26240
rect 26510 26188 26516 26240
rect 26568 26228 26574 26240
rect 27264 26228 27292 26268
rect 29546 26256 29552 26308
rect 29604 26256 29610 26308
rect 29840 26296 29868 26327
rect 30466 26324 30472 26336
rect 30524 26324 30530 26376
rect 30650 26324 30656 26376
rect 30708 26364 30714 26376
rect 30745 26367 30803 26373
rect 30745 26364 30757 26367
rect 30708 26336 30757 26364
rect 30708 26324 30714 26336
rect 30745 26333 30757 26336
rect 30791 26364 30803 26367
rect 31036 26364 31064 26392
rect 30791 26336 31064 26364
rect 30791 26333 30803 26336
rect 30745 26327 30803 26333
rect 29914 26296 29920 26308
rect 29840 26268 29920 26296
rect 29914 26256 29920 26268
rect 29972 26256 29978 26308
rect 30193 26299 30251 26305
rect 30193 26265 30205 26299
rect 30239 26296 30251 26299
rect 31018 26296 31024 26308
rect 30239 26268 31024 26296
rect 30239 26265 30251 26268
rect 30193 26259 30251 26265
rect 31018 26256 31024 26268
rect 31076 26256 31082 26308
rect 26568 26200 27292 26228
rect 26568 26188 26574 26200
rect 1104 26138 32016 26160
rect 1104 26086 6102 26138
rect 6154 26086 6166 26138
rect 6218 26086 6230 26138
rect 6282 26086 6294 26138
rect 6346 26086 6358 26138
rect 6410 26086 16405 26138
rect 16457 26086 16469 26138
rect 16521 26086 16533 26138
rect 16585 26086 16597 26138
rect 16649 26086 16661 26138
rect 16713 26086 26709 26138
rect 26761 26086 26773 26138
rect 26825 26086 26837 26138
rect 26889 26086 26901 26138
rect 26953 26086 26965 26138
rect 27017 26086 32016 26138
rect 1104 26064 32016 26086
rect 1394 26024 1400 26036
rect 1355 25996 1400 26024
rect 1394 25984 1400 25996
rect 1452 25984 1458 26036
rect 5166 26024 5172 26036
rect 5127 25996 5172 26024
rect 5166 25984 5172 25996
rect 5224 25984 5230 26036
rect 6822 26024 6828 26036
rect 6783 25996 6828 26024
rect 6822 25984 6828 25996
rect 6880 25984 6886 26036
rect 8202 26024 8208 26036
rect 8163 25996 8208 26024
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 12802 25984 12808 26036
rect 12860 26024 12866 26036
rect 13078 26024 13084 26036
rect 12860 25996 13084 26024
rect 12860 25984 12866 25996
rect 13078 25984 13084 25996
rect 13136 25984 13142 26036
rect 14185 26027 14243 26033
rect 14185 25993 14197 26027
rect 14231 26024 14243 26027
rect 14274 26024 14280 26036
rect 14231 25996 14280 26024
rect 14231 25993 14243 25996
rect 14185 25987 14243 25993
rect 14274 25984 14280 25996
rect 14332 25984 14338 26036
rect 14366 25984 14372 26036
rect 14424 26024 14430 26036
rect 15013 26027 15071 26033
rect 15013 26024 15025 26027
rect 14424 25996 15025 26024
rect 14424 25984 14430 25996
rect 15013 25993 15025 25996
rect 15059 25993 15071 26027
rect 16114 26024 16120 26036
rect 16075 25996 16120 26024
rect 15013 25987 15071 25993
rect 16114 25984 16120 25996
rect 16172 25984 16178 26036
rect 16942 25984 16948 26036
rect 17000 26024 17006 26036
rect 17865 26027 17923 26033
rect 17865 26024 17877 26027
rect 17000 25996 17877 26024
rect 17000 25984 17006 25996
rect 17865 25993 17877 25996
rect 17911 25993 17923 26027
rect 19702 26024 19708 26036
rect 19663 25996 19708 26024
rect 17865 25987 17923 25993
rect 19702 25984 19708 25996
rect 19760 25984 19766 26036
rect 21450 25984 21456 26036
rect 21508 26024 21514 26036
rect 21545 26027 21603 26033
rect 21545 26024 21557 26027
rect 21508 25996 21557 26024
rect 21508 25984 21514 25996
rect 21545 25993 21557 25996
rect 21591 25993 21603 26027
rect 21545 25987 21603 25993
rect 22465 26027 22523 26033
rect 22465 25993 22477 26027
rect 22511 26024 22523 26027
rect 22554 26024 22560 26036
rect 22511 25996 22560 26024
rect 22511 25993 22523 25996
rect 22465 25987 22523 25993
rect 22554 25984 22560 25996
rect 22612 25984 22618 26036
rect 22649 26027 22707 26033
rect 22649 25993 22661 26027
rect 22695 26024 22707 26027
rect 22738 26024 22744 26036
rect 22695 25996 22744 26024
rect 22695 25993 22707 25996
rect 22649 25987 22707 25993
rect 22738 25984 22744 25996
rect 22796 25984 22802 26036
rect 27522 26024 27528 26036
rect 26896 25996 27528 26024
rect 10870 25916 10876 25968
rect 10928 25956 10934 25968
rect 11609 25959 11667 25965
rect 11609 25956 11621 25959
rect 10928 25928 11621 25956
rect 10928 25916 10934 25928
rect 11609 25925 11621 25928
rect 11655 25956 11667 25959
rect 11974 25956 11980 25968
rect 11655 25928 11980 25956
rect 11655 25925 11667 25928
rect 11609 25919 11667 25925
rect 11974 25916 11980 25928
rect 12032 25916 12038 25968
rect 14918 25916 14924 25968
rect 14976 25956 14982 25968
rect 15470 25956 15476 25968
rect 14976 25928 15476 25956
rect 14976 25916 14982 25928
rect 15470 25916 15476 25928
rect 15528 25956 15534 25968
rect 18046 25956 18052 25968
rect 15528 25928 18052 25956
rect 15528 25916 15534 25928
rect 18046 25916 18052 25928
rect 18104 25916 18110 25968
rect 18506 25956 18512 25968
rect 18248 25928 18512 25956
rect 6638 25848 6644 25900
rect 6696 25888 6702 25900
rect 7285 25891 7343 25897
rect 7285 25888 7297 25891
rect 6696 25860 7297 25888
rect 6696 25848 6702 25860
rect 7285 25857 7297 25860
rect 7331 25857 7343 25891
rect 7285 25851 7343 25857
rect 7742 25848 7748 25900
rect 7800 25848 7806 25900
rect 9030 25888 9036 25900
rect 8991 25860 9036 25888
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 18248 25897 18276 25928
rect 18506 25916 18512 25928
rect 18564 25916 18570 25968
rect 22094 25916 22100 25968
rect 22152 25956 22158 25968
rect 23201 25959 23259 25965
rect 23201 25956 23213 25959
rect 22152 25928 23213 25956
rect 22152 25916 22158 25928
rect 23201 25925 23213 25928
rect 23247 25925 23259 25959
rect 23201 25919 23259 25925
rect 26418 25916 26424 25968
rect 26476 25956 26482 25968
rect 26694 25956 26700 25968
rect 26476 25928 26700 25956
rect 26476 25916 26482 25928
rect 26694 25916 26700 25928
rect 26752 25916 26758 25968
rect 18233 25891 18291 25897
rect 18233 25888 18245 25891
rect 14568 25860 18245 25888
rect 2498 25820 2504 25832
rect 2556 25829 2562 25832
rect 2468 25792 2504 25820
rect 2498 25780 2504 25792
rect 2556 25783 2568 25829
rect 2556 25780 2562 25783
rect 2774 25780 2780 25832
rect 2832 25820 2838 25832
rect 3789 25823 3847 25829
rect 3789 25820 3801 25823
rect 2832 25792 3801 25820
rect 2832 25780 2838 25792
rect 3789 25789 3801 25792
rect 3835 25820 3847 25823
rect 4798 25820 4804 25832
rect 3835 25792 4804 25820
rect 3835 25789 3847 25792
rect 3789 25783 3847 25789
rect 4798 25780 4804 25792
rect 4856 25780 4862 25832
rect 7006 25820 7012 25832
rect 6967 25792 7012 25820
rect 7006 25780 7012 25792
rect 7064 25780 7070 25832
rect 7190 25820 7196 25832
rect 7151 25792 7196 25820
rect 7190 25780 7196 25792
rect 7248 25780 7254 25832
rect 7377 25823 7435 25829
rect 7377 25820 7389 25823
rect 7300 25792 7389 25820
rect 7300 25764 7328 25792
rect 7377 25789 7389 25792
rect 7423 25789 7435 25823
rect 7377 25783 7435 25789
rect 7561 25823 7619 25829
rect 7561 25789 7573 25823
rect 7607 25820 7619 25823
rect 7760 25820 7788 25848
rect 8018 25820 8024 25832
rect 7607 25792 7788 25820
rect 7979 25792 8024 25820
rect 7607 25789 7619 25792
rect 7561 25783 7619 25789
rect 8018 25780 8024 25792
rect 8076 25780 8082 25832
rect 9306 25829 9312 25832
rect 9300 25820 9312 25829
rect 9267 25792 9312 25820
rect 9300 25783 9312 25792
rect 9306 25780 9312 25783
rect 9364 25780 9370 25832
rect 12434 25780 12440 25832
rect 12492 25820 12498 25832
rect 12722 25823 12780 25829
rect 12722 25820 12734 25823
rect 12492 25792 12734 25820
rect 12492 25780 12498 25792
rect 12722 25789 12734 25792
rect 12768 25789 12780 25823
rect 12986 25820 12992 25832
rect 12899 25792 12992 25820
rect 12722 25783 12780 25789
rect 12986 25780 12992 25792
rect 13044 25820 13050 25832
rect 13538 25820 13544 25832
rect 13044 25792 13544 25820
rect 13044 25780 13050 25792
rect 13538 25780 13544 25792
rect 13596 25780 13602 25832
rect 4062 25761 4068 25764
rect 4056 25752 4068 25761
rect 4023 25724 4068 25752
rect 4056 25715 4068 25724
rect 4062 25712 4068 25715
rect 4120 25712 4126 25764
rect 6914 25712 6920 25764
rect 6972 25752 6978 25764
rect 7282 25752 7288 25764
rect 6972 25724 7288 25752
rect 6972 25712 6978 25724
rect 7282 25712 7288 25724
rect 7340 25712 7346 25764
rect 7742 25712 7748 25764
rect 7800 25752 7806 25764
rect 14568 25752 14596 25860
rect 18233 25857 18245 25860
rect 18279 25857 18291 25891
rect 18233 25851 18291 25857
rect 18325 25891 18383 25897
rect 18325 25857 18337 25891
rect 18371 25888 18383 25891
rect 21085 25891 21143 25897
rect 18371 25860 20116 25888
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 14642 25780 14648 25832
rect 14700 25820 14706 25832
rect 18049 25823 18107 25829
rect 14700 25792 14745 25820
rect 14700 25780 14706 25792
rect 18049 25789 18061 25823
rect 18095 25820 18107 25823
rect 18138 25820 18144 25832
rect 18095 25792 18144 25820
rect 18095 25789 18107 25792
rect 18049 25783 18107 25789
rect 18138 25780 18144 25792
rect 18196 25780 18202 25832
rect 18414 25820 18420 25832
rect 18375 25792 18420 25820
rect 18414 25780 18420 25792
rect 18472 25780 18478 25832
rect 18598 25820 18604 25832
rect 18559 25792 18604 25820
rect 18598 25780 18604 25792
rect 18656 25780 18662 25832
rect 20088 25820 20116 25860
rect 21085 25857 21097 25891
rect 21131 25888 21143 25891
rect 22186 25888 22192 25900
rect 21131 25860 22192 25888
rect 21131 25857 21143 25860
rect 21085 25851 21143 25857
rect 22186 25848 22192 25860
rect 22244 25888 22250 25900
rect 22738 25888 22744 25900
rect 22244 25860 22744 25888
rect 22244 25848 22250 25860
rect 22738 25848 22744 25860
rect 22796 25848 22802 25900
rect 25409 25891 25467 25897
rect 25409 25857 25421 25891
rect 25455 25888 25467 25891
rect 25682 25888 25688 25900
rect 25455 25860 25688 25888
rect 25455 25857 25467 25860
rect 25409 25851 25467 25857
rect 25682 25848 25688 25860
rect 25740 25848 25746 25900
rect 26510 25848 26516 25900
rect 26568 25888 26574 25900
rect 26896 25897 26924 25996
rect 27522 25984 27528 25996
rect 27580 25984 27586 26036
rect 27706 26024 27712 26036
rect 27667 25996 27712 26024
rect 27706 25984 27712 25996
rect 27764 25984 27770 26036
rect 27338 25956 27344 25968
rect 26988 25928 27344 25956
rect 26789 25891 26847 25897
rect 26789 25888 26801 25891
rect 26568 25860 26801 25888
rect 26568 25848 26574 25860
rect 26789 25857 26801 25860
rect 26835 25857 26847 25891
rect 26789 25851 26847 25857
rect 26881 25891 26939 25897
rect 26881 25857 26893 25891
rect 26927 25857 26939 25891
rect 26881 25851 26939 25857
rect 20254 25820 20260 25832
rect 20088 25792 20260 25820
rect 20254 25780 20260 25792
rect 20312 25780 20318 25832
rect 22097 25823 22155 25829
rect 22097 25789 22109 25823
rect 22143 25820 22155 25823
rect 22278 25820 22284 25832
rect 22143 25792 22284 25820
rect 22143 25789 22155 25792
rect 22097 25783 22155 25789
rect 22278 25780 22284 25792
rect 22336 25780 22342 25832
rect 23109 25823 23167 25829
rect 23109 25789 23121 25823
rect 23155 25820 23167 25823
rect 23290 25820 23296 25832
rect 23155 25792 23296 25820
rect 23155 25789 23167 25792
rect 23109 25783 23167 25789
rect 23290 25780 23296 25792
rect 23348 25780 23354 25832
rect 24581 25823 24639 25829
rect 24581 25789 24593 25823
rect 24627 25789 24639 25823
rect 24581 25783 24639 25789
rect 15010 25752 15016 25764
rect 7800 25724 14596 25752
rect 14971 25724 15016 25752
rect 7800 25712 7806 25724
rect 15010 25712 15016 25724
rect 15068 25712 15074 25764
rect 17405 25755 17463 25761
rect 15120 25724 17356 25752
rect 5534 25644 5540 25696
rect 5592 25684 5598 25696
rect 5629 25687 5687 25693
rect 5629 25684 5641 25687
rect 5592 25656 5641 25684
rect 5592 25644 5598 25656
rect 5629 25653 5641 25656
rect 5675 25653 5687 25687
rect 5629 25647 5687 25653
rect 6365 25687 6423 25693
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 6822 25684 6828 25696
rect 6411 25656 6828 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 8202 25644 8208 25696
rect 8260 25684 8266 25696
rect 8478 25684 8484 25696
rect 8260 25656 8484 25684
rect 8260 25644 8266 25656
rect 8478 25644 8484 25656
rect 8536 25644 8542 25696
rect 10410 25684 10416 25696
rect 10371 25656 10416 25684
rect 10410 25644 10416 25656
rect 10468 25644 10474 25696
rect 11054 25684 11060 25696
rect 11015 25656 11060 25684
rect 11054 25644 11060 25656
rect 11112 25644 11118 25696
rect 13262 25644 13268 25696
rect 13320 25684 13326 25696
rect 13449 25687 13507 25693
rect 13449 25684 13461 25687
rect 13320 25656 13461 25684
rect 13320 25644 13326 25656
rect 13449 25653 13461 25656
rect 13495 25653 13507 25687
rect 13449 25647 13507 25653
rect 14458 25644 14464 25696
rect 14516 25684 14522 25696
rect 15120 25684 15148 25724
rect 14516 25656 15148 25684
rect 15197 25687 15255 25693
rect 14516 25644 14522 25656
rect 15197 25653 15209 25687
rect 15243 25684 15255 25687
rect 15378 25684 15384 25696
rect 15243 25656 15384 25684
rect 15243 25653 15255 25656
rect 15197 25647 15255 25653
rect 15378 25644 15384 25656
rect 15436 25644 15442 25696
rect 17328 25684 17356 25724
rect 17405 25721 17417 25755
rect 17451 25752 17463 25755
rect 18874 25752 18880 25764
rect 17451 25724 18880 25752
rect 17451 25721 17463 25724
rect 17405 25715 17463 25721
rect 18874 25712 18880 25724
rect 18932 25712 18938 25764
rect 20070 25712 20076 25764
rect 20128 25752 20134 25764
rect 20818 25755 20876 25761
rect 20818 25752 20830 25755
rect 20128 25724 20830 25752
rect 20128 25712 20134 25724
rect 20818 25721 20830 25724
rect 20864 25721 20876 25755
rect 20818 25715 20876 25721
rect 21910 25712 21916 25764
rect 21968 25752 21974 25764
rect 22465 25755 22523 25761
rect 22465 25752 22477 25755
rect 21968 25724 22477 25752
rect 21968 25712 21974 25724
rect 22465 25721 22477 25724
rect 22511 25721 22523 25755
rect 24596 25752 24624 25783
rect 24670 25780 24676 25832
rect 24728 25820 24734 25832
rect 24728 25792 24773 25820
rect 24728 25780 24734 25792
rect 25038 25780 25044 25832
rect 25096 25820 25102 25832
rect 25501 25823 25559 25829
rect 25501 25820 25513 25823
rect 25096 25792 25513 25820
rect 25096 25780 25102 25792
rect 25501 25789 25513 25792
rect 25547 25789 25559 25823
rect 25501 25783 25559 25789
rect 25593 25823 25651 25829
rect 25593 25789 25605 25823
rect 25639 25820 25651 25823
rect 25866 25820 25872 25832
rect 25639 25792 25872 25820
rect 25639 25789 25651 25792
rect 25593 25783 25651 25789
rect 25866 25780 25872 25792
rect 25924 25780 25930 25832
rect 26050 25780 26056 25832
rect 26108 25820 26114 25832
rect 26988 25829 27016 25928
rect 27338 25916 27344 25928
rect 27396 25916 27402 25968
rect 27430 25916 27436 25968
rect 27488 25956 27494 25968
rect 28169 25959 28227 25965
rect 28169 25956 28181 25959
rect 27488 25928 28181 25956
rect 27488 25916 27494 25928
rect 28169 25925 28181 25928
rect 28215 25925 28227 25959
rect 28169 25919 28227 25925
rect 27246 25848 27252 25900
rect 27304 25888 27310 25900
rect 27304 25860 28028 25888
rect 27304 25848 27310 25860
rect 28000 25829 28028 25860
rect 28810 25848 28816 25900
rect 28868 25888 28874 25900
rect 28868 25860 28948 25888
rect 28868 25848 28874 25860
rect 26605 25823 26663 25829
rect 26605 25820 26617 25823
rect 26108 25792 26617 25820
rect 26108 25780 26114 25792
rect 26605 25789 26617 25792
rect 26651 25789 26663 25823
rect 26605 25783 26663 25789
rect 26973 25823 27031 25829
rect 26973 25789 26985 25823
rect 27019 25789 27031 25823
rect 26973 25783 27031 25789
rect 27157 25823 27215 25829
rect 27157 25789 27169 25823
rect 27203 25789 27215 25823
rect 27157 25783 27215 25789
rect 27893 25823 27951 25829
rect 27893 25789 27905 25823
rect 27939 25789 27951 25823
rect 27893 25783 27951 25789
rect 27985 25823 28043 25829
rect 27985 25789 27997 25823
rect 28031 25789 28043 25823
rect 28258 25820 28264 25832
rect 28219 25792 28264 25820
rect 27985 25783 28043 25789
rect 24762 25752 24768 25764
rect 24596 25724 24768 25752
rect 22465 25715 22523 25721
rect 24762 25712 24768 25724
rect 24820 25712 24826 25764
rect 26510 25712 26516 25764
rect 26568 25752 26574 25764
rect 27172 25752 27200 25783
rect 26568 25724 27200 25752
rect 27908 25752 27936 25783
rect 28258 25780 28264 25792
rect 28316 25780 28322 25832
rect 28920 25829 28948 25860
rect 28905 25823 28963 25829
rect 28905 25789 28917 25823
rect 28951 25789 28963 25823
rect 28905 25783 28963 25789
rect 31018 25780 31024 25832
rect 31076 25829 31082 25832
rect 31076 25820 31088 25829
rect 31076 25792 31121 25820
rect 31076 25783 31088 25792
rect 31076 25780 31082 25783
rect 31202 25780 31208 25832
rect 31260 25820 31266 25832
rect 31297 25823 31355 25829
rect 31297 25820 31309 25823
rect 31260 25792 31309 25820
rect 31260 25780 31266 25792
rect 31297 25789 31309 25792
rect 31343 25789 31355 25823
rect 31297 25783 31355 25789
rect 28813 25755 28871 25761
rect 28813 25752 28825 25755
rect 27908 25724 28825 25752
rect 26568 25712 26574 25724
rect 28813 25721 28825 25724
rect 28859 25721 28871 25755
rect 28813 25715 28871 25721
rect 20162 25684 20168 25696
rect 17328 25656 20168 25684
rect 20162 25644 20168 25656
rect 20220 25644 20226 25696
rect 20530 25644 20536 25696
rect 20588 25684 20594 25696
rect 22002 25684 22008 25696
rect 20588 25656 22008 25684
rect 20588 25644 20594 25656
rect 22002 25644 22008 25656
rect 22060 25644 22066 25696
rect 23845 25687 23903 25693
rect 23845 25653 23857 25687
rect 23891 25684 23903 25687
rect 24026 25684 24032 25696
rect 23891 25656 24032 25684
rect 23891 25653 23903 25656
rect 23845 25647 23903 25653
rect 24026 25644 24032 25656
rect 24084 25644 24090 25696
rect 24397 25687 24455 25693
rect 24397 25653 24409 25687
rect 24443 25684 24455 25687
rect 24578 25684 24584 25696
rect 24443 25656 24584 25684
rect 24443 25653 24455 25656
rect 24397 25647 24455 25653
rect 24578 25644 24584 25656
rect 24636 25644 24642 25696
rect 25958 25684 25964 25696
rect 25919 25656 25964 25684
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 26418 25684 26424 25696
rect 26379 25656 26424 25684
rect 26418 25644 26424 25656
rect 26476 25644 26482 25696
rect 29454 25644 29460 25696
rect 29512 25684 29518 25696
rect 29917 25687 29975 25693
rect 29917 25684 29929 25687
rect 29512 25656 29929 25684
rect 29512 25644 29518 25656
rect 29917 25653 29929 25656
rect 29963 25684 29975 25687
rect 30006 25684 30012 25696
rect 29963 25656 30012 25684
rect 29963 25653 29975 25656
rect 29917 25647 29975 25653
rect 30006 25644 30012 25656
rect 30064 25644 30070 25696
rect 1104 25594 32016 25616
rect 0 25548 800 25562
rect 0 25520 1072 25548
rect 1104 25542 11253 25594
rect 11305 25542 11317 25594
rect 11369 25542 11381 25594
rect 11433 25542 11445 25594
rect 11497 25542 11509 25594
rect 11561 25542 21557 25594
rect 21609 25542 21621 25594
rect 21673 25542 21685 25594
rect 21737 25542 21749 25594
rect 21801 25542 21813 25594
rect 21865 25542 32016 25594
rect 32320 25548 33120 25562
rect 1104 25520 32016 25542
rect 32048 25520 33120 25548
rect 0 25506 800 25520
rect 1044 25344 1072 25520
rect 1581 25483 1639 25489
rect 1581 25449 1593 25483
rect 1627 25480 1639 25483
rect 1627 25452 2774 25480
rect 1627 25449 1639 25452
rect 1581 25443 1639 25449
rect 2746 25412 2774 25452
rect 3418 25440 3424 25492
rect 3476 25480 3482 25492
rect 3697 25483 3755 25489
rect 3697 25480 3709 25483
rect 3476 25452 3709 25480
rect 3476 25440 3482 25452
rect 3697 25449 3709 25452
rect 3743 25449 3755 25483
rect 3697 25443 3755 25449
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 5074 25480 5080 25492
rect 4120 25452 5080 25480
rect 4120 25440 4126 25452
rect 5074 25440 5080 25452
rect 5132 25440 5138 25492
rect 5902 25440 5908 25492
rect 5960 25480 5966 25492
rect 6546 25480 6552 25492
rect 5960 25452 6552 25480
rect 5960 25440 5966 25452
rect 6546 25440 6552 25452
rect 6604 25480 6610 25492
rect 6825 25483 6883 25489
rect 6825 25480 6837 25483
rect 6604 25452 6837 25480
rect 6604 25440 6610 25452
rect 6825 25449 6837 25452
rect 6871 25449 6883 25483
rect 6825 25443 6883 25449
rect 13357 25483 13415 25489
rect 13357 25449 13369 25483
rect 13403 25480 13415 25483
rect 13630 25480 13636 25492
rect 13403 25452 13636 25480
rect 13403 25449 13415 25452
rect 13357 25443 13415 25449
rect 13630 25440 13636 25452
rect 13688 25440 13694 25492
rect 15654 25440 15660 25492
rect 15712 25480 15718 25492
rect 16853 25483 16911 25489
rect 16853 25480 16865 25483
rect 15712 25452 16865 25480
rect 15712 25440 15718 25452
rect 16853 25449 16865 25452
rect 16899 25480 16911 25483
rect 17126 25480 17132 25492
rect 16899 25452 17132 25480
rect 16899 25449 16911 25452
rect 16853 25443 16911 25449
rect 17126 25440 17132 25452
rect 17184 25480 17190 25492
rect 17184 25452 18092 25480
rect 17184 25440 17190 25452
rect 3326 25412 3332 25424
rect 2746 25384 3332 25412
rect 3326 25372 3332 25384
rect 3384 25412 3390 25424
rect 5718 25412 5724 25424
rect 3384 25384 5724 25412
rect 3384 25372 3390 25384
rect 5718 25372 5724 25384
rect 5776 25372 5782 25424
rect 8478 25372 8484 25424
rect 8536 25412 8542 25424
rect 9490 25412 9496 25424
rect 8536 25384 9496 25412
rect 8536 25372 8542 25384
rect 9490 25372 9496 25384
rect 9548 25372 9554 25424
rect 9674 25412 9680 25424
rect 9587 25384 9680 25412
rect 9674 25372 9680 25384
rect 9732 25412 9738 25424
rect 10410 25412 10416 25424
rect 9732 25384 10416 25412
rect 9732 25372 9738 25384
rect 10410 25372 10416 25384
rect 10468 25372 10474 25424
rect 10594 25372 10600 25424
rect 10652 25412 10658 25424
rect 10689 25415 10747 25421
rect 10689 25412 10701 25415
rect 10652 25384 10701 25412
rect 10652 25372 10658 25384
rect 10689 25381 10701 25384
rect 10735 25381 10747 25415
rect 10689 25375 10747 25381
rect 12894 25372 12900 25424
rect 12952 25412 12958 25424
rect 13170 25412 13176 25424
rect 12952 25384 13176 25412
rect 12952 25372 12958 25384
rect 13170 25372 13176 25384
rect 13228 25372 13234 25424
rect 17770 25421 17776 25424
rect 13817 25415 13875 25421
rect 13817 25381 13829 25415
rect 13863 25412 13875 25415
rect 17764 25412 17776 25421
rect 13863 25384 15056 25412
rect 17731 25384 17776 25412
rect 13863 25381 13875 25384
rect 13817 25375 13875 25381
rect 1397 25347 1455 25353
rect 1397 25344 1409 25347
rect 1044 25316 1409 25344
rect 1397 25313 1409 25316
rect 1443 25344 1455 25347
rect 2866 25344 2872 25356
rect 1443 25316 2872 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2866 25304 2872 25316
rect 2924 25304 2930 25356
rect 6822 25344 6828 25356
rect 6783 25316 6828 25344
rect 6822 25304 6828 25316
rect 6880 25304 6886 25356
rect 7834 25304 7840 25356
rect 7892 25344 7898 25356
rect 8021 25347 8079 25353
rect 8021 25344 8033 25347
rect 7892 25316 8033 25344
rect 7892 25304 7898 25316
rect 8021 25313 8033 25316
rect 8067 25313 8079 25347
rect 8294 25344 8300 25356
rect 8255 25316 8300 25344
rect 8021 25307 8079 25313
rect 8294 25304 8300 25316
rect 8352 25304 8358 25356
rect 8757 25347 8815 25353
rect 8757 25313 8769 25347
rect 8803 25313 8815 25347
rect 8757 25307 8815 25313
rect 8941 25347 8999 25353
rect 8941 25313 8953 25347
rect 8987 25344 8999 25347
rect 9582 25344 9588 25356
rect 8987 25316 9588 25344
rect 8987 25313 8999 25316
rect 8941 25307 8999 25313
rect 2317 25279 2375 25285
rect 2317 25245 2329 25279
rect 2363 25276 2375 25279
rect 2409 25279 2467 25285
rect 2409 25276 2421 25279
rect 2363 25248 2421 25276
rect 2363 25245 2375 25248
rect 2317 25239 2375 25245
rect 2409 25245 2421 25248
rect 2455 25245 2467 25279
rect 2409 25239 2467 25245
rect 2685 25279 2743 25285
rect 2685 25245 2697 25279
rect 2731 25245 2743 25279
rect 8772 25276 8800 25307
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 10873 25347 10931 25353
rect 10873 25313 10885 25347
rect 10919 25344 10931 25347
rect 11054 25344 11060 25356
rect 10919 25316 11060 25344
rect 10919 25313 10931 25316
rect 10873 25307 10931 25313
rect 11054 25304 11060 25316
rect 11112 25304 11118 25356
rect 11974 25304 11980 25356
rect 12032 25344 12038 25356
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 12032 25316 12817 25344
rect 12032 25304 12038 25316
rect 12805 25313 12817 25316
rect 12851 25313 12863 25347
rect 12805 25307 12863 25313
rect 13446 25304 13452 25356
rect 13504 25344 13510 25356
rect 13630 25344 13636 25356
rect 13504 25316 13636 25344
rect 13504 25304 13510 25316
rect 13630 25304 13636 25316
rect 13688 25304 13694 25356
rect 14001 25347 14059 25353
rect 14001 25313 14013 25347
rect 14047 25313 14059 25347
rect 14182 25344 14188 25356
rect 14143 25316 14188 25344
rect 14001 25307 14059 25313
rect 9030 25276 9036 25288
rect 8772 25248 9036 25276
rect 2685 25239 2743 25245
rect 1946 25168 1952 25220
rect 2004 25208 2010 25220
rect 2700 25208 2728 25239
rect 9030 25236 9036 25248
rect 9088 25236 9094 25288
rect 12066 25276 12072 25288
rect 12027 25248 12072 25276
rect 12066 25236 12072 25248
rect 12124 25236 12130 25288
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25276 12403 25279
rect 13906 25276 13912 25288
rect 12391 25248 13912 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 13906 25236 13912 25248
rect 13964 25236 13970 25288
rect 2004 25180 2728 25208
rect 2004 25168 2010 25180
rect 3694 25168 3700 25220
rect 3752 25208 3758 25220
rect 5169 25211 5227 25217
rect 5169 25208 5181 25211
rect 3752 25180 5181 25208
rect 3752 25168 3758 25180
rect 5169 25177 5181 25180
rect 5215 25177 5227 25211
rect 5169 25171 5227 25177
rect 8941 25211 8999 25217
rect 8941 25177 8953 25211
rect 8987 25208 8999 25211
rect 9766 25208 9772 25220
rect 8987 25180 9772 25208
rect 8987 25177 8999 25180
rect 8941 25171 8999 25177
rect 9766 25168 9772 25180
rect 9824 25168 9830 25220
rect 1486 25100 1492 25152
rect 1544 25140 1550 25152
rect 2317 25143 2375 25149
rect 2317 25140 2329 25143
rect 1544 25112 2329 25140
rect 1544 25100 1550 25112
rect 2317 25109 2329 25112
rect 2363 25140 2375 25143
rect 3418 25140 3424 25152
rect 2363 25112 3424 25140
rect 2363 25109 2375 25112
rect 2317 25103 2375 25109
rect 3418 25100 3424 25112
rect 3476 25100 3482 25152
rect 4338 25100 4344 25152
rect 4396 25140 4402 25152
rect 4617 25143 4675 25149
rect 4617 25140 4629 25143
rect 4396 25112 4629 25140
rect 4396 25100 4402 25112
rect 4617 25109 4629 25112
rect 4663 25109 4675 25143
rect 4617 25103 4675 25109
rect 5258 25100 5264 25152
rect 5316 25140 5322 25152
rect 5721 25143 5779 25149
rect 5721 25140 5733 25143
rect 5316 25112 5733 25140
rect 5316 25100 5322 25112
rect 5721 25109 5733 25112
rect 5767 25140 5779 25143
rect 7742 25140 7748 25152
rect 5767 25112 7748 25140
rect 5767 25109 5779 25112
rect 5721 25103 5779 25109
rect 7742 25100 7748 25112
rect 7800 25100 7806 25152
rect 12710 25100 12716 25152
rect 12768 25140 12774 25152
rect 13173 25143 13231 25149
rect 13173 25140 13185 25143
rect 12768 25112 13185 25140
rect 12768 25100 12774 25112
rect 13173 25109 13185 25112
rect 13219 25109 13231 25143
rect 14016 25140 14044 25307
rect 14182 25304 14188 25316
rect 14240 25304 14246 25356
rect 14366 25344 14372 25356
rect 14327 25316 14372 25344
rect 14366 25304 14372 25316
rect 14424 25304 14430 25356
rect 15028 25353 15056 25384
rect 17764 25375 17776 25384
rect 17770 25372 17776 25375
rect 17828 25372 17834 25424
rect 18064 25412 18092 25452
rect 18138 25440 18144 25492
rect 18196 25480 18202 25492
rect 18877 25483 18935 25489
rect 18877 25480 18889 25483
rect 18196 25452 18889 25480
rect 18196 25440 18202 25452
rect 18877 25449 18889 25452
rect 18923 25449 18935 25483
rect 21266 25480 21272 25492
rect 18877 25443 18935 25449
rect 18984 25452 21272 25480
rect 18984 25412 19012 25452
rect 21266 25440 21272 25452
rect 21324 25440 21330 25492
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25480 23075 25483
rect 24486 25480 24492 25492
rect 23063 25452 24256 25480
rect 24447 25452 24492 25480
rect 23063 25449 23075 25452
rect 23017 25443 23075 25449
rect 18064 25384 19012 25412
rect 20714 25372 20720 25424
rect 20772 25412 20778 25424
rect 24118 25412 24124 25424
rect 20772 25384 24124 25412
rect 20772 25372 20778 25384
rect 14553 25347 14611 25353
rect 14553 25313 14565 25347
rect 14599 25313 14611 25347
rect 14553 25307 14611 25313
rect 15013 25347 15071 25353
rect 15013 25313 15025 25347
rect 15059 25313 15071 25347
rect 15378 25344 15384 25356
rect 15339 25316 15384 25344
rect 15013 25307 15071 25313
rect 14090 25236 14096 25288
rect 14148 25276 14154 25288
rect 14277 25279 14335 25285
rect 14277 25276 14289 25279
rect 14148 25248 14289 25276
rect 14148 25236 14154 25248
rect 14277 25245 14289 25248
rect 14323 25276 14335 25279
rect 14458 25276 14464 25288
rect 14323 25248 14464 25276
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 14568 25276 14596 25307
rect 15378 25304 15384 25316
rect 15436 25304 15442 25356
rect 15841 25347 15899 25353
rect 15841 25344 15853 25347
rect 15764 25316 15853 25344
rect 14642 25276 14648 25288
rect 14568 25248 14648 25276
rect 14642 25236 14648 25248
rect 14700 25276 14706 25288
rect 15562 25276 15568 25288
rect 14700 25248 15568 25276
rect 14700 25236 14706 25248
rect 15562 25236 15568 25248
rect 15620 25236 15626 25288
rect 14182 25168 14188 25220
rect 14240 25208 14246 25220
rect 15764 25208 15792 25316
rect 15841 25313 15853 25316
rect 15887 25344 15899 25347
rect 15930 25344 15936 25356
rect 15887 25316 15936 25344
rect 15887 25313 15899 25316
rect 15841 25307 15899 25313
rect 15930 25304 15936 25316
rect 15988 25304 15994 25356
rect 16669 25347 16727 25353
rect 16669 25313 16681 25347
rect 16715 25313 16727 25347
rect 16669 25307 16727 25313
rect 16684 25276 16712 25307
rect 16758 25304 16764 25356
rect 16816 25344 16822 25356
rect 17497 25347 17555 25353
rect 17497 25344 17509 25347
rect 16816 25316 17509 25344
rect 16816 25304 16822 25316
rect 17497 25313 17509 25316
rect 17543 25313 17555 25347
rect 17497 25307 17555 25313
rect 18782 25304 18788 25356
rect 18840 25344 18846 25356
rect 20450 25347 20508 25353
rect 20450 25344 20462 25347
rect 18840 25316 20462 25344
rect 18840 25304 18846 25316
rect 20450 25313 20462 25316
rect 20496 25313 20508 25347
rect 20450 25307 20508 25313
rect 20990 25304 20996 25356
rect 21048 25344 21054 25356
rect 21821 25347 21879 25353
rect 21821 25344 21833 25347
rect 21048 25316 21833 25344
rect 21048 25304 21054 25316
rect 21821 25313 21833 25316
rect 21867 25313 21879 25347
rect 21821 25307 21879 25313
rect 22005 25347 22063 25353
rect 22005 25313 22017 25347
rect 22051 25313 22063 25347
rect 22005 25307 22063 25313
rect 20717 25279 20775 25285
rect 16684 25248 16988 25276
rect 15930 25208 15936 25220
rect 14240 25180 15792 25208
rect 15891 25180 15936 25208
rect 14240 25168 14246 25180
rect 15930 25168 15936 25180
rect 15988 25168 15994 25220
rect 16960 25152 16988 25248
rect 20717 25245 20729 25279
rect 20763 25245 20775 25279
rect 20717 25239 20775 25245
rect 18598 25168 18604 25220
rect 18656 25208 18662 25220
rect 19337 25211 19395 25217
rect 19337 25208 19349 25211
rect 18656 25180 19349 25208
rect 18656 25168 18662 25180
rect 19337 25177 19349 25180
rect 19383 25177 19395 25211
rect 20732 25208 20760 25239
rect 20898 25236 20904 25288
rect 20956 25276 20962 25288
rect 22020 25276 22048 25307
rect 22278 25304 22284 25356
rect 22336 25344 22342 25356
rect 23124 25353 23152 25384
rect 24118 25372 24124 25384
rect 24176 25372 24182 25424
rect 24228 25412 24256 25452
rect 24486 25440 24492 25452
rect 24544 25440 24550 25492
rect 25958 25440 25964 25492
rect 26016 25480 26022 25492
rect 26211 25483 26269 25489
rect 26211 25480 26223 25483
rect 26016 25452 26223 25480
rect 26016 25440 26022 25452
rect 26211 25449 26223 25452
rect 26257 25449 26269 25483
rect 26211 25443 26269 25449
rect 31297 25483 31355 25489
rect 31297 25449 31309 25483
rect 31343 25480 31355 25483
rect 32048 25480 32076 25520
rect 32320 25506 33120 25520
rect 31343 25452 32076 25480
rect 31343 25449 31355 25452
rect 31297 25443 31355 25449
rect 24228 25384 24532 25412
rect 22373 25347 22431 25353
rect 22373 25344 22385 25347
rect 22336 25316 22385 25344
rect 22336 25304 22342 25316
rect 22373 25313 22385 25316
rect 22419 25344 22431 25347
rect 23017 25347 23075 25353
rect 23017 25344 23029 25347
rect 22419 25316 23029 25344
rect 22419 25313 22431 25316
rect 22373 25307 22431 25313
rect 23017 25313 23029 25316
rect 23063 25313 23075 25347
rect 23017 25307 23075 25313
rect 23109 25347 23167 25353
rect 23109 25313 23121 25347
rect 23155 25313 23167 25347
rect 23109 25307 23167 25313
rect 23376 25347 23434 25353
rect 23376 25313 23388 25347
rect 23422 25344 23434 25347
rect 24394 25344 24400 25356
rect 23422 25316 24400 25344
rect 23422 25313 23434 25316
rect 23376 25307 23434 25313
rect 24394 25304 24400 25316
rect 24452 25304 24458 25356
rect 20956 25248 22048 25276
rect 24504 25276 24532 25384
rect 24762 25372 24768 25424
rect 24820 25412 24826 25424
rect 25216 25415 25274 25421
rect 25216 25412 25228 25415
rect 24820 25384 25228 25412
rect 24820 25372 24826 25384
rect 25216 25381 25228 25384
rect 25262 25412 25274 25415
rect 26421 25415 26479 25421
rect 25262 25384 26096 25412
rect 25262 25381 25274 25384
rect 25216 25375 25274 25381
rect 24946 25344 24952 25356
rect 24907 25316 24952 25344
rect 24946 25304 24952 25316
rect 25004 25304 25010 25356
rect 25038 25304 25044 25356
rect 25096 25344 25102 25356
rect 25314 25344 25320 25356
rect 25096 25316 25320 25344
rect 25096 25304 25102 25316
rect 25314 25304 25320 25316
rect 25372 25304 25378 25356
rect 25406 25304 25412 25356
rect 25464 25344 25470 25356
rect 25593 25347 25651 25353
rect 25593 25344 25605 25347
rect 25464 25316 25605 25344
rect 25464 25304 25470 25316
rect 25593 25313 25605 25316
rect 25639 25313 25651 25347
rect 25593 25307 25651 25313
rect 25866 25276 25872 25288
rect 24504 25248 25872 25276
rect 20956 25236 20962 25248
rect 25866 25236 25872 25248
rect 25924 25236 25930 25288
rect 22094 25208 22100 25220
rect 20732 25180 22100 25208
rect 19337 25171 19395 25177
rect 22094 25168 22100 25180
rect 22152 25168 22158 25220
rect 25958 25208 25964 25220
rect 25056 25180 25964 25208
rect 16758 25140 16764 25152
rect 14016 25112 16764 25140
rect 13173 25103 13231 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 16942 25100 16948 25152
rect 17000 25140 17006 25152
rect 21177 25143 21235 25149
rect 21177 25140 21189 25143
rect 17000 25112 21189 25140
rect 17000 25100 17006 25112
rect 21177 25109 21189 25112
rect 21223 25109 21235 25143
rect 21177 25103 21235 25109
rect 22281 25143 22339 25149
rect 22281 25109 22293 25143
rect 22327 25140 22339 25143
rect 25056 25140 25084 25180
rect 25958 25168 25964 25180
rect 26016 25168 26022 25220
rect 26068 25217 26096 25384
rect 26421 25381 26433 25415
rect 26467 25381 26479 25415
rect 30561 25415 30619 25421
rect 30561 25412 30573 25415
rect 26421 25375 26479 25381
rect 26988 25384 30573 25412
rect 26142 25304 26148 25356
rect 26200 25344 26206 25356
rect 26436 25344 26464 25375
rect 26988 25353 27016 25384
rect 30561 25381 30573 25384
rect 30607 25381 30619 25415
rect 30561 25375 30619 25381
rect 26200 25316 26464 25344
rect 26973 25347 27031 25353
rect 26200 25304 26206 25316
rect 26973 25313 26985 25347
rect 27019 25313 27031 25347
rect 27246 25344 27252 25356
rect 27207 25316 27252 25344
rect 26973 25307 27031 25313
rect 27246 25304 27252 25316
rect 27304 25304 27310 25356
rect 27341 25347 27399 25353
rect 27341 25313 27353 25347
rect 27387 25344 27399 25347
rect 28810 25344 28816 25356
rect 27387 25316 28816 25344
rect 27387 25313 27399 25316
rect 27341 25307 27399 25313
rect 28810 25304 28816 25316
rect 28868 25304 28874 25356
rect 29270 25344 29276 25356
rect 29231 25316 29276 25344
rect 29270 25304 29276 25316
rect 29328 25304 29334 25356
rect 29454 25344 29460 25356
rect 29415 25316 29460 25344
rect 29454 25304 29460 25316
rect 29512 25304 29518 25356
rect 29546 25304 29552 25356
rect 29604 25344 29610 25356
rect 29604 25316 29649 25344
rect 29604 25304 29610 25316
rect 29730 25304 29736 25356
rect 29788 25344 29794 25356
rect 29825 25347 29883 25353
rect 29825 25344 29837 25347
rect 29788 25316 29837 25344
rect 29788 25304 29794 25316
rect 29825 25313 29837 25316
rect 29871 25313 29883 25347
rect 30466 25344 30472 25356
rect 30427 25316 30472 25344
rect 29825 25307 29883 25313
rect 30466 25304 30472 25316
rect 30524 25304 30530 25356
rect 31113 25347 31171 25353
rect 31113 25313 31125 25347
rect 31159 25344 31171 25347
rect 31294 25344 31300 25356
rect 31159 25316 31300 25344
rect 31159 25313 31171 25316
rect 31113 25307 31171 25313
rect 31294 25304 31300 25316
rect 31352 25304 31358 25356
rect 27982 25276 27988 25288
rect 27943 25248 27988 25276
rect 27982 25236 27988 25248
rect 28040 25236 28046 25288
rect 28261 25279 28319 25285
rect 28261 25245 28273 25279
rect 28307 25276 28319 25279
rect 28534 25276 28540 25288
rect 28307 25248 28540 25276
rect 28307 25245 28319 25248
rect 28261 25239 28319 25245
rect 28534 25236 28540 25248
rect 28592 25276 28598 25288
rect 29641 25279 29699 25285
rect 29641 25276 29653 25279
rect 28592 25248 29653 25276
rect 28592 25236 28598 25248
rect 29641 25245 29653 25248
rect 29687 25245 29699 25279
rect 29641 25239 29699 25245
rect 26053 25211 26111 25217
rect 26053 25177 26065 25211
rect 26099 25177 26111 25211
rect 26694 25208 26700 25220
rect 26053 25171 26111 25177
rect 26252 25180 26700 25208
rect 25222 25140 25228 25152
rect 22327 25112 25084 25140
rect 25183 25112 25228 25140
rect 22327 25109 22339 25112
rect 22281 25103 22339 25109
rect 25222 25100 25228 25112
rect 25280 25100 25286 25152
rect 25406 25100 25412 25152
rect 25464 25140 25470 25152
rect 26252 25149 26280 25180
rect 26694 25168 26700 25180
rect 26752 25168 26758 25220
rect 26237 25143 26295 25149
rect 26237 25140 26249 25143
rect 25464 25112 26249 25140
rect 25464 25100 25470 25112
rect 26237 25109 26249 25112
rect 26283 25109 26295 25143
rect 26237 25103 26295 25109
rect 27065 25143 27123 25149
rect 27065 25109 27077 25143
rect 27111 25140 27123 25143
rect 27430 25140 27436 25152
rect 27111 25112 27436 25140
rect 27111 25109 27123 25112
rect 27065 25103 27123 25109
rect 27430 25100 27436 25112
rect 27488 25100 27494 25152
rect 27525 25143 27583 25149
rect 27525 25109 27537 25143
rect 27571 25140 27583 25143
rect 27614 25140 27620 25152
rect 27571 25112 27620 25140
rect 27571 25109 27583 25112
rect 27525 25103 27583 25109
rect 27614 25100 27620 25112
rect 27672 25100 27678 25152
rect 30009 25143 30067 25149
rect 30009 25109 30021 25143
rect 30055 25140 30067 25143
rect 30374 25140 30380 25152
rect 30055 25112 30380 25140
rect 30055 25109 30067 25112
rect 30009 25103 30067 25109
rect 30374 25100 30380 25112
rect 30432 25100 30438 25152
rect 1104 25050 32016 25072
rect 1104 24998 6102 25050
rect 6154 24998 6166 25050
rect 6218 24998 6230 25050
rect 6282 24998 6294 25050
rect 6346 24998 6358 25050
rect 6410 24998 16405 25050
rect 16457 24998 16469 25050
rect 16521 24998 16533 25050
rect 16585 24998 16597 25050
rect 16649 24998 16661 25050
rect 16713 24998 26709 25050
rect 26761 24998 26773 25050
rect 26825 24998 26837 25050
rect 26889 24998 26901 25050
rect 26953 24998 26965 25050
rect 27017 24998 32016 25050
rect 1104 24976 32016 24998
rect 5350 24896 5356 24948
rect 5408 24936 5414 24948
rect 5408 24908 6500 24936
rect 5408 24896 5414 24908
rect 4338 24828 4344 24880
rect 4396 24828 4402 24880
rect 2774 24760 2780 24812
rect 2832 24800 2838 24812
rect 4356 24800 4384 24828
rect 2832 24772 2877 24800
rect 3896 24772 4384 24800
rect 2832 24760 2838 24772
rect 1946 24692 1952 24744
rect 2004 24732 2010 24744
rect 3789 24735 3847 24741
rect 3789 24732 3801 24735
rect 2004 24704 3801 24732
rect 2004 24692 2010 24704
rect 3789 24701 3801 24704
rect 3835 24701 3847 24735
rect 3896 24730 3924 24772
rect 4798 24760 4804 24812
rect 4856 24800 4862 24812
rect 4985 24803 5043 24809
rect 4985 24800 4997 24803
rect 4856 24772 4997 24800
rect 4856 24760 4862 24772
rect 4985 24769 4997 24772
rect 5031 24769 5043 24803
rect 4985 24763 5043 24769
rect 3973 24735 4031 24741
rect 3973 24730 3985 24735
rect 3896 24702 3985 24730
rect 3789 24695 3847 24701
rect 3973 24701 3985 24702
rect 4019 24701 4031 24735
rect 3973 24695 4031 24701
rect 4065 24735 4123 24741
rect 4065 24701 4077 24735
rect 4111 24701 4123 24735
rect 4065 24695 4123 24701
rect 1854 24624 1860 24676
rect 1912 24664 1918 24676
rect 2130 24664 2136 24676
rect 1912 24636 2136 24664
rect 1912 24624 1918 24636
rect 2130 24624 2136 24636
rect 2188 24624 2194 24676
rect 2498 24664 2504 24676
rect 2556 24673 2562 24676
rect 2468 24636 2504 24664
rect 2498 24624 2504 24636
rect 2556 24627 2568 24673
rect 2556 24624 2562 24627
rect 3694 24624 3700 24676
rect 3752 24664 3758 24676
rect 4080 24664 4108 24695
rect 4154 24692 4160 24744
rect 4212 24732 4218 24744
rect 4341 24735 4399 24741
rect 4212 24704 4257 24732
rect 4212 24692 4218 24704
rect 4341 24701 4353 24735
rect 4387 24701 4399 24735
rect 6472 24732 6500 24908
rect 10410 24896 10416 24948
rect 10468 24936 10474 24948
rect 11330 24936 11336 24948
rect 10468 24908 11336 24936
rect 10468 24896 10474 24908
rect 11330 24896 11336 24908
rect 11388 24896 11394 24948
rect 13906 24896 13912 24948
rect 13964 24936 13970 24948
rect 15194 24936 15200 24948
rect 13964 24908 15200 24936
rect 13964 24896 13970 24908
rect 15194 24896 15200 24908
rect 15252 24936 15258 24948
rect 16117 24939 16175 24945
rect 16117 24936 16129 24939
rect 15252 24908 16129 24936
rect 15252 24896 15258 24908
rect 16117 24905 16129 24908
rect 16163 24905 16175 24939
rect 16117 24899 16175 24905
rect 16206 24896 16212 24948
rect 16264 24936 16270 24948
rect 22278 24936 22284 24948
rect 16264 24908 22284 24936
rect 16264 24896 16270 24908
rect 22278 24896 22284 24908
rect 22336 24896 22342 24948
rect 22462 24896 22468 24948
rect 22520 24936 22526 24948
rect 23290 24936 23296 24948
rect 22520 24908 23296 24936
rect 22520 24896 22526 24908
rect 23290 24896 23296 24908
rect 23348 24896 23354 24948
rect 23566 24896 23572 24948
rect 23624 24936 23630 24948
rect 23753 24939 23811 24945
rect 23753 24936 23765 24939
rect 23624 24908 23765 24936
rect 23624 24896 23630 24908
rect 23753 24905 23765 24908
rect 23799 24905 23811 24939
rect 24394 24936 24400 24948
rect 24355 24908 24400 24936
rect 23753 24899 23811 24905
rect 24394 24896 24400 24908
rect 24452 24896 24458 24948
rect 24486 24896 24492 24948
rect 24544 24936 24550 24948
rect 26602 24936 26608 24948
rect 24544 24908 26608 24936
rect 24544 24896 24550 24908
rect 10318 24828 10324 24880
rect 10376 24868 10382 24880
rect 10778 24868 10784 24880
rect 10376 24840 10784 24868
rect 10376 24828 10382 24840
rect 10778 24828 10784 24840
rect 10836 24828 10842 24880
rect 14090 24828 14096 24880
rect 14148 24828 14154 24880
rect 20898 24868 20904 24880
rect 19720 24840 20904 24868
rect 6546 24760 6552 24812
rect 6604 24800 6610 24812
rect 7101 24803 7159 24809
rect 7101 24800 7113 24803
rect 6604 24772 7113 24800
rect 6604 24760 6610 24772
rect 7101 24769 7113 24772
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 7466 24760 7472 24812
rect 7524 24800 7530 24812
rect 8113 24803 8171 24809
rect 8113 24800 8125 24803
rect 7524 24772 8125 24800
rect 7524 24760 7530 24772
rect 8113 24769 8125 24772
rect 8159 24769 8171 24803
rect 8113 24763 8171 24769
rect 9582 24760 9588 24812
rect 9640 24800 9646 24812
rect 9677 24803 9735 24809
rect 9677 24800 9689 24803
rect 9640 24772 9689 24800
rect 9640 24760 9646 24772
rect 9677 24769 9689 24772
rect 9723 24769 9735 24803
rect 9677 24763 9735 24769
rect 10594 24760 10600 24812
rect 10652 24800 10658 24812
rect 11057 24803 11115 24809
rect 11057 24800 11069 24803
rect 10652 24772 11069 24800
rect 10652 24760 10658 24772
rect 11057 24769 11069 24772
rect 11103 24769 11115 24803
rect 11057 24763 11115 24769
rect 12621 24803 12679 24809
rect 12621 24769 12633 24803
rect 12667 24800 12679 24803
rect 14108 24800 14136 24828
rect 12667 24772 14136 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 6825 24735 6883 24741
rect 6825 24732 6837 24735
rect 6472 24704 6837 24732
rect 4341 24695 4399 24701
rect 6825 24701 6837 24704
rect 6871 24732 6883 24735
rect 8018 24732 8024 24744
rect 6871 24704 8024 24732
rect 6871 24701 6883 24704
rect 6825 24695 6883 24701
rect 4356 24664 4384 24695
rect 8018 24692 8024 24704
rect 8076 24732 8082 24744
rect 8297 24735 8355 24741
rect 8297 24732 8309 24735
rect 8076 24704 8309 24732
rect 8076 24692 8082 24704
rect 8297 24701 8309 24704
rect 8343 24701 8355 24735
rect 8297 24695 8355 24701
rect 8754 24692 8760 24744
rect 8812 24732 8818 24744
rect 8941 24735 8999 24741
rect 8941 24732 8953 24735
rect 8812 24704 8953 24732
rect 8812 24692 8818 24704
rect 8941 24701 8953 24704
rect 8987 24732 8999 24735
rect 9490 24732 9496 24744
rect 8987 24704 9496 24732
rect 8987 24701 8999 24704
rect 8941 24695 8999 24701
rect 9490 24692 9496 24704
rect 9548 24692 9554 24744
rect 9769 24735 9827 24741
rect 9769 24701 9781 24735
rect 9815 24732 9827 24735
rect 9950 24732 9956 24744
rect 9815 24704 9956 24732
rect 9815 24701 9827 24704
rect 9769 24695 9827 24701
rect 9950 24692 9956 24704
rect 10008 24732 10014 24744
rect 10226 24732 10232 24744
rect 10008 24704 10232 24732
rect 10008 24692 10014 24704
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 10781 24735 10839 24741
rect 10781 24701 10793 24735
rect 10827 24701 10839 24735
rect 10962 24732 10968 24744
rect 10923 24704 10968 24732
rect 10781 24695 10839 24701
rect 3752 24636 4108 24664
rect 4264 24636 4384 24664
rect 3752 24624 3758 24636
rect 1397 24599 1455 24605
rect 1397 24565 1409 24599
rect 1443 24596 1455 24599
rect 2038 24596 2044 24608
rect 1443 24568 2044 24596
rect 1443 24565 1455 24568
rect 1397 24559 1455 24565
rect 2038 24556 2044 24568
rect 2096 24556 2102 24608
rect 2406 24556 2412 24608
rect 2464 24596 2470 24608
rect 2774 24596 2780 24608
rect 2464 24568 2780 24596
rect 2464 24556 2470 24568
rect 2774 24556 2780 24568
rect 2832 24556 2838 24608
rect 3510 24556 3516 24608
rect 3568 24596 3574 24608
rect 4264 24596 4292 24636
rect 5074 24624 5080 24676
rect 5132 24664 5138 24676
rect 5230 24667 5288 24673
rect 5230 24664 5242 24667
rect 5132 24636 5242 24664
rect 5132 24624 5138 24636
rect 5230 24633 5242 24636
rect 5276 24633 5288 24667
rect 10796 24664 10824 24695
rect 10962 24692 10968 24704
rect 11020 24692 11026 24744
rect 11146 24732 11152 24744
rect 11107 24704 11152 24732
rect 11146 24692 11152 24704
rect 11204 24692 11210 24744
rect 11330 24732 11336 24744
rect 11291 24704 11336 24732
rect 11330 24692 11336 24704
rect 11388 24732 11394 24744
rect 12342 24732 12348 24744
rect 11388 24704 12348 24732
rect 11388 24692 11394 24704
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 12526 24732 12532 24744
rect 12487 24704 12532 24732
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 12066 24664 12072 24676
rect 10796 24636 12072 24664
rect 5230 24627 5288 24633
rect 12066 24624 12072 24636
rect 12124 24624 12130 24676
rect 4522 24596 4528 24608
rect 3568 24568 4292 24596
rect 4483 24568 4528 24596
rect 3568 24556 3574 24568
rect 4522 24556 4528 24568
rect 4580 24556 4586 24608
rect 6362 24596 6368 24608
rect 6323 24568 6368 24596
rect 6362 24556 6368 24568
rect 6420 24556 6426 24608
rect 9030 24596 9036 24608
rect 8991 24568 9036 24596
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 10321 24599 10379 24605
rect 10321 24565 10333 24599
rect 10367 24596 10379 24599
rect 10778 24596 10784 24608
rect 10367 24568 10784 24596
rect 10367 24565 10379 24568
rect 10321 24559 10379 24565
rect 10778 24556 10784 24568
rect 10836 24556 10842 24608
rect 11517 24599 11575 24605
rect 11517 24565 11529 24599
rect 11563 24596 11575 24599
rect 11698 24596 11704 24608
rect 11563 24568 11704 24596
rect 11563 24565 11575 24568
rect 11517 24559 11575 24565
rect 11698 24556 11704 24568
rect 11756 24556 11762 24608
rect 11790 24556 11796 24608
rect 11848 24596 11854 24608
rect 12636 24596 12664 24763
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 19720 24809 19748 24840
rect 20898 24828 20904 24840
rect 20956 24828 20962 24880
rect 23198 24868 23204 24880
rect 23159 24840 23204 24868
rect 23198 24828 23204 24840
rect 23256 24828 23262 24880
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 18380 24772 19717 24800
rect 18380 24760 18386 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 20070 24800 20076 24812
rect 20031 24772 20076 24800
rect 19705 24763 19763 24769
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20438 24760 20444 24812
rect 20496 24800 20502 24812
rect 20625 24803 20683 24809
rect 20625 24800 20637 24803
rect 20496 24772 20637 24800
rect 20496 24760 20502 24772
rect 20625 24769 20637 24772
rect 20671 24769 20683 24803
rect 20625 24763 20683 24769
rect 22649 24803 22707 24809
rect 22649 24769 22661 24803
rect 22695 24800 22707 24803
rect 22738 24800 22744 24812
rect 22695 24772 22744 24800
rect 22695 24769 22707 24772
rect 22649 24763 22707 24769
rect 22738 24760 22744 24772
rect 22796 24760 22802 24812
rect 25130 24800 25136 24812
rect 25091 24772 25136 24800
rect 25130 24760 25136 24772
rect 25188 24760 25194 24812
rect 25424 24809 25452 24908
rect 25409 24803 25467 24809
rect 25409 24769 25421 24803
rect 25455 24769 25467 24803
rect 25409 24763 25467 24769
rect 25501 24803 25559 24809
rect 25501 24769 25513 24803
rect 25547 24800 25559 24803
rect 26237 24803 26295 24809
rect 25547 24772 25748 24800
rect 25547 24769 25559 24772
rect 25501 24763 25559 24769
rect 12713 24735 12771 24741
rect 12713 24701 12725 24735
rect 12759 24732 12771 24735
rect 12802 24732 12808 24744
rect 12759 24704 12808 24732
rect 12759 24701 12771 24704
rect 12713 24695 12771 24701
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 12897 24735 12955 24741
rect 12897 24701 12909 24735
rect 12943 24732 12955 24735
rect 13446 24732 13452 24744
rect 12943 24704 13452 24732
rect 12943 24701 12955 24704
rect 12897 24695 12955 24701
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 13538 24692 13544 24744
rect 13596 24732 13602 24744
rect 14093 24735 14151 24741
rect 14093 24732 14105 24735
rect 13596 24704 14105 24732
rect 13596 24692 13602 24704
rect 14093 24701 14105 24704
rect 14139 24701 14151 24735
rect 14093 24695 14151 24701
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 17678 24732 17684 24744
rect 14792 24704 17684 24732
rect 14792 24692 14798 24704
rect 17678 24692 17684 24704
rect 17736 24692 17742 24744
rect 18690 24732 18696 24744
rect 18651 24704 18696 24732
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 19334 24692 19340 24744
rect 19392 24732 19398 24744
rect 19521 24735 19579 24741
rect 19392 24704 19437 24732
rect 19392 24692 19398 24704
rect 19521 24701 19533 24735
rect 19567 24701 19579 24735
rect 19521 24695 19579 24701
rect 14360 24667 14418 24673
rect 14360 24633 14372 24667
rect 14406 24664 14418 24667
rect 14458 24664 14464 24676
rect 14406 24636 14464 24664
rect 14406 24633 14418 24636
rect 14360 24627 14418 24633
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 15102 24624 15108 24676
rect 15160 24664 15166 24676
rect 16025 24667 16083 24673
rect 16025 24664 16037 24667
rect 15160 24636 16037 24664
rect 15160 24624 15166 24636
rect 16025 24633 16037 24636
rect 16071 24633 16083 24667
rect 17034 24664 17040 24676
rect 16995 24636 17040 24664
rect 16025 24627 16083 24633
rect 17034 24624 17040 24636
rect 17092 24624 17098 24676
rect 19536 24664 19564 24695
rect 19610 24692 19616 24744
rect 19668 24732 19674 24744
rect 19668 24704 19713 24732
rect 19668 24692 19674 24704
rect 19794 24692 19800 24744
rect 19852 24732 19858 24744
rect 19889 24735 19947 24741
rect 19889 24732 19901 24735
rect 19852 24704 19901 24732
rect 19852 24692 19858 24704
rect 19889 24701 19901 24704
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 20717 24735 20775 24741
rect 20717 24701 20729 24735
rect 20763 24732 20775 24735
rect 20806 24732 20812 24744
rect 20763 24704 20812 24732
rect 20763 24701 20775 24704
rect 20717 24695 20775 24701
rect 20732 24664 20760 24695
rect 20806 24692 20812 24704
rect 20864 24692 20870 24744
rect 22382 24735 22440 24741
rect 22382 24732 22394 24735
rect 22066 24704 22394 24732
rect 21082 24664 21088 24676
rect 19536 24636 21088 24664
rect 21082 24624 21088 24636
rect 21140 24664 21146 24676
rect 21140 24636 21312 24664
rect 21140 24624 21146 24636
rect 11848 24568 12664 24596
rect 11848 24556 11854 24568
rect 12986 24556 12992 24608
rect 13044 24596 13050 24608
rect 13081 24599 13139 24605
rect 13081 24596 13093 24599
rect 13044 24568 13093 24596
rect 13044 24556 13050 24568
rect 13081 24565 13093 24568
rect 13127 24565 13139 24599
rect 13081 24559 13139 24565
rect 15473 24599 15531 24605
rect 15473 24565 15485 24599
rect 15519 24596 15531 24599
rect 15562 24596 15568 24608
rect 15519 24568 15568 24596
rect 15519 24565 15531 24568
rect 15473 24559 15531 24565
rect 15562 24556 15568 24568
rect 15620 24556 15626 24608
rect 21284 24605 21312 24636
rect 21358 24624 21364 24676
rect 21416 24664 21422 24676
rect 22066 24664 22094 24704
rect 22382 24701 22394 24704
rect 22428 24701 22440 24735
rect 22382 24695 22440 24701
rect 23106 24692 23112 24744
rect 23164 24732 23170 24744
rect 23293 24735 23351 24741
rect 23293 24732 23305 24735
rect 23164 24704 23305 24732
rect 23164 24692 23170 24704
rect 23293 24701 23305 24704
rect 23339 24701 23351 24735
rect 24578 24732 24584 24744
rect 24539 24704 24584 24732
rect 23293 24695 23351 24701
rect 24578 24692 24584 24704
rect 24636 24692 24642 24744
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24732 25099 24735
rect 25317 24735 25375 24741
rect 25317 24732 25329 24735
rect 25087 24704 25329 24732
rect 25087 24701 25099 24704
rect 25041 24695 25099 24701
rect 25317 24701 25329 24704
rect 25363 24701 25375 24735
rect 25317 24695 25375 24701
rect 25593 24735 25651 24741
rect 25593 24701 25605 24735
rect 25639 24701 25651 24735
rect 25593 24695 25651 24701
rect 24118 24664 24124 24676
rect 21416 24636 22094 24664
rect 22397 24636 24124 24664
rect 21416 24624 21422 24636
rect 21269 24599 21327 24605
rect 21269 24565 21281 24599
rect 21315 24565 21327 24599
rect 21269 24559 21327 24565
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 22397 24596 22425 24636
rect 24118 24624 24124 24636
rect 24176 24624 24182 24676
rect 24946 24624 24952 24676
rect 25004 24664 25010 24676
rect 25608 24664 25636 24695
rect 25004 24636 25636 24664
rect 25720 24664 25748 24772
rect 26237 24769 26249 24803
rect 26283 24769 26295 24803
rect 26344 24800 26372 24908
rect 26602 24896 26608 24908
rect 26660 24896 26666 24948
rect 26418 24828 26424 24880
rect 26476 24868 26482 24880
rect 26476 24840 26740 24868
rect 26476 24828 26482 24840
rect 26712 24809 26740 24840
rect 26513 24803 26571 24809
rect 26513 24800 26525 24803
rect 26344 24772 26525 24800
rect 26237 24763 26295 24769
rect 26513 24769 26525 24772
rect 26559 24769 26571 24803
rect 26513 24763 26571 24769
rect 26697 24803 26755 24809
rect 26697 24769 26709 24803
rect 26743 24769 26755 24803
rect 26697 24763 26755 24769
rect 25777 24735 25835 24741
rect 25777 24701 25789 24735
rect 25823 24732 25835 24735
rect 26252 24732 26280 24763
rect 27522 24760 27528 24812
rect 27580 24800 27586 24812
rect 27893 24803 27951 24809
rect 27893 24800 27905 24803
rect 27580 24772 27905 24800
rect 27580 24760 27586 24772
rect 27893 24769 27905 24772
rect 27939 24769 27951 24803
rect 27893 24763 27951 24769
rect 27985 24803 28043 24809
rect 27985 24769 27997 24803
rect 28031 24800 28043 24803
rect 28074 24800 28080 24812
rect 28031 24772 28080 24800
rect 28031 24769 28043 24772
rect 27985 24763 28043 24769
rect 25823 24704 26280 24732
rect 25823 24701 25835 24704
rect 25777 24695 25835 24701
rect 26418 24692 26424 24744
rect 26476 24732 26482 24744
rect 26476 24704 26521 24732
rect 26476 24692 26482 24704
rect 26602 24692 26608 24744
rect 26660 24732 26666 24744
rect 26881 24735 26939 24741
rect 26660 24704 26705 24732
rect 26660 24692 26666 24704
rect 26881 24701 26893 24735
rect 26927 24732 26939 24735
rect 27062 24732 27068 24744
rect 26927 24704 27068 24732
rect 26927 24701 26939 24704
rect 26881 24695 26939 24701
rect 27062 24692 27068 24704
rect 27120 24692 27126 24744
rect 27614 24732 27620 24744
rect 27575 24704 27620 24732
rect 27614 24692 27620 24704
rect 27672 24692 27678 24744
rect 27798 24732 27804 24744
rect 27759 24704 27804 24732
rect 27798 24692 27804 24704
rect 27856 24692 27862 24744
rect 26234 24664 26240 24676
rect 25720 24636 26240 24664
rect 25004 24624 25010 24636
rect 26234 24624 26240 24636
rect 26292 24624 26298 24676
rect 27154 24664 27160 24676
rect 26629 24636 27160 24664
rect 21968 24568 22425 24596
rect 21968 24556 21974 24568
rect 22462 24556 22468 24608
rect 22520 24596 22526 24608
rect 23382 24596 23388 24608
rect 22520 24568 23388 24596
rect 22520 24556 22526 24568
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 25041 24599 25099 24605
rect 25041 24565 25053 24599
rect 25087 24596 25099 24599
rect 26629 24596 26657 24636
rect 27154 24624 27160 24636
rect 27212 24624 27218 24676
rect 27338 24624 27344 24676
rect 27396 24664 27402 24676
rect 28000 24664 28028 24763
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24800 30987 24803
rect 31202 24800 31208 24812
rect 30975 24772 31208 24800
rect 30975 24769 30987 24772
rect 30929 24763 30987 24769
rect 31202 24760 31208 24772
rect 31260 24760 31266 24812
rect 28169 24735 28227 24741
rect 28169 24701 28181 24735
rect 28215 24732 28227 24735
rect 28905 24735 28963 24741
rect 28905 24732 28917 24735
rect 28215 24704 28917 24732
rect 28215 24701 28227 24704
rect 28169 24695 28227 24701
rect 28905 24701 28917 24704
rect 28951 24701 28963 24735
rect 28905 24695 28963 24701
rect 28994 24692 29000 24744
rect 29052 24732 29058 24744
rect 29052 24704 29097 24732
rect 29052 24692 29058 24704
rect 30374 24692 30380 24744
rect 30432 24732 30438 24744
rect 30662 24735 30720 24741
rect 30662 24732 30674 24735
rect 30432 24704 30674 24732
rect 30432 24692 30438 24704
rect 30662 24701 30674 24704
rect 30708 24701 30720 24735
rect 30662 24695 30720 24701
rect 27396 24636 28028 24664
rect 27396 24624 27402 24636
rect 25087 24568 26657 24596
rect 25087 24565 25099 24568
rect 25041 24559 25099 24565
rect 26694 24556 26700 24608
rect 26752 24596 26758 24608
rect 28353 24599 28411 24605
rect 28353 24596 28365 24599
rect 26752 24568 28365 24596
rect 26752 24556 26758 24568
rect 28353 24565 28365 24568
rect 28399 24565 28411 24599
rect 28353 24559 28411 24565
rect 28994 24556 29000 24608
rect 29052 24596 29058 24608
rect 29549 24599 29607 24605
rect 29549 24596 29561 24599
rect 29052 24568 29561 24596
rect 29052 24556 29058 24568
rect 29549 24565 29561 24568
rect 29595 24596 29607 24599
rect 29730 24596 29736 24608
rect 29595 24568 29736 24596
rect 29595 24565 29607 24568
rect 29549 24559 29607 24565
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 1104 24506 32016 24528
rect 1104 24454 11253 24506
rect 11305 24454 11317 24506
rect 11369 24454 11381 24506
rect 11433 24454 11445 24506
rect 11497 24454 11509 24506
rect 11561 24454 21557 24506
rect 21609 24454 21621 24506
rect 21673 24454 21685 24506
rect 21737 24454 21749 24506
rect 21801 24454 21813 24506
rect 21865 24454 32016 24506
rect 1104 24432 32016 24454
rect 1946 24392 1952 24404
rect 1872 24364 1952 24392
rect 1872 24265 1900 24364
rect 1946 24352 1952 24364
rect 2004 24352 2010 24404
rect 2038 24352 2044 24404
rect 2096 24352 2102 24404
rect 2498 24352 2504 24404
rect 2556 24392 2562 24404
rect 2593 24395 2651 24401
rect 2593 24392 2605 24395
rect 2556 24364 2605 24392
rect 2556 24352 2562 24364
rect 2593 24361 2605 24364
rect 2639 24361 2651 24395
rect 5074 24392 5080 24404
rect 5035 24364 5080 24392
rect 2593 24355 2651 24361
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 7926 24352 7932 24404
rect 7984 24392 7990 24404
rect 7984 24364 8064 24392
rect 7984 24352 7990 24364
rect 2056 24324 2084 24352
rect 4154 24324 4160 24336
rect 2056 24296 2452 24324
rect 1857 24259 1915 24265
rect 1857 24225 1869 24259
rect 1903 24225 1915 24259
rect 2038 24256 2044 24268
rect 1999 24228 2044 24256
rect 1857 24219 1915 24225
rect 2038 24216 2044 24228
rect 2096 24216 2102 24268
rect 2424 24265 2452 24296
rect 3896 24296 4160 24324
rect 2409 24259 2467 24265
rect 2409 24225 2421 24259
rect 2455 24225 2467 24259
rect 2409 24219 2467 24225
rect 2130 24188 2136 24200
rect 2091 24160 2136 24188
rect 2130 24148 2136 24160
rect 2188 24148 2194 24200
rect 3896 24197 3924 24296
rect 4154 24284 4160 24296
rect 4212 24284 4218 24336
rect 4798 24284 4804 24336
rect 4856 24324 4862 24336
rect 8036 24324 8064 24364
rect 8110 24352 8116 24404
rect 8168 24392 8174 24404
rect 10781 24395 10839 24401
rect 8168 24364 10732 24392
rect 8168 24352 8174 24364
rect 9490 24324 9496 24336
rect 4856 24296 7972 24324
rect 8036 24296 9076 24324
rect 4856 24284 4862 24296
rect 5261 24259 5319 24265
rect 5261 24225 5273 24259
rect 5307 24256 5319 24259
rect 5307 24228 5396 24256
rect 5307 24225 5319 24228
rect 5261 24219 5319 24225
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 3881 24191 3939 24197
rect 3881 24188 3893 24191
rect 2271 24160 3893 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 3881 24157 3893 24160
rect 3927 24157 3939 24191
rect 4154 24188 4160 24200
rect 4115 24160 4160 24188
rect 3881 24151 3939 24157
rect 4154 24148 4160 24160
rect 4212 24148 4218 24200
rect 2038 24080 2044 24132
rect 2096 24120 2102 24132
rect 4246 24120 4252 24132
rect 2096 24092 4252 24120
rect 2096 24080 2102 24092
rect 4246 24080 4252 24092
rect 4304 24080 4310 24132
rect 5368 24120 5396 24228
rect 5442 24216 5448 24268
rect 5500 24256 5506 24268
rect 5626 24256 5632 24268
rect 5500 24228 5545 24256
rect 5587 24228 5632 24256
rect 5500 24216 5506 24228
rect 5626 24216 5632 24228
rect 5684 24216 5690 24268
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 5994 24256 6000 24268
rect 5859 24228 6000 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 5994 24216 6000 24228
rect 6052 24216 6058 24268
rect 7673 24259 7731 24265
rect 7673 24225 7685 24259
rect 7719 24256 7731 24259
rect 7834 24256 7840 24268
rect 7719 24228 7840 24256
rect 7719 24225 7731 24228
rect 7673 24219 7731 24225
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 7944 24265 7972 24296
rect 9048 24265 9076 24296
rect 9223 24296 9496 24324
rect 7929 24259 7987 24265
rect 7929 24225 7941 24259
rect 7975 24225 7987 24259
rect 8941 24259 8999 24265
rect 8941 24256 8953 24259
rect 8936 24254 8953 24256
rect 7929 24219 7987 24225
rect 8864 24226 8953 24254
rect 5537 24191 5595 24197
rect 5537 24157 5549 24191
rect 5583 24188 5595 24191
rect 6546 24188 6552 24200
rect 5583 24160 6552 24188
rect 5583 24157 5595 24160
rect 5537 24151 5595 24157
rect 6546 24148 6552 24160
rect 6604 24148 6610 24200
rect 8570 24148 8576 24200
rect 8628 24188 8634 24200
rect 8665 24191 8723 24197
rect 8665 24188 8677 24191
rect 8628 24160 8677 24188
rect 8628 24148 8634 24160
rect 8665 24157 8677 24160
rect 8711 24157 8723 24191
rect 8665 24151 8723 24157
rect 5810 24120 5816 24132
rect 5368 24092 5816 24120
rect 5810 24080 5816 24092
rect 5868 24120 5874 24132
rect 6362 24120 6368 24132
rect 5868 24092 6368 24120
rect 5868 24080 5874 24092
rect 6362 24080 6368 24092
rect 6420 24080 6426 24132
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 7006 24052 7012 24064
rect 6595 24024 7012 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 7006 24012 7012 24024
rect 7064 24012 7070 24064
rect 8864 24052 8892 24226
rect 8941 24225 8953 24226
rect 8987 24225 8999 24259
rect 8941 24219 8999 24225
rect 9033 24259 9091 24265
rect 9033 24225 9045 24259
rect 9079 24225 9091 24259
rect 9033 24219 9091 24225
rect 9125 24259 9183 24265
rect 9125 24225 9137 24259
rect 9171 24258 9183 24259
rect 9223 24258 9251 24296
rect 9490 24284 9496 24296
rect 9548 24324 9554 24336
rect 9548 24296 9812 24324
rect 9548 24284 9554 24296
rect 9171 24230 9251 24258
rect 9309 24259 9367 24265
rect 9171 24225 9183 24230
rect 9125 24219 9183 24225
rect 9309 24225 9321 24259
rect 9355 24256 9367 24259
rect 9582 24256 9588 24268
rect 9355 24228 9588 24256
rect 9355 24225 9367 24228
rect 9309 24219 9367 24225
rect 9582 24216 9588 24228
rect 9640 24216 9646 24268
rect 9784 24265 9812 24296
rect 9769 24259 9827 24265
rect 9769 24225 9781 24259
rect 9815 24225 9827 24259
rect 9950 24256 9956 24268
rect 9911 24228 9956 24256
rect 9769 24219 9827 24225
rect 9950 24216 9956 24228
rect 10008 24216 10014 24268
rect 10704 24188 10732 24364
rect 10781 24361 10793 24395
rect 10827 24392 10839 24395
rect 11146 24392 11152 24404
rect 10827 24364 11152 24392
rect 10827 24361 10839 24364
rect 10781 24355 10839 24361
rect 11146 24352 11152 24364
rect 11204 24352 11210 24404
rect 15286 24352 15292 24404
rect 15344 24392 15350 24404
rect 16022 24392 16028 24404
rect 15344 24364 16028 24392
rect 15344 24352 15350 24364
rect 16022 24352 16028 24364
rect 16080 24352 16086 24404
rect 18693 24395 18751 24401
rect 18693 24361 18705 24395
rect 18739 24392 18751 24395
rect 18782 24392 18788 24404
rect 18739 24364 18788 24392
rect 18739 24361 18751 24364
rect 18693 24355 18751 24361
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 19334 24352 19340 24404
rect 19392 24352 19398 24404
rect 19518 24352 19524 24404
rect 19576 24392 19582 24404
rect 21269 24395 21327 24401
rect 19576 24364 21220 24392
rect 19576 24352 19582 24364
rect 10962 24284 10968 24336
rect 11020 24324 11026 24336
rect 12526 24324 12532 24336
rect 11020 24296 12532 24324
rect 11020 24284 11026 24296
rect 12526 24284 12532 24296
rect 12584 24324 12590 24336
rect 12710 24324 12716 24336
rect 12584 24296 12716 24324
rect 12584 24284 12590 24296
rect 12710 24284 12716 24296
rect 12768 24284 12774 24336
rect 13262 24284 13268 24336
rect 13320 24324 13326 24336
rect 15102 24324 15108 24336
rect 13320 24296 15108 24324
rect 13320 24284 13326 24296
rect 15102 24284 15108 24296
rect 15160 24324 15166 24336
rect 15381 24327 15439 24333
rect 15381 24324 15393 24327
rect 15160 24296 15393 24324
rect 15160 24284 15166 24296
rect 15381 24293 15393 24296
rect 15427 24293 15439 24327
rect 19352 24324 19380 24352
rect 15381 24287 15439 24293
rect 17972 24296 20576 24324
rect 10778 24216 10784 24268
rect 10836 24256 10842 24268
rect 10873 24259 10931 24265
rect 10873 24256 10885 24259
rect 10836 24228 10885 24256
rect 10836 24216 10842 24228
rect 10873 24225 10885 24228
rect 10919 24225 10931 24259
rect 10873 24219 10931 24225
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11514 24256 11520 24268
rect 11112 24228 11520 24256
rect 11112 24216 11118 24228
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 12986 24256 12992 24268
rect 12947 24228 12992 24256
rect 12986 24216 12992 24228
rect 13044 24216 13050 24268
rect 13170 24256 13176 24268
rect 13131 24228 13176 24256
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 13725 24259 13783 24265
rect 13725 24225 13737 24259
rect 13771 24256 13783 24259
rect 13814 24256 13820 24268
rect 13771 24228 13820 24256
rect 13771 24225 13783 24228
rect 13725 24219 13783 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 14182 24216 14188 24268
rect 14240 24256 14246 24268
rect 14369 24259 14427 24265
rect 14369 24256 14381 24259
rect 14240 24228 14381 24256
rect 14240 24216 14246 24228
rect 14369 24225 14381 24228
rect 14415 24256 14427 24259
rect 16942 24256 16948 24268
rect 14415 24228 16948 24256
rect 14415 24225 14427 24228
rect 14369 24219 14427 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17221 24259 17279 24265
rect 17221 24225 17233 24259
rect 17267 24256 17279 24259
rect 17402 24256 17408 24268
rect 17267 24228 17408 24256
rect 17267 24225 17279 24228
rect 17221 24219 17279 24225
rect 17402 24216 17408 24228
rect 17460 24216 17466 24268
rect 17972 24265 18000 24296
rect 17957 24259 18015 24265
rect 17957 24225 17969 24259
rect 18003 24225 18015 24259
rect 18138 24256 18144 24268
rect 18099 24228 18144 24256
rect 17957 24219 18015 24225
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 18230 24216 18236 24268
rect 18288 24256 18294 24268
rect 18509 24259 18567 24265
rect 18288 24228 18333 24256
rect 18288 24216 18294 24228
rect 18509 24225 18521 24259
rect 18555 24256 18567 24259
rect 18598 24256 18604 24268
rect 18555 24228 18604 24256
rect 18555 24225 18567 24228
rect 18509 24219 18567 24225
rect 18598 24216 18604 24228
rect 18656 24216 18662 24268
rect 19426 24256 19432 24268
rect 19387 24228 19432 24256
rect 19426 24216 19432 24228
rect 19484 24216 19490 24268
rect 19797 24259 19855 24265
rect 19797 24256 19809 24259
rect 19536 24228 19809 24256
rect 14642 24188 14648 24200
rect 10704 24160 13952 24188
rect 14603 24160 14648 24188
rect 11606 24080 11612 24132
rect 11664 24120 11670 24132
rect 13633 24123 13691 24129
rect 11664 24092 13400 24120
rect 11664 24080 11670 24092
rect 9214 24052 9220 24064
rect 8864 24024 9220 24052
rect 9214 24012 9220 24024
rect 9272 24012 9278 24064
rect 9950 24052 9956 24064
rect 9911 24024 9956 24052
rect 9950 24012 9956 24024
rect 10008 24012 10014 24064
rect 10594 24012 10600 24064
rect 10652 24052 10658 24064
rect 11054 24052 11060 24064
rect 10652 24024 11060 24052
rect 10652 24012 10658 24024
rect 11054 24012 11060 24024
rect 11112 24052 11118 24064
rect 11747 24055 11805 24061
rect 11747 24052 11759 24055
rect 11112 24024 11759 24052
rect 11112 24012 11118 24024
rect 11747 24021 11759 24024
rect 11793 24021 11805 24055
rect 13372 24052 13400 24092
rect 13633 24089 13645 24123
rect 13679 24089 13691 24123
rect 13924 24120 13952 24160
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 15565 24191 15623 24197
rect 15565 24157 15577 24191
rect 15611 24188 15623 24191
rect 16206 24188 16212 24200
rect 15611 24160 16212 24188
rect 15611 24157 15623 24160
rect 15565 24151 15623 24157
rect 16206 24148 16212 24160
rect 16264 24188 16270 24200
rect 17497 24191 17555 24197
rect 17497 24188 17509 24191
rect 16264 24160 17509 24188
rect 16264 24148 16270 24160
rect 17497 24157 17509 24160
rect 17543 24157 17555 24191
rect 18322 24188 18328 24200
rect 18283 24160 18328 24188
rect 17497 24151 17555 24157
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 19150 24148 19156 24200
rect 19208 24188 19214 24200
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 19208 24160 19257 24188
rect 19208 24148 19214 24160
rect 19245 24157 19257 24160
rect 19291 24157 19303 24191
rect 19245 24151 19303 24157
rect 18782 24120 18788 24132
rect 13924 24092 18788 24120
rect 13633 24083 13691 24089
rect 13648 24052 13676 24083
rect 18782 24080 18788 24092
rect 18840 24080 18846 24132
rect 13372 24024 13676 24052
rect 11747 24015 11805 24021
rect 16298 24012 16304 24064
rect 16356 24052 16362 24064
rect 19536 24052 19564 24228
rect 19797 24225 19809 24228
rect 19843 24256 19855 24259
rect 19886 24256 19892 24268
rect 19843 24228 19892 24256
rect 19843 24225 19855 24228
rect 19797 24219 19855 24225
rect 19886 24216 19892 24228
rect 19944 24216 19950 24268
rect 20548 24265 20576 24296
rect 20806 24284 20812 24336
rect 20864 24284 20870 24336
rect 21192 24324 21220 24364
rect 21269 24361 21281 24395
rect 21315 24392 21327 24395
rect 21358 24392 21364 24404
rect 21315 24364 21364 24392
rect 21315 24361 21327 24364
rect 21269 24355 21327 24361
rect 21358 24352 21364 24364
rect 21416 24352 21422 24404
rect 21913 24395 21971 24401
rect 21913 24361 21925 24395
rect 21959 24392 21971 24395
rect 23842 24392 23848 24404
rect 21959 24364 23848 24392
rect 21959 24361 21971 24364
rect 21913 24355 21971 24361
rect 23842 24352 23848 24364
rect 23900 24352 23906 24404
rect 23937 24395 23995 24401
rect 23937 24361 23949 24395
rect 23983 24392 23995 24395
rect 24118 24392 24124 24404
rect 23983 24364 24124 24392
rect 23983 24361 23995 24364
rect 23937 24355 23995 24361
rect 24118 24352 24124 24364
rect 24176 24352 24182 24404
rect 26418 24392 26424 24404
rect 26252 24364 26424 24392
rect 23382 24324 23388 24336
rect 21192 24296 23388 24324
rect 20533 24259 20591 24265
rect 20533 24225 20545 24259
rect 20579 24256 20591 24259
rect 20622 24256 20628 24268
rect 20579 24228 20628 24256
rect 20579 24225 20591 24228
rect 20533 24219 20591 24225
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 20717 24259 20775 24265
rect 20717 24225 20729 24259
rect 20763 24256 20775 24259
rect 20824 24256 20852 24284
rect 20763 24228 20852 24256
rect 20763 24225 20775 24228
rect 20717 24219 20775 24225
rect 20898 24216 20904 24268
rect 20956 24256 20962 24268
rect 20956 24228 21001 24256
rect 20956 24216 20962 24228
rect 21082 24216 21088 24268
rect 21140 24256 21146 24268
rect 22373 24259 22431 24265
rect 21140 24228 21185 24256
rect 21140 24216 21146 24228
rect 22373 24225 22385 24259
rect 22419 24225 22431 24259
rect 22373 24219 22431 24225
rect 19610 24148 19616 24200
rect 19668 24188 19674 24200
rect 19978 24188 19984 24200
rect 19668 24160 19984 24188
rect 19668 24148 19674 24160
rect 19978 24148 19984 24160
rect 20036 24188 20042 24200
rect 20818 24191 20876 24197
rect 20818 24188 20830 24191
rect 20036 24160 20830 24188
rect 20036 24148 20042 24160
rect 20818 24157 20830 24160
rect 20864 24157 20876 24191
rect 20818 24151 20876 24157
rect 19705 24123 19763 24129
rect 19705 24089 19717 24123
rect 19751 24120 19763 24123
rect 22278 24120 22284 24132
rect 19751 24092 22284 24120
rect 19751 24089 19763 24092
rect 19705 24083 19763 24089
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 16356 24024 19564 24052
rect 16356 24012 16362 24024
rect 21542 24012 21548 24064
rect 21600 24052 21606 24064
rect 22397 24052 22425 24219
rect 22480 24188 22508 24296
rect 23382 24284 23388 24296
rect 23440 24324 23446 24336
rect 23440 24296 23796 24324
rect 23440 24284 23446 24296
rect 22554 24216 22560 24268
rect 22612 24256 22618 24268
rect 22940 24265 23060 24266
rect 22925 24259 23060 24265
rect 22612 24228 22657 24256
rect 22612 24216 22618 24228
rect 22925 24225 22937 24259
rect 22971 24258 23060 24259
rect 22971 24256 23152 24258
rect 23198 24256 23204 24268
rect 22971 24238 23204 24256
rect 22971 24225 22983 24238
rect 23032 24230 23204 24238
rect 23124 24228 23204 24230
rect 22925 24219 22983 24225
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 22649 24191 22707 24197
rect 22649 24188 22661 24191
rect 22480 24160 22661 24188
rect 22649 24157 22661 24160
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 22741 24191 22799 24197
rect 22741 24157 22753 24191
rect 22787 24188 22799 24191
rect 22787 24160 22876 24188
rect 22787 24157 22799 24160
rect 22741 24151 22799 24157
rect 22848 24120 22876 24160
rect 23014 24148 23020 24200
rect 23072 24148 23078 24200
rect 23106 24148 23112 24200
rect 23164 24188 23170 24200
rect 23164 24160 23209 24188
rect 23164 24148 23170 24160
rect 23032 24120 23060 24148
rect 23569 24123 23627 24129
rect 23569 24120 23581 24123
rect 22848 24092 23060 24120
rect 23124 24092 23581 24120
rect 22738 24052 22744 24064
rect 21600 24024 22744 24052
rect 21600 24012 21606 24024
rect 22738 24012 22744 24024
rect 22796 24052 22802 24064
rect 23124 24052 23152 24092
rect 23569 24089 23581 24092
rect 23615 24089 23627 24123
rect 23768 24120 23796 24296
rect 24302 24284 24308 24336
rect 24360 24324 24366 24336
rect 25682 24324 25688 24336
rect 24360 24296 25688 24324
rect 24360 24284 24366 24296
rect 25682 24284 25688 24296
rect 25740 24284 25746 24336
rect 24854 24256 24860 24268
rect 24767 24228 24860 24256
rect 24854 24216 24860 24228
rect 24912 24256 24918 24268
rect 25314 24256 25320 24268
rect 24912 24228 25320 24256
rect 24912 24216 24918 24228
rect 25314 24216 25320 24228
rect 25372 24216 25378 24268
rect 25958 24216 25964 24268
rect 26016 24256 26022 24268
rect 26252 24265 26280 24364
rect 26418 24352 26424 24364
rect 26476 24352 26482 24404
rect 27062 24352 27068 24404
rect 27120 24392 27126 24404
rect 27341 24395 27399 24401
rect 27341 24392 27353 24395
rect 27120 24364 27353 24392
rect 27120 24352 27126 24364
rect 27341 24361 27353 24364
rect 27387 24361 27399 24395
rect 27341 24355 27399 24361
rect 27798 24352 27804 24404
rect 27856 24392 27862 24404
rect 28169 24395 28227 24401
rect 28169 24392 28181 24395
rect 27856 24364 28181 24392
rect 27856 24352 27862 24364
rect 28169 24361 28181 24364
rect 28215 24361 28227 24395
rect 28810 24392 28816 24404
rect 28771 24364 28816 24392
rect 28169 24355 28227 24361
rect 28810 24352 28816 24364
rect 28868 24352 28874 24404
rect 29822 24352 29828 24404
rect 29880 24392 29886 24404
rect 29917 24395 29975 24401
rect 29917 24392 29929 24395
rect 29880 24364 29929 24392
rect 29880 24352 29886 24364
rect 29917 24361 29929 24364
rect 29963 24361 29975 24395
rect 30558 24392 30564 24404
rect 30519 24364 30564 24392
rect 29917 24355 29975 24361
rect 30558 24352 30564 24364
rect 30616 24392 30622 24404
rect 30834 24392 30840 24404
rect 30616 24364 30840 24392
rect 30616 24352 30622 24364
rect 30834 24352 30840 24364
rect 30892 24352 30898 24404
rect 26326 24284 26332 24336
rect 26384 24324 26390 24336
rect 26973 24327 27031 24333
rect 26973 24324 26985 24327
rect 26384 24296 26985 24324
rect 26384 24284 26390 24296
rect 26973 24293 26985 24296
rect 27019 24293 27031 24327
rect 27154 24324 27160 24336
rect 27115 24296 27160 24324
rect 26973 24287 27031 24293
rect 27154 24284 27160 24296
rect 27212 24284 27218 24336
rect 29365 24327 29423 24333
rect 29365 24293 29377 24327
rect 29411 24324 29423 24327
rect 30282 24324 30288 24336
rect 29411 24296 30288 24324
rect 29411 24293 29423 24296
rect 29365 24287 29423 24293
rect 30282 24284 30288 24296
rect 30340 24324 30346 24336
rect 31294 24324 31300 24336
rect 30340 24296 31300 24324
rect 30340 24284 30346 24296
rect 31294 24284 31300 24296
rect 31352 24284 31358 24336
rect 26237 24259 26295 24265
rect 26237 24256 26249 24259
rect 26016 24228 26249 24256
rect 26016 24216 26022 24228
rect 26237 24225 26249 24228
rect 26283 24225 26295 24259
rect 26237 24219 26295 24225
rect 26421 24259 26479 24265
rect 26421 24225 26433 24259
rect 26467 24256 26479 24259
rect 26694 24256 26700 24268
rect 26467 24228 26700 24256
rect 26467 24225 26479 24228
rect 26421 24219 26479 24225
rect 26694 24216 26700 24228
rect 26752 24216 26758 24268
rect 28261 24259 28319 24265
rect 28261 24225 28273 24259
rect 28307 24256 28319 24259
rect 28810 24256 28816 24268
rect 28307 24228 28816 24256
rect 28307 24225 28319 24228
rect 28261 24219 28319 24225
rect 28810 24216 28816 24228
rect 28868 24216 28874 24268
rect 28905 24259 28963 24265
rect 28905 24225 28917 24259
rect 28951 24256 28963 24259
rect 29454 24256 29460 24268
rect 28951 24228 29460 24256
rect 28951 24225 28963 24228
rect 28905 24219 28963 24225
rect 29454 24216 29460 24228
rect 29512 24216 29518 24268
rect 31110 24256 31116 24268
rect 31071 24228 31116 24256
rect 31110 24216 31116 24228
rect 31168 24216 31174 24268
rect 24210 24148 24216 24200
rect 24268 24188 24274 24200
rect 24762 24188 24768 24200
rect 24268 24160 24768 24188
rect 24268 24148 24274 24160
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 25130 24148 25136 24200
rect 25188 24188 25194 24200
rect 25406 24188 25412 24200
rect 25188 24160 25412 24188
rect 25188 24148 25194 24160
rect 25406 24148 25412 24160
rect 25464 24188 25470 24200
rect 25501 24191 25559 24197
rect 25501 24188 25513 24191
rect 25464 24160 25513 24188
rect 25464 24148 25470 24160
rect 25501 24157 25513 24160
rect 25547 24157 25559 24191
rect 25501 24151 25559 24157
rect 31018 24120 31024 24132
rect 23768 24092 31024 24120
rect 23569 24083 23627 24089
rect 31018 24080 31024 24092
rect 31076 24080 31082 24132
rect 22796 24024 23152 24052
rect 22796 24012 22802 24024
rect 23198 24012 23204 24064
rect 23256 24052 23262 24064
rect 23937 24055 23995 24061
rect 23937 24052 23949 24055
rect 23256 24024 23949 24052
rect 23256 24012 23262 24024
rect 23937 24021 23949 24024
rect 23983 24021 23995 24055
rect 23937 24015 23995 24021
rect 24121 24055 24179 24061
rect 24121 24021 24133 24055
rect 24167 24052 24179 24055
rect 24578 24052 24584 24064
rect 24167 24024 24584 24052
rect 24167 24021 24179 24024
rect 24121 24015 24179 24021
rect 24578 24012 24584 24024
rect 24636 24012 24642 24064
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 26053 24055 26111 24061
rect 26053 24052 26065 24055
rect 25004 24024 26065 24052
rect 25004 24012 25010 24024
rect 26053 24021 26065 24024
rect 26099 24021 26111 24055
rect 26326 24052 26332 24064
rect 26287 24024 26332 24052
rect 26053 24015 26111 24021
rect 26326 24012 26332 24024
rect 26384 24012 26390 24064
rect 31297 24055 31355 24061
rect 31297 24021 31309 24055
rect 31343 24052 31355 24055
rect 31343 24024 32352 24052
rect 31343 24021 31355 24024
rect 31297 24015 31355 24021
rect 1104 23962 32016 23984
rect 1104 23910 6102 23962
rect 6154 23910 6166 23962
rect 6218 23910 6230 23962
rect 6282 23910 6294 23962
rect 6346 23910 6358 23962
rect 6410 23910 16405 23962
rect 16457 23910 16469 23962
rect 16521 23910 16533 23962
rect 16585 23910 16597 23962
rect 16649 23910 16661 23962
rect 16713 23910 26709 23962
rect 26761 23910 26773 23962
rect 26825 23910 26837 23962
rect 26889 23910 26901 23962
rect 26953 23910 26965 23962
rect 27017 23910 32016 23962
rect 1104 23888 32016 23910
rect 1964 23820 2774 23848
rect 1854 23644 1860 23656
rect 860 23616 1860 23644
rect 0 23508 800 23522
rect 860 23508 888 23616
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 0 23480 888 23508
rect 0 23466 800 23480
rect 1578 23468 1584 23520
rect 1636 23508 1642 23520
rect 1964 23517 1992 23820
rect 2746 23780 2774 23820
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 3789 23851 3847 23857
rect 3789 23848 3801 23851
rect 3568 23820 3801 23848
rect 3568 23808 3574 23820
rect 3789 23817 3801 23820
rect 3835 23817 3847 23851
rect 5534 23848 5540 23860
rect 3789 23811 3847 23817
rect 4264 23820 5540 23848
rect 3142 23780 3148 23792
rect 2746 23752 3148 23780
rect 3142 23740 3148 23752
rect 3200 23780 3206 23792
rect 4264 23780 4292 23820
rect 5534 23808 5540 23820
rect 5592 23808 5598 23860
rect 7834 23808 7840 23860
rect 7892 23848 7898 23860
rect 8113 23851 8171 23857
rect 8113 23848 8125 23851
rect 7892 23820 8125 23848
rect 7892 23808 7898 23820
rect 8113 23817 8125 23820
rect 8159 23817 8171 23851
rect 8113 23811 8171 23817
rect 8266 23820 12572 23848
rect 8266 23792 8294 23820
rect 3200 23752 4292 23780
rect 3200 23740 3206 23752
rect 6730 23740 6736 23792
rect 6788 23780 6794 23792
rect 6788 23752 7788 23780
rect 6788 23740 6794 23752
rect 5994 23672 6000 23724
rect 6052 23712 6058 23724
rect 6052 23684 7420 23712
rect 6052 23672 6058 23684
rect 4522 23604 4528 23656
rect 4580 23644 4586 23656
rect 4902 23647 4960 23653
rect 4902 23644 4914 23647
rect 4580 23616 4914 23644
rect 4580 23604 4586 23616
rect 4902 23613 4914 23616
rect 4948 23613 4960 23647
rect 5166 23644 5172 23656
rect 5127 23616 5172 23644
rect 4902 23607 4960 23613
rect 5166 23604 5172 23616
rect 5224 23604 5230 23656
rect 5902 23604 5908 23656
rect 5960 23644 5966 23656
rect 6089 23647 6147 23653
rect 6089 23644 6101 23647
rect 5960 23616 6101 23644
rect 5960 23604 5966 23616
rect 6089 23613 6101 23616
rect 6135 23613 6147 23647
rect 6089 23607 6147 23613
rect 6365 23647 6423 23653
rect 6365 23613 6377 23647
rect 6411 23644 6423 23647
rect 6730 23644 6736 23656
rect 6411 23616 6736 23644
rect 6411 23613 6423 23616
rect 6365 23607 6423 23613
rect 5534 23536 5540 23588
rect 5592 23576 5598 23588
rect 6380 23576 6408 23607
rect 6730 23604 6736 23616
rect 6788 23604 6794 23656
rect 7392 23653 7420 23684
rect 7466 23672 7472 23724
rect 7524 23712 7530 23724
rect 7760 23721 7788 23752
rect 8202 23740 8208 23792
rect 8260 23752 8294 23792
rect 8260 23740 8266 23752
rect 12342 23740 12348 23792
rect 12400 23780 12406 23792
rect 12437 23783 12495 23789
rect 12437 23780 12449 23783
rect 12400 23752 12449 23780
rect 12400 23740 12406 23752
rect 12437 23749 12449 23752
rect 12483 23749 12495 23783
rect 12544 23780 12572 23820
rect 12710 23808 12716 23860
rect 12768 23848 12774 23860
rect 12805 23851 12863 23857
rect 12805 23848 12817 23851
rect 12768 23820 12817 23848
rect 12768 23808 12774 23820
rect 12805 23817 12817 23820
rect 12851 23817 12863 23851
rect 12805 23811 12863 23817
rect 12989 23851 13047 23857
rect 12989 23817 13001 23851
rect 13035 23848 13047 23851
rect 13170 23848 13176 23860
rect 13035 23820 13176 23848
rect 13035 23817 13047 23820
rect 12989 23811 13047 23817
rect 13170 23808 13176 23820
rect 13228 23808 13234 23860
rect 13262 23808 13268 23860
rect 13320 23848 13326 23860
rect 13449 23851 13507 23857
rect 13449 23848 13461 23851
rect 13320 23820 13461 23848
rect 13320 23808 13326 23820
rect 13449 23817 13461 23820
rect 13495 23848 13507 23851
rect 13906 23848 13912 23860
rect 13495 23820 13912 23848
rect 13495 23817 13507 23820
rect 13449 23811 13507 23817
rect 13906 23808 13912 23820
rect 13964 23808 13970 23860
rect 16117 23851 16175 23857
rect 16117 23817 16129 23851
rect 16163 23848 16175 23851
rect 17954 23848 17960 23860
rect 16163 23820 17960 23848
rect 16163 23817 16175 23820
rect 16117 23811 16175 23817
rect 17954 23808 17960 23820
rect 18012 23808 18018 23860
rect 18693 23851 18751 23857
rect 18693 23817 18705 23851
rect 18739 23848 18751 23851
rect 19150 23848 19156 23860
rect 18739 23820 19156 23848
rect 18739 23817 18751 23820
rect 18693 23811 18751 23817
rect 19150 23808 19156 23820
rect 19208 23808 19214 23860
rect 19426 23848 19432 23860
rect 19387 23820 19432 23848
rect 19426 23808 19432 23820
rect 19484 23808 19490 23860
rect 19610 23848 19616 23860
rect 19571 23820 19616 23848
rect 19610 23808 19616 23820
rect 19668 23808 19674 23860
rect 20068 23820 22968 23848
rect 13354 23780 13360 23792
rect 12544 23752 13360 23780
rect 12437 23743 12495 23749
rect 13354 23740 13360 23752
rect 13412 23740 13418 23792
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 16298 23780 16304 23792
rect 14700 23752 16304 23780
rect 14700 23740 14706 23752
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 17037 23783 17095 23789
rect 17037 23749 17049 23783
rect 17083 23780 17095 23783
rect 20068 23780 20096 23820
rect 21542 23780 21548 23792
rect 17083 23752 20096 23780
rect 21503 23752 21548 23780
rect 17083 23749 17095 23752
rect 17037 23743 17095 23749
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7524 23684 7665 23712
rect 7524 23672 7530 23684
rect 7653 23681 7665 23684
rect 7699 23681 7711 23715
rect 7653 23675 7711 23681
rect 7745 23715 7803 23721
rect 7745 23681 7757 23715
rect 7791 23681 7803 23715
rect 7745 23675 7803 23681
rect 9030 23672 9036 23724
rect 9088 23712 9094 23724
rect 9088 23684 9444 23712
rect 9088 23672 9094 23684
rect 7377 23647 7435 23653
rect 7377 23613 7389 23647
rect 7423 23613 7435 23647
rect 7377 23607 7435 23613
rect 7561 23647 7619 23653
rect 7561 23613 7573 23647
rect 7607 23613 7619 23647
rect 7561 23607 7619 23613
rect 5592 23548 6408 23576
rect 5592 23536 5598 23548
rect 7190 23536 7196 23588
rect 7248 23576 7254 23588
rect 7576 23576 7604 23607
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 7929 23647 7987 23653
rect 7929 23644 7941 23647
rect 7892 23616 7941 23644
rect 7892 23604 7898 23616
rect 7929 23613 7941 23616
rect 7975 23613 7987 23647
rect 9214 23644 9220 23656
rect 9175 23616 9220 23644
rect 7929 23607 7987 23613
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 9416 23653 9444 23684
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 12802 23712 12808 23724
rect 12584 23684 12808 23712
rect 12584 23672 12590 23684
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 13262 23672 13268 23724
rect 13320 23712 13326 23724
rect 13814 23712 13820 23724
rect 13320 23684 13820 23712
rect 13320 23672 13326 23684
rect 13814 23672 13820 23684
rect 13872 23672 13878 23724
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23712 14887 23715
rect 15746 23712 15752 23724
rect 14875 23684 15752 23712
rect 14875 23681 14887 23684
rect 14829 23675 14887 23681
rect 15746 23672 15752 23684
rect 15804 23672 15810 23724
rect 9309 23647 9367 23653
rect 9309 23613 9321 23647
rect 9355 23613 9367 23647
rect 9309 23607 9367 23613
rect 9401 23647 9459 23653
rect 9401 23613 9413 23647
rect 9447 23613 9459 23647
rect 9401 23607 9459 23613
rect 9585 23647 9643 23653
rect 9585 23613 9597 23647
rect 9631 23644 9643 23647
rect 9858 23644 9864 23656
rect 9631 23616 9864 23644
rect 9631 23613 9643 23616
rect 9585 23607 9643 23613
rect 7248 23548 7604 23576
rect 7248 23536 7254 23548
rect 9122 23536 9128 23588
rect 9180 23576 9186 23588
rect 9324 23576 9352 23607
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 11698 23604 11704 23656
rect 11756 23653 11762 23656
rect 11756 23644 11768 23653
rect 11756 23616 11801 23644
rect 11756 23607 11768 23616
rect 11756 23604 11762 23607
rect 11882 23604 11888 23656
rect 11940 23644 11946 23656
rect 11977 23647 12035 23653
rect 11977 23644 11989 23647
rect 11940 23616 11989 23644
rect 11940 23604 11946 23616
rect 11977 23613 11989 23616
rect 12023 23613 12035 23647
rect 11977 23607 12035 23613
rect 14366 23604 14372 23656
rect 14424 23644 14430 23656
rect 14645 23647 14703 23653
rect 14645 23644 14657 23647
rect 14424 23616 14657 23644
rect 14424 23604 14430 23616
rect 14645 23613 14657 23616
rect 14691 23644 14703 23647
rect 14734 23644 14740 23656
rect 14691 23616 14740 23644
rect 14691 23613 14703 23616
rect 14645 23607 14703 23613
rect 14734 23604 14740 23616
rect 14792 23604 14798 23656
rect 14927 23647 14985 23653
rect 14927 23613 14939 23647
rect 14973 23613 14985 23647
rect 14927 23607 14985 23613
rect 15025 23647 15083 23653
rect 15025 23613 15037 23647
rect 15071 23613 15083 23647
rect 15025 23607 15083 23613
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23644 15255 23647
rect 15378 23644 15384 23656
rect 15243 23616 15384 23644
rect 15243 23613 15255 23616
rect 15197 23607 15255 23613
rect 9180 23548 9352 23576
rect 10137 23579 10195 23585
rect 9180 23536 9186 23548
rect 10137 23545 10149 23579
rect 10183 23576 10195 23579
rect 11514 23576 11520 23588
rect 10183 23548 11520 23576
rect 10183 23545 10195 23548
rect 10137 23539 10195 23545
rect 11514 23536 11520 23548
rect 11572 23576 11578 23588
rect 12342 23576 12348 23588
rect 11572 23548 12348 23576
rect 11572 23536 11578 23548
rect 12342 23536 12348 23548
rect 12400 23536 12406 23588
rect 14936 23520 14964 23607
rect 15028 23520 15056 23607
rect 15378 23604 15384 23616
rect 15436 23604 15442 23656
rect 15838 23604 15844 23656
rect 15896 23644 15902 23656
rect 15933 23647 15991 23653
rect 15933 23644 15945 23647
rect 15896 23616 15945 23644
rect 15896 23604 15902 23616
rect 15933 23613 15945 23616
rect 15979 23613 15991 23647
rect 15933 23607 15991 23613
rect 16025 23647 16083 23653
rect 16025 23613 16037 23647
rect 16071 23613 16083 23647
rect 16025 23607 16083 23613
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 16850 23644 16856 23656
rect 16255 23616 16856 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 16040 23576 16068 23607
rect 16850 23604 16856 23616
rect 16908 23604 16914 23656
rect 17126 23604 17132 23656
rect 17184 23604 17190 23656
rect 16298 23576 16304 23588
rect 16040 23548 16304 23576
rect 16298 23536 16304 23548
rect 16356 23536 16362 23588
rect 16761 23579 16819 23585
rect 16761 23545 16773 23579
rect 16807 23576 16819 23579
rect 17144 23576 17172 23604
rect 16807 23548 17172 23576
rect 16807 23545 16819 23548
rect 16761 23539 16819 23545
rect 1949 23511 2007 23517
rect 1949 23508 1961 23511
rect 1636 23480 1961 23508
rect 1636 23468 1642 23480
rect 1949 23477 1961 23480
rect 1995 23477 2007 23511
rect 1949 23471 2007 23477
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 2832 23480 2877 23508
rect 2832 23468 2838 23480
rect 2958 23468 2964 23520
rect 3016 23508 3022 23520
rect 7374 23508 7380 23520
rect 3016 23480 7380 23508
rect 3016 23468 3022 23480
rect 7374 23468 7380 23480
rect 7432 23468 7438 23520
rect 8386 23468 8392 23520
rect 8444 23508 8450 23520
rect 8941 23511 8999 23517
rect 8941 23508 8953 23511
rect 8444 23480 8953 23508
rect 8444 23468 8450 23480
rect 8941 23477 8953 23480
rect 8987 23477 8999 23511
rect 8941 23471 8999 23477
rect 10410 23468 10416 23520
rect 10468 23508 10474 23520
rect 10597 23511 10655 23517
rect 10597 23508 10609 23511
rect 10468 23480 10609 23508
rect 10468 23468 10474 23480
rect 10597 23477 10609 23480
rect 10643 23477 10655 23511
rect 10597 23471 10655 23477
rect 11974 23468 11980 23520
rect 12032 23508 12038 23520
rect 12805 23511 12863 23517
rect 12805 23508 12817 23511
rect 12032 23480 12817 23508
rect 12032 23468 12038 23480
rect 12805 23477 12817 23480
rect 12851 23477 12863 23511
rect 12805 23471 12863 23477
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 14461 23511 14519 23517
rect 14461 23508 14473 23511
rect 13872 23480 14473 23508
rect 13872 23468 13878 23480
rect 14461 23477 14473 23480
rect 14507 23477 14519 23511
rect 14461 23471 14519 23477
rect 14918 23468 14924 23520
rect 14976 23468 14982 23520
rect 15010 23468 15016 23520
rect 15068 23468 15074 23520
rect 15654 23468 15660 23520
rect 15712 23508 15718 23520
rect 17126 23508 17132 23520
rect 15712 23480 17132 23508
rect 15712 23468 15718 23480
rect 17126 23468 17132 23480
rect 17184 23508 17190 23520
rect 17236 23508 17264 23752
rect 21542 23740 21548 23752
rect 21600 23740 21606 23792
rect 22940 23780 22968 23820
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 23477 23851 23535 23857
rect 23477 23848 23489 23851
rect 23348 23820 23489 23848
rect 23348 23808 23354 23820
rect 23477 23817 23489 23820
rect 23523 23817 23535 23851
rect 23477 23811 23535 23817
rect 24486 23808 24492 23860
rect 24544 23848 24550 23860
rect 24857 23851 24915 23857
rect 24857 23848 24869 23851
rect 24544 23820 24869 23848
rect 24544 23808 24550 23820
rect 24857 23817 24869 23820
rect 24903 23817 24915 23851
rect 24857 23811 24915 23817
rect 27246 23808 27252 23860
rect 27304 23848 27310 23860
rect 27433 23851 27491 23857
rect 27433 23848 27445 23851
rect 27304 23820 27445 23848
rect 27304 23808 27310 23820
rect 27433 23817 27445 23820
rect 27479 23817 27491 23851
rect 27433 23811 27491 23817
rect 25777 23783 25835 23789
rect 22940 23752 24992 23780
rect 19981 23715 20039 23721
rect 19981 23712 19993 23715
rect 17972 23684 19993 23712
rect 17972 23653 18000 23684
rect 19981 23681 19993 23684
rect 20027 23712 20039 23715
rect 20438 23712 20444 23724
rect 20027 23684 20444 23712
rect 20027 23681 20039 23684
rect 19981 23675 20039 23681
rect 20438 23672 20444 23684
rect 20496 23712 20502 23724
rect 20990 23712 20996 23724
rect 20496 23684 20996 23712
rect 20496 23672 20502 23684
rect 20990 23672 20996 23684
rect 21048 23672 21054 23724
rect 17957 23647 18015 23653
rect 17957 23613 17969 23647
rect 18003 23613 18015 23647
rect 18138 23644 18144 23656
rect 18099 23616 18144 23644
rect 17957 23607 18015 23613
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 18233 23647 18291 23653
rect 18233 23613 18245 23647
rect 18279 23613 18291 23647
rect 18233 23607 18291 23613
rect 18325 23647 18383 23653
rect 18325 23613 18337 23647
rect 18371 23613 18383 23647
rect 18325 23607 18383 23613
rect 18509 23647 18567 23653
rect 18509 23613 18521 23647
rect 18555 23644 18567 23647
rect 19610 23644 19616 23656
rect 18555 23616 19616 23644
rect 18555 23613 18567 23616
rect 18509 23607 18567 23613
rect 17586 23536 17592 23588
rect 17644 23576 17650 23588
rect 18248 23576 18276 23607
rect 17644 23548 18276 23576
rect 17644 23536 17650 23548
rect 17184 23480 17264 23508
rect 17184 23468 17190 23480
rect 17678 23468 17684 23520
rect 17736 23508 17742 23520
rect 18340 23508 18368 23607
rect 19610 23604 19616 23616
rect 19668 23604 19674 23656
rect 20622 23604 20628 23656
rect 20680 23644 20686 23656
rect 20717 23647 20775 23653
rect 20717 23644 20729 23647
rect 20680 23616 20729 23644
rect 20680 23604 20686 23616
rect 20717 23613 20729 23616
rect 20763 23613 20775 23647
rect 20717 23607 20775 23613
rect 20806 23604 20812 23656
rect 20864 23644 20870 23656
rect 21560 23644 21588 23740
rect 23106 23672 23112 23724
rect 23164 23712 23170 23724
rect 24397 23715 24455 23721
rect 24397 23712 24409 23715
rect 23164 23684 24409 23712
rect 23164 23672 23170 23684
rect 24397 23681 24409 23684
rect 24443 23681 24455 23715
rect 24397 23675 24455 23681
rect 20864 23616 21588 23644
rect 20864 23604 20870 23616
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22925 23647 22983 23653
rect 22925 23644 22937 23647
rect 22152 23616 22937 23644
rect 22152 23604 22158 23616
rect 22925 23613 22937 23616
rect 22971 23613 22983 23647
rect 22925 23607 22983 23613
rect 23569 23647 23627 23653
rect 23569 23613 23581 23647
rect 23615 23613 23627 23647
rect 24578 23644 24584 23656
rect 24539 23616 24584 23644
rect 23569 23607 23627 23613
rect 20070 23536 20076 23588
rect 20128 23576 20134 23588
rect 20533 23579 20591 23585
rect 20533 23576 20545 23579
rect 20128 23548 20545 23576
rect 20128 23536 20134 23548
rect 20533 23545 20545 23548
rect 20579 23545 20591 23579
rect 22462 23576 22468 23588
rect 20533 23539 20591 23545
rect 20640 23548 22468 23576
rect 17736 23480 18368 23508
rect 17736 23468 17742 23480
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19613 23511 19671 23517
rect 19613 23508 19625 23511
rect 19392 23480 19625 23508
rect 19392 23468 19398 23480
rect 19613 23477 19625 23480
rect 19659 23508 19671 23511
rect 20640 23508 20668 23548
rect 22462 23536 22468 23548
rect 22520 23536 22526 23588
rect 22554 23536 22560 23588
rect 22612 23576 22618 23588
rect 22658 23579 22716 23585
rect 22658 23576 22670 23579
rect 22612 23548 22670 23576
rect 22612 23536 22618 23548
rect 22658 23545 22670 23548
rect 22704 23545 22716 23579
rect 22658 23539 22716 23545
rect 23106 23536 23112 23588
rect 23164 23576 23170 23588
rect 23584 23576 23612 23607
rect 24578 23604 24584 23616
rect 24636 23604 24642 23656
rect 24964 23653 24992 23752
rect 25777 23749 25789 23783
rect 25823 23780 25835 23783
rect 27062 23780 27068 23792
rect 25823 23752 27068 23780
rect 25823 23749 25835 23752
rect 25777 23743 25835 23749
rect 27062 23740 27068 23752
rect 27120 23780 27126 23792
rect 27338 23780 27344 23792
rect 27120 23752 27344 23780
rect 27120 23740 27126 23752
rect 27338 23740 27344 23752
rect 27396 23740 27402 23792
rect 28994 23712 29000 23724
rect 28368 23684 29000 23712
rect 24949 23647 25007 23653
rect 24949 23613 24961 23647
rect 24995 23644 25007 23647
rect 25038 23644 25044 23656
rect 24995 23616 25044 23644
rect 24995 23613 25007 23616
rect 24949 23607 25007 23613
rect 25038 23604 25044 23616
rect 25096 23604 25102 23656
rect 26237 23647 26295 23653
rect 26237 23644 26249 23647
rect 25424 23616 26249 23644
rect 23164 23548 23612 23576
rect 23164 23536 23170 23548
rect 25314 23536 25320 23588
rect 25372 23576 25378 23588
rect 25424 23585 25452 23616
rect 26237 23613 26249 23616
rect 26283 23613 26295 23647
rect 26237 23607 26295 23613
rect 26421 23647 26479 23653
rect 26421 23613 26433 23647
rect 26467 23644 26479 23647
rect 28166 23644 28172 23656
rect 26467 23616 27200 23644
rect 28127 23616 28172 23644
rect 26467 23613 26479 23616
rect 26421 23607 26479 23613
rect 27172 23588 27200 23616
rect 28166 23604 28172 23616
rect 28224 23604 28230 23656
rect 28368 23653 28396 23684
rect 28994 23672 29000 23684
rect 29052 23672 29058 23724
rect 28353 23647 28411 23653
rect 28353 23613 28365 23647
rect 28399 23613 28411 23647
rect 28353 23607 28411 23613
rect 28448 23647 28506 23653
rect 28448 23613 28460 23647
rect 28494 23613 28506 23647
rect 28448 23607 28506 23613
rect 25409 23579 25467 23585
rect 25409 23576 25421 23579
rect 25372 23548 25421 23576
rect 25372 23536 25378 23548
rect 25409 23545 25421 23548
rect 25455 23545 25467 23579
rect 25409 23539 25467 23545
rect 25593 23579 25651 23585
rect 25593 23545 25605 23579
rect 25639 23545 25651 23579
rect 25593 23539 25651 23545
rect 19659 23480 20668 23508
rect 19659 23477 19671 23480
rect 19613 23471 19671 23477
rect 22278 23468 22284 23520
rect 22336 23508 22342 23520
rect 25608 23508 25636 23539
rect 26050 23536 26056 23588
rect 26108 23576 26114 23588
rect 27065 23579 27123 23585
rect 27065 23576 27077 23579
rect 26108 23548 27077 23576
rect 26108 23536 26114 23548
rect 27065 23545 27077 23548
rect 27111 23545 27123 23579
rect 27065 23539 27123 23545
rect 27154 23536 27160 23588
rect 27212 23576 27218 23588
rect 27249 23579 27307 23585
rect 27249 23576 27261 23579
rect 27212 23548 27261 23576
rect 27212 23536 27218 23548
rect 27249 23545 27261 23548
rect 27295 23545 27307 23579
rect 27249 23539 27307 23545
rect 28460 23520 28488 23607
rect 28534 23604 28540 23656
rect 28592 23644 28598 23656
rect 28721 23647 28779 23653
rect 28592 23616 28637 23644
rect 28592 23604 28598 23616
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 28810 23644 28816 23656
rect 28767 23616 28816 23644
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 28810 23604 28816 23616
rect 28868 23604 28874 23656
rect 30926 23644 30932 23656
rect 30887 23616 30932 23644
rect 30926 23604 30932 23616
rect 30984 23604 30990 23656
rect 32324 23644 32352 24024
rect 32232 23616 32352 23644
rect 28905 23579 28963 23585
rect 28905 23545 28917 23579
rect 28951 23576 28963 23579
rect 30662 23579 30720 23585
rect 30662 23576 30674 23579
rect 28951 23548 30674 23576
rect 28951 23545 28963 23548
rect 28905 23539 28963 23545
rect 30662 23545 30674 23548
rect 30708 23545 30720 23579
rect 30662 23539 30720 23545
rect 26326 23508 26332 23520
rect 22336 23480 26332 23508
rect 22336 23468 22342 23480
rect 26326 23468 26332 23480
rect 26384 23468 26390 23520
rect 26605 23511 26663 23517
rect 26605 23477 26617 23511
rect 26651 23508 26663 23511
rect 26694 23508 26700 23520
rect 26651 23480 26700 23508
rect 26651 23477 26663 23480
rect 26605 23471 26663 23477
rect 26694 23468 26700 23480
rect 26752 23468 26758 23520
rect 28442 23468 28448 23520
rect 28500 23468 28506 23520
rect 28810 23468 28816 23520
rect 28868 23508 28874 23520
rect 29549 23511 29607 23517
rect 29549 23508 29561 23511
rect 28868 23480 29561 23508
rect 28868 23468 28874 23480
rect 29549 23477 29561 23480
rect 29595 23477 29607 23511
rect 32232 23508 32260 23616
rect 32320 23508 33120 23522
rect 32232 23480 33120 23508
rect 29549 23471 29607 23477
rect 32320 23466 33120 23480
rect 1104 23418 32016 23440
rect 1104 23366 11253 23418
rect 11305 23366 11317 23418
rect 11369 23366 11381 23418
rect 11433 23366 11445 23418
rect 11497 23366 11509 23418
rect 11561 23366 21557 23418
rect 21609 23366 21621 23418
rect 21673 23366 21685 23418
rect 21737 23366 21749 23418
rect 21801 23366 21813 23418
rect 21865 23366 32016 23418
rect 1104 23344 32016 23366
rect 2222 23264 2228 23316
rect 2280 23304 2286 23316
rect 2406 23304 2412 23316
rect 2280 23276 2412 23304
rect 2280 23264 2286 23276
rect 2406 23264 2412 23276
rect 2464 23304 2470 23316
rect 3237 23307 3295 23313
rect 3237 23304 3249 23307
rect 2464 23276 3249 23304
rect 2464 23264 2470 23276
rect 3237 23273 3249 23276
rect 3283 23273 3295 23307
rect 3237 23267 3295 23273
rect 3881 23307 3939 23313
rect 3881 23273 3893 23307
rect 3927 23304 3939 23307
rect 4430 23304 4436 23316
rect 3927 23276 4436 23304
rect 3927 23273 3939 23276
rect 3881 23267 3939 23273
rect 4430 23264 4436 23276
rect 4488 23264 4494 23316
rect 6822 23264 6828 23316
rect 6880 23304 6886 23316
rect 7466 23304 7472 23316
rect 6880 23276 7472 23304
rect 6880 23264 6886 23276
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 7653 23307 7711 23313
rect 7653 23273 7665 23307
rect 7699 23304 7711 23307
rect 8018 23304 8024 23316
rect 7699 23276 8024 23304
rect 7699 23273 7711 23276
rect 7653 23267 7711 23273
rect 8018 23264 8024 23276
rect 8076 23264 8082 23316
rect 12986 23264 12992 23316
rect 13044 23304 13050 23316
rect 16942 23304 16948 23316
rect 13044 23276 16948 23304
rect 13044 23264 13050 23276
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 18230 23264 18236 23316
rect 18288 23304 18294 23316
rect 18874 23304 18880 23316
rect 18288 23276 18880 23304
rect 18288 23264 18294 23276
rect 18874 23264 18880 23276
rect 18932 23264 18938 23316
rect 19978 23304 19984 23316
rect 19939 23276 19984 23304
rect 19978 23264 19984 23276
rect 20036 23304 20042 23316
rect 20036 23276 20852 23304
rect 20036 23264 20042 23276
rect 5166 23236 5172 23248
rect 1872 23208 5172 23236
rect 1394 23060 1400 23112
rect 1452 23100 1458 23112
rect 1872 23109 1900 23208
rect 2124 23171 2182 23177
rect 2124 23137 2136 23171
rect 2170 23168 2182 23171
rect 2590 23168 2596 23180
rect 2170 23140 2596 23168
rect 2170 23137 2182 23140
rect 2124 23131 2182 23137
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 4356 23177 4384 23208
rect 5166 23196 5172 23208
rect 5224 23196 5230 23248
rect 7006 23236 7012 23248
rect 6564 23208 7012 23236
rect 4341 23171 4399 23177
rect 4341 23137 4353 23171
rect 4387 23137 4399 23171
rect 4597 23171 4655 23177
rect 4597 23168 4609 23171
rect 4341 23131 4399 23137
rect 4448 23140 4609 23168
rect 1857 23103 1915 23109
rect 1857 23100 1869 23103
rect 1452 23072 1869 23100
rect 1452 23060 1458 23072
rect 1857 23069 1869 23072
rect 1903 23069 1915 23103
rect 1857 23063 1915 23069
rect 3234 23060 3240 23112
rect 3292 23100 3298 23112
rect 4448 23100 4476 23140
rect 4597 23137 4609 23140
rect 4643 23137 4655 23171
rect 4597 23131 4655 23137
rect 5994 23128 6000 23180
rect 6052 23168 6058 23180
rect 6564 23177 6592 23208
rect 7006 23196 7012 23208
rect 7064 23236 7070 23248
rect 7834 23236 7840 23248
rect 7064 23208 7840 23236
rect 7064 23196 7070 23208
rect 7834 23196 7840 23208
rect 7892 23196 7898 23248
rect 8938 23196 8944 23248
rect 8996 23236 9002 23248
rect 17589 23239 17647 23245
rect 17589 23236 17601 23239
rect 8996 23208 17601 23236
rect 8996 23196 9002 23208
rect 17589 23205 17601 23208
rect 17635 23205 17647 23239
rect 17589 23199 17647 23205
rect 20438 23196 20444 23248
rect 20496 23236 20502 23248
rect 20496 23208 20760 23236
rect 20496 23196 20502 23208
rect 6365 23171 6423 23177
rect 6365 23168 6377 23171
rect 6052 23140 6377 23168
rect 6052 23128 6058 23140
rect 6365 23137 6377 23140
rect 6411 23137 6423 23171
rect 6365 23131 6423 23137
rect 6549 23171 6607 23177
rect 6549 23137 6561 23171
rect 6595 23137 6607 23171
rect 6730 23168 6736 23180
rect 6691 23140 6736 23168
rect 6549 23131 6607 23137
rect 6730 23128 6736 23140
rect 6788 23128 6794 23180
rect 6914 23168 6920 23180
rect 6875 23140 6920 23168
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 7466 23128 7472 23180
rect 7524 23168 7530 23180
rect 7745 23171 7803 23177
rect 7745 23168 7757 23171
rect 7524 23140 7757 23168
rect 7524 23128 7530 23140
rect 7745 23137 7757 23140
rect 7791 23137 7803 23171
rect 7745 23131 7803 23137
rect 8297 23171 8355 23177
rect 8297 23137 8309 23171
rect 8343 23168 8355 23171
rect 8478 23168 8484 23180
rect 8343 23140 8484 23168
rect 8343 23137 8355 23140
rect 8297 23131 8355 23137
rect 8478 23128 8484 23140
rect 8536 23128 8542 23180
rect 9306 23168 9312 23180
rect 9267 23140 9312 23168
rect 9306 23128 9312 23140
rect 9364 23128 9370 23180
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 9953 23171 10011 23177
rect 9953 23168 9965 23171
rect 9548 23140 9965 23168
rect 9548 23128 9554 23140
rect 9953 23137 9965 23140
rect 9999 23137 10011 23171
rect 9953 23131 10011 23137
rect 10042 23128 10048 23180
rect 10100 23168 10106 23180
rect 11517 23171 11575 23177
rect 11517 23168 11529 23171
rect 10100 23140 11529 23168
rect 10100 23128 10106 23140
rect 11517 23137 11529 23140
rect 11563 23137 11575 23171
rect 11517 23131 11575 23137
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 12621 23171 12679 23177
rect 12621 23168 12633 23171
rect 12492 23140 12633 23168
rect 12492 23128 12498 23140
rect 12621 23137 12633 23140
rect 12667 23137 12679 23171
rect 12621 23131 12679 23137
rect 12897 23171 12955 23177
rect 12897 23137 12909 23171
rect 12943 23168 12955 23171
rect 12986 23168 12992 23180
rect 12943 23140 12992 23168
rect 12943 23137 12955 23140
rect 12897 23131 12955 23137
rect 6641 23103 6699 23109
rect 6641 23100 6653 23103
rect 3292 23072 4476 23100
rect 6564 23072 6653 23100
rect 3292 23060 3298 23072
rect 6564 23044 6592 23072
rect 6641 23069 6653 23072
rect 6687 23069 6699 23103
rect 6641 23063 6699 23069
rect 8110 23060 8116 23112
rect 8168 23100 8174 23112
rect 8389 23103 8447 23109
rect 8389 23100 8401 23103
rect 8168 23072 8401 23100
rect 8168 23060 8174 23072
rect 8389 23069 8401 23072
rect 8435 23069 8447 23103
rect 8570 23100 8576 23112
rect 8531 23072 8576 23100
rect 8389 23063 8447 23069
rect 5902 23032 5908 23044
rect 5276 23004 5908 23032
rect 4246 22924 4252 22976
rect 4304 22964 4310 22976
rect 5276 22964 5304 23004
rect 5902 22992 5908 23004
rect 5960 22992 5966 23044
rect 6546 22992 6552 23044
rect 6604 22992 6610 23044
rect 5718 22964 5724 22976
rect 4304 22936 5304 22964
rect 5679 22936 5724 22964
rect 4304 22924 4310 22936
rect 5718 22924 5724 22936
rect 5776 22924 5782 22976
rect 6822 22924 6828 22976
rect 6880 22964 6886 22976
rect 7101 22967 7159 22973
rect 7101 22964 7113 22967
rect 6880 22936 7113 22964
rect 6880 22924 6886 22936
rect 7101 22933 7113 22936
rect 7147 22933 7159 22967
rect 8404 22964 8432 23063
rect 8570 23060 8576 23072
rect 8628 23060 8634 23112
rect 9585 23103 9643 23109
rect 9585 23100 9597 23103
rect 8956 23072 9597 23100
rect 8481 23035 8539 23041
rect 8481 23001 8493 23035
rect 8527 23032 8539 23035
rect 8956 23032 8984 23072
rect 9585 23069 9597 23072
rect 9631 23069 9643 23103
rect 9585 23063 9643 23069
rect 10321 23103 10379 23109
rect 10321 23069 10333 23103
rect 10367 23100 10379 23103
rect 11609 23103 11667 23109
rect 11609 23100 11621 23103
rect 10367 23072 11621 23100
rect 10367 23069 10379 23072
rect 10321 23063 10379 23069
rect 11609 23069 11621 23072
rect 11655 23069 11667 23103
rect 11609 23063 11667 23069
rect 8527 23004 8984 23032
rect 9769 23035 9827 23041
rect 8527 23001 8539 23004
rect 8481 22995 8539 23001
rect 9769 23001 9781 23035
rect 9815 23032 9827 23035
rect 10502 23032 10508 23044
rect 9815 23004 10508 23032
rect 9815 23001 9827 23004
rect 9769 22995 9827 23001
rect 10502 22992 10508 23004
rect 10560 22992 10566 23044
rect 8570 22964 8576 22976
rect 8404 22936 8576 22964
rect 7101 22927 7159 22933
rect 8570 22924 8576 22936
rect 8628 22924 8634 22976
rect 12636 22964 12664 23131
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 13538 23168 13544 23180
rect 13499 23140 13544 23168
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 13814 23177 13820 23180
rect 13808 23168 13820 23177
rect 13775 23140 13820 23168
rect 13808 23131 13820 23140
rect 13814 23128 13820 23131
rect 13872 23128 13878 23180
rect 14366 23128 14372 23180
rect 14424 23168 14430 23180
rect 15378 23168 15384 23180
rect 14424 23140 15240 23168
rect 15339 23140 15384 23168
rect 14424 23128 14430 23140
rect 15212 23100 15240 23140
rect 15378 23128 15384 23140
rect 15436 23128 15442 23180
rect 15562 23168 15568 23180
rect 15475 23140 15568 23168
rect 15562 23128 15568 23140
rect 15620 23128 15626 23180
rect 15746 23168 15752 23180
rect 15707 23140 15752 23168
rect 15746 23128 15752 23140
rect 15804 23128 15810 23180
rect 15838 23128 15844 23180
rect 15896 23168 15902 23180
rect 15933 23171 15991 23177
rect 15933 23168 15945 23171
rect 15896 23140 15945 23168
rect 15896 23128 15902 23140
rect 15933 23137 15945 23140
rect 15979 23137 15991 23171
rect 15933 23131 15991 23137
rect 16022 23128 16028 23180
rect 16080 23168 16086 23180
rect 17037 23171 17095 23177
rect 17037 23168 17049 23171
rect 16080 23140 17049 23168
rect 16080 23128 16086 23140
rect 17037 23137 17049 23140
rect 17083 23168 17095 23171
rect 19889 23171 19947 23177
rect 19889 23168 19901 23171
rect 17083 23140 19901 23168
rect 17083 23137 17095 23140
rect 17037 23131 17095 23137
rect 19889 23137 19901 23140
rect 19935 23137 19947 23171
rect 19889 23131 19947 23137
rect 20533 23171 20591 23177
rect 20533 23137 20545 23171
rect 20579 23168 20591 23171
rect 20622 23168 20628 23180
rect 20579 23140 20628 23168
rect 20579 23137 20591 23140
rect 20533 23131 20591 23137
rect 15580 23100 15608 23128
rect 15212 23072 15608 23100
rect 15657 23103 15715 23109
rect 15657 23069 15669 23103
rect 15703 23100 15715 23103
rect 15703 23072 16988 23100
rect 15703 23069 15715 23072
rect 15657 23063 15715 23069
rect 14182 22964 14188 22976
rect 12636 22936 14188 22964
rect 14182 22924 14188 22936
rect 14240 22924 14246 22976
rect 14734 22924 14740 22976
rect 14792 22964 14798 22976
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 14792 22936 14933 22964
rect 14792 22924 14798 22936
rect 14921 22933 14933 22936
rect 14967 22964 14979 22967
rect 15102 22964 15108 22976
rect 14967 22936 15108 22964
rect 14967 22933 14979 22936
rect 14921 22927 14979 22933
rect 15102 22924 15108 22936
rect 15160 22924 15166 22976
rect 16022 22924 16028 22976
rect 16080 22964 16086 22976
rect 16960 22973 16988 23072
rect 18046 23060 18052 23112
rect 18104 23100 18110 23112
rect 18506 23100 18512 23112
rect 18104 23072 18512 23100
rect 18104 23060 18110 23072
rect 18506 23060 18512 23072
rect 18564 23060 18570 23112
rect 16117 22967 16175 22973
rect 16117 22964 16129 22967
rect 16080 22936 16129 22964
rect 16080 22924 16086 22936
rect 16117 22933 16129 22936
rect 16163 22933 16175 22967
rect 16117 22927 16175 22933
rect 16945 22967 17003 22973
rect 16945 22933 16957 22967
rect 16991 22964 17003 22967
rect 18598 22964 18604 22976
rect 16991 22936 18604 22964
rect 16991 22933 17003 22936
rect 16945 22927 17003 22933
rect 18598 22924 18604 22936
rect 18656 22924 18662 22976
rect 19904 22964 19932 23131
rect 20548 23032 20576 23131
rect 20622 23128 20628 23140
rect 20680 23128 20686 23180
rect 20732 23177 20760 23208
rect 20824 23177 20852 23276
rect 20898 23264 20904 23316
rect 20956 23304 20962 23316
rect 22554 23304 22560 23316
rect 20956 23276 22324 23304
rect 22515 23276 22560 23304
rect 20956 23264 20962 23276
rect 20916 23177 20944 23264
rect 21100 23208 22048 23236
rect 21100 23177 21128 23208
rect 22020 23180 22048 23208
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23137 20775 23171
rect 20717 23131 20775 23137
rect 20809 23171 20867 23177
rect 20809 23137 20821 23171
rect 20855 23137 20867 23171
rect 20809 23131 20867 23137
rect 20901 23171 20959 23177
rect 20901 23137 20913 23171
rect 20947 23137 20959 23171
rect 20901 23131 20959 23137
rect 21085 23171 21143 23177
rect 21085 23137 21097 23171
rect 21131 23137 21143 23171
rect 21266 23168 21272 23180
rect 21227 23140 21272 23168
rect 21085 23131 21143 23137
rect 20824 23100 20852 23131
rect 21266 23128 21272 23140
rect 21324 23128 21330 23180
rect 21818 23168 21824 23180
rect 21779 23140 21824 23168
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 22002 23128 22008 23180
rect 22060 23168 22066 23180
rect 22189 23171 22247 23177
rect 22060 23140 22153 23168
rect 22060 23128 22066 23140
rect 22189 23137 22201 23171
rect 22235 23168 22247 23171
rect 22296 23168 22324 23276
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 24946 23304 24952 23316
rect 24859 23276 24952 23304
rect 24946 23264 24952 23276
rect 25004 23304 25010 23316
rect 25222 23304 25228 23316
rect 25004 23276 25228 23304
rect 25004 23264 25010 23276
rect 25222 23264 25228 23276
rect 25280 23264 25286 23316
rect 26421 23307 26479 23313
rect 26421 23273 26433 23307
rect 26467 23304 26479 23307
rect 26510 23304 26516 23316
rect 26467 23276 26516 23304
rect 26467 23273 26479 23276
rect 26421 23267 26479 23273
rect 26510 23264 26516 23276
rect 26568 23264 26574 23316
rect 30282 23304 30288 23316
rect 26620 23276 29776 23304
rect 30243 23276 30288 23304
rect 24486 23196 24492 23248
rect 24544 23236 24550 23248
rect 26620 23236 26648 23276
rect 29748 23245 29776 23276
rect 30282 23264 30288 23276
rect 30340 23264 30346 23316
rect 31110 23264 31116 23316
rect 31168 23304 31174 23316
rect 31297 23307 31355 23313
rect 31297 23304 31309 23307
rect 31168 23276 31309 23304
rect 31168 23264 31174 23276
rect 31297 23273 31309 23276
rect 31343 23273 31355 23307
rect 31297 23267 31355 23273
rect 29089 23239 29147 23245
rect 29089 23236 29101 23239
rect 24544 23208 26648 23236
rect 27540 23208 29101 23236
rect 24544 23196 24550 23208
rect 22235 23140 22324 23168
rect 22373 23171 22431 23177
rect 22235 23137 22247 23140
rect 22189 23131 22247 23137
rect 22373 23137 22385 23171
rect 22419 23168 22431 23171
rect 22738 23168 22744 23180
rect 22419 23140 22744 23168
rect 22419 23137 22431 23140
rect 22373 23131 22431 23137
rect 22738 23128 22744 23140
rect 22796 23128 22802 23180
rect 23836 23171 23894 23177
rect 23836 23137 23848 23171
rect 23882 23168 23894 23171
rect 24394 23168 24400 23180
rect 23882 23140 24400 23168
rect 23882 23137 23894 23140
rect 23836 23131 23894 23137
rect 24394 23128 24400 23140
rect 24452 23128 24458 23180
rect 25774 23128 25780 23180
rect 25832 23168 25838 23180
rect 27540 23177 27568 23208
rect 29089 23205 29101 23208
rect 29135 23205 29147 23239
rect 29089 23199 29147 23205
rect 29733 23239 29791 23245
rect 29733 23205 29745 23239
rect 29779 23236 29791 23239
rect 30190 23236 30196 23248
rect 29779 23208 30196 23236
rect 29779 23205 29791 23208
rect 29733 23199 29791 23205
rect 30190 23196 30196 23208
rect 30248 23196 30254 23248
rect 25869 23171 25927 23177
rect 25869 23168 25881 23171
rect 25832 23140 25881 23168
rect 25832 23128 25838 23140
rect 25869 23137 25881 23140
rect 25915 23137 25927 23171
rect 25869 23131 25927 23137
rect 27525 23171 27583 23177
rect 27525 23137 27537 23171
rect 27571 23137 27583 23171
rect 27525 23131 27583 23137
rect 27617 23171 27675 23177
rect 27617 23137 27629 23171
rect 27663 23137 27675 23171
rect 27617 23131 27675 23137
rect 27893 23171 27951 23177
rect 27893 23137 27905 23171
rect 27939 23168 27951 23171
rect 28445 23171 28503 23177
rect 28445 23168 28457 23171
rect 27939 23140 28457 23168
rect 27939 23137 27951 23140
rect 27893 23131 27951 23137
rect 28445 23137 28457 23140
rect 28491 23137 28503 23171
rect 28445 23131 28503 23137
rect 28537 23171 28595 23177
rect 28537 23137 28549 23171
rect 28583 23137 28595 23171
rect 28537 23131 28595 23137
rect 22097 23103 22155 23109
rect 22097 23100 22109 23103
rect 20824 23072 22109 23100
rect 22097 23069 22109 23072
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 23290 23060 23296 23112
rect 23348 23100 23354 23112
rect 23569 23103 23627 23109
rect 23569 23100 23581 23103
rect 23348 23072 23581 23100
rect 23348 23060 23354 23072
rect 23569 23069 23581 23072
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 26145 23103 26203 23109
rect 26145 23069 26157 23103
rect 26191 23100 26203 23103
rect 27154 23100 27160 23112
rect 26191 23072 27160 23100
rect 26191 23069 26203 23072
rect 26145 23063 26203 23069
rect 27154 23060 27160 23072
rect 27212 23060 27218 23112
rect 27246 23060 27252 23112
rect 27304 23100 27310 23112
rect 27632 23100 27660 23131
rect 27304 23072 27660 23100
rect 28552 23100 28580 23131
rect 28626 23128 28632 23180
rect 28684 23168 28690 23180
rect 28997 23171 29055 23177
rect 28997 23168 29009 23171
rect 28684 23140 29009 23168
rect 28684 23128 28690 23140
rect 28997 23137 29009 23140
rect 29043 23137 29055 23171
rect 28997 23131 29055 23137
rect 31018 23128 31024 23180
rect 31076 23168 31082 23180
rect 31113 23171 31171 23177
rect 31113 23168 31125 23171
rect 31076 23140 31125 23168
rect 31076 23128 31082 23140
rect 31113 23137 31125 23140
rect 31159 23168 31171 23171
rect 31294 23168 31300 23180
rect 31159 23140 31300 23168
rect 31159 23137 31171 23140
rect 31113 23131 31171 23137
rect 31294 23128 31300 23140
rect 31352 23128 31358 23180
rect 28718 23100 28724 23112
rect 28552 23072 28724 23100
rect 27304 23060 27310 23072
rect 28718 23060 28724 23072
rect 28776 23060 28782 23112
rect 21818 23032 21824 23044
rect 20548 23004 21824 23032
rect 21818 22992 21824 23004
rect 21876 22992 21882 23044
rect 22002 22992 22008 23044
rect 22060 23032 22066 23044
rect 23106 23032 23112 23044
rect 22060 23004 23112 23032
rect 22060 22992 22066 23004
rect 23106 22992 23112 23004
rect 23164 22992 23170 23044
rect 26694 22992 26700 23044
rect 26752 23032 26758 23044
rect 27430 23032 27436 23044
rect 26752 23004 27436 23032
rect 26752 22992 26758 23004
rect 27430 22992 27436 23004
rect 27488 23032 27494 23044
rect 27801 23035 27859 23041
rect 27801 23032 27813 23035
rect 27488 23004 27813 23032
rect 27488 22992 27494 23004
rect 27801 23001 27813 23004
rect 27847 23001 27859 23035
rect 27801 22995 27859 23001
rect 20898 22964 20904 22976
rect 19904 22936 20904 22964
rect 20898 22924 20904 22936
rect 20956 22964 20962 22976
rect 23017 22967 23075 22973
rect 23017 22964 23029 22967
rect 20956 22936 23029 22964
rect 20956 22924 20962 22936
rect 23017 22933 23029 22936
rect 23063 22933 23075 22967
rect 26050 22964 26056 22976
rect 26011 22936 26056 22964
rect 23017 22927 23075 22933
rect 26050 22924 26056 22936
rect 26108 22924 26114 22976
rect 27246 22924 27252 22976
rect 27304 22964 27310 22976
rect 27341 22967 27399 22973
rect 27341 22964 27353 22967
rect 27304 22936 27353 22964
rect 27304 22924 27310 22936
rect 27341 22933 27353 22936
rect 27387 22933 27399 22967
rect 27341 22927 27399 22933
rect 1104 22874 32016 22896
rect 1104 22822 6102 22874
rect 6154 22822 6166 22874
rect 6218 22822 6230 22874
rect 6282 22822 6294 22874
rect 6346 22822 6358 22874
rect 6410 22822 16405 22874
rect 16457 22822 16469 22874
rect 16521 22822 16533 22874
rect 16585 22822 16597 22874
rect 16649 22822 16661 22874
rect 16713 22822 26709 22874
rect 26761 22822 26773 22874
rect 26825 22822 26837 22874
rect 26889 22822 26901 22874
rect 26953 22822 26965 22874
rect 27017 22822 32016 22874
rect 1104 22800 32016 22822
rect 1946 22720 1952 22772
rect 2004 22760 2010 22772
rect 2590 22760 2596 22772
rect 2004 22732 2268 22760
rect 2551 22732 2596 22760
rect 2004 22720 2010 22732
rect 2240 22633 2268 22732
rect 2590 22720 2596 22732
rect 2648 22720 2654 22772
rect 5166 22720 5172 22772
rect 5224 22760 5230 22772
rect 5902 22760 5908 22772
rect 5224 22732 5908 22760
rect 5224 22720 5230 22732
rect 5902 22720 5908 22732
rect 5960 22720 5966 22772
rect 8297 22763 8355 22769
rect 8297 22729 8309 22763
rect 8343 22760 8355 22763
rect 9306 22760 9312 22772
rect 8343 22732 9312 22760
rect 8343 22729 8355 22732
rect 8297 22723 8355 22729
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 10042 22760 10048 22772
rect 10003 22732 10048 22760
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 10870 22760 10876 22772
rect 10796 22732 10876 22760
rect 5626 22652 5632 22704
rect 5684 22692 5690 22704
rect 6730 22692 6736 22704
rect 5684 22664 6736 22692
rect 5684 22652 5690 22664
rect 6730 22652 6736 22664
rect 6788 22692 6794 22704
rect 8478 22692 8484 22704
rect 6788 22664 7236 22692
rect 6788 22652 6794 22664
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22593 2283 22627
rect 2225 22587 2283 22593
rect 6270 22584 6276 22636
rect 6328 22624 6334 22636
rect 6546 22624 6552 22636
rect 6328 22596 6552 22624
rect 6328 22584 6334 22596
rect 6546 22584 6552 22596
rect 6604 22624 6610 22636
rect 7208 22633 7236 22664
rect 8128 22664 8484 22692
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 6604 22596 7113 22624
rect 6604 22584 6610 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 7558 22584 7564 22636
rect 7616 22624 7622 22636
rect 7616 22596 7880 22624
rect 7616 22584 7622 22596
rect 2038 22556 2044 22568
rect 2096 22565 2102 22568
rect 1845 22549 1903 22555
rect 1845 22546 1857 22549
rect 1780 22518 1857 22546
rect 1780 22420 1808 22518
rect 1845 22515 1857 22518
rect 1891 22515 1903 22549
rect 2003 22528 2044 22556
rect 2038 22516 2044 22528
rect 2096 22519 2103 22565
rect 2096 22516 2102 22519
rect 2133 22516 2139 22568
rect 2191 22565 2197 22568
rect 2191 22556 2200 22565
rect 2406 22556 2412 22568
rect 2191 22528 2236 22556
rect 2367 22528 2412 22556
rect 2191 22519 2200 22528
rect 2191 22516 2197 22519
rect 2406 22516 2412 22528
rect 2464 22516 2470 22568
rect 3973 22559 4031 22565
rect 3973 22525 3985 22559
rect 4019 22556 4031 22559
rect 4246 22556 4252 22568
rect 4019 22528 4252 22556
rect 4019 22525 4031 22528
rect 3973 22519 4031 22525
rect 4246 22516 4252 22528
rect 4304 22516 4310 22568
rect 4614 22556 4620 22568
rect 4575 22528 4620 22556
rect 4614 22516 4620 22528
rect 4672 22556 4678 22568
rect 5442 22556 5448 22568
rect 4672 22528 5448 22556
rect 4672 22516 4678 22528
rect 5442 22516 5448 22528
rect 5500 22516 5506 22568
rect 5994 22516 6000 22568
rect 6052 22556 6058 22568
rect 6454 22556 6460 22568
rect 6052 22528 6460 22556
rect 6052 22516 6058 22528
rect 6454 22516 6460 22528
rect 6512 22556 6518 22568
rect 6825 22559 6883 22565
rect 6825 22556 6837 22559
rect 6512 22528 6837 22556
rect 6512 22516 6518 22528
rect 6825 22525 6837 22528
rect 6871 22525 6883 22559
rect 6825 22519 6883 22525
rect 6914 22516 6920 22568
rect 6972 22556 6978 22568
rect 7009 22559 7067 22565
rect 7009 22556 7021 22559
rect 6972 22528 7021 22556
rect 6972 22516 6978 22528
rect 7009 22525 7021 22528
rect 7055 22525 7067 22559
rect 7009 22519 7067 22525
rect 7377 22559 7435 22565
rect 7377 22525 7389 22559
rect 7423 22556 7435 22559
rect 7650 22556 7656 22568
rect 7423 22528 7656 22556
rect 7423 22525 7435 22528
rect 7377 22519 7435 22525
rect 1845 22509 1903 22515
rect 3237 22491 3295 22497
rect 3237 22457 3249 22491
rect 3283 22488 3295 22491
rect 7024 22488 7052 22519
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 7742 22488 7748 22500
rect 3283 22460 5488 22488
rect 7024 22460 7748 22488
rect 3283 22457 3295 22460
rect 3237 22451 3295 22457
rect 2222 22420 2228 22432
rect 1780 22392 2228 22420
rect 2222 22380 2228 22392
rect 2280 22380 2286 22432
rect 3881 22423 3939 22429
rect 3881 22389 3893 22423
rect 3927 22420 3939 22423
rect 4154 22420 4160 22432
rect 3927 22392 4160 22420
rect 3927 22389 3939 22392
rect 3881 22383 3939 22389
rect 4154 22380 4160 22392
rect 4212 22420 4218 22432
rect 4798 22420 4804 22432
rect 4212 22392 4804 22420
rect 4212 22380 4218 22392
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 5460 22420 5488 22460
rect 7742 22448 7748 22460
rect 7800 22448 7806 22500
rect 7852 22488 7880 22596
rect 8128 22565 8156 22664
rect 8478 22652 8484 22664
rect 8536 22692 8542 22704
rect 9122 22692 9128 22704
rect 8536 22664 9128 22692
rect 8536 22652 8542 22664
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 9674 22692 9680 22704
rect 9508 22664 9680 22692
rect 8386 22624 8392 22636
rect 8347 22596 8392 22624
rect 8386 22584 8392 22596
rect 8444 22584 8450 22636
rect 9508 22633 9536 22664
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22593 9551 22627
rect 9493 22587 9551 22593
rect 9585 22627 9643 22633
rect 9585 22593 9597 22627
rect 9631 22624 9643 22627
rect 9950 22624 9956 22636
rect 9631 22596 9956 22624
rect 9631 22593 9643 22596
rect 9585 22587 9643 22593
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 8113 22559 8171 22565
rect 8113 22525 8125 22559
rect 8159 22525 8171 22559
rect 8113 22519 8171 22525
rect 8205 22559 8263 22565
rect 8205 22525 8217 22559
rect 8251 22556 8263 22559
rect 8754 22556 8760 22568
rect 8251 22528 8760 22556
rect 8251 22525 8263 22528
rect 8205 22519 8263 22525
rect 8220 22488 8248 22519
rect 8754 22516 8760 22528
rect 8812 22516 8818 22568
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 9766 22556 9772 22568
rect 9723 22528 9772 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 9766 22516 9772 22528
rect 9824 22516 9830 22568
rect 10226 22516 10232 22568
rect 10284 22556 10290 22568
rect 10796 22565 10824 22732
rect 10870 22720 10876 22732
rect 10928 22720 10934 22772
rect 12710 22760 12716 22772
rect 11164 22732 12716 22760
rect 10873 22627 10931 22633
rect 10873 22593 10885 22627
rect 10919 22624 10931 22627
rect 11054 22624 11060 22636
rect 10919 22596 11060 22624
rect 10919 22593 10931 22596
rect 10873 22587 10931 22593
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 10597 22559 10655 22565
rect 10597 22556 10609 22559
rect 10284 22528 10609 22556
rect 10284 22516 10290 22528
rect 10597 22525 10609 22528
rect 10643 22525 10655 22559
rect 10597 22519 10655 22525
rect 10781 22559 10839 22565
rect 10781 22525 10793 22559
rect 10827 22525 10839 22559
rect 10781 22519 10839 22525
rect 10962 22516 10968 22568
rect 11020 22556 11026 22568
rect 11164 22565 11192 22732
rect 12710 22720 12716 22732
rect 12768 22760 12774 22772
rect 13354 22760 13360 22772
rect 12768 22732 13360 22760
rect 12768 22720 12774 22732
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 13538 22720 13544 22772
rect 13596 22760 13602 22772
rect 19518 22760 19524 22772
rect 13596 22732 19524 22760
rect 13596 22720 13602 22732
rect 19518 22720 19524 22732
rect 19576 22720 19582 22772
rect 19613 22763 19671 22769
rect 19613 22729 19625 22763
rect 19659 22760 19671 22763
rect 19702 22760 19708 22772
rect 19659 22732 19708 22760
rect 19659 22729 19671 22732
rect 19613 22723 19671 22729
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 21358 22760 21364 22772
rect 20088 22732 21364 22760
rect 18414 22652 18420 22704
rect 18472 22692 18478 22704
rect 20088 22692 20116 22732
rect 21358 22720 21364 22732
rect 21416 22720 21422 22772
rect 22094 22760 22100 22772
rect 21744 22732 22100 22760
rect 18472 22664 20116 22692
rect 18472 22652 18478 22664
rect 14737 22627 14795 22633
rect 14737 22593 14749 22627
rect 14783 22624 14795 22627
rect 14918 22624 14924 22636
rect 14783 22596 14924 22624
rect 14783 22593 14795 22596
rect 14737 22587 14795 22593
rect 14918 22584 14924 22596
rect 14976 22584 14982 22636
rect 18690 22584 18696 22636
rect 18748 22584 18754 22636
rect 21744 22633 21772 22732
rect 22094 22720 22100 22732
rect 22152 22720 22158 22772
rect 22370 22720 22376 22772
rect 22428 22760 22434 22772
rect 22922 22760 22928 22772
rect 22428 22732 22928 22760
rect 22428 22720 22434 22732
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 23106 22760 23112 22772
rect 23067 22732 23112 22760
rect 23106 22720 23112 22732
rect 23164 22720 23170 22772
rect 23845 22763 23903 22769
rect 23845 22729 23857 22763
rect 23891 22760 23903 22763
rect 24397 22763 24455 22769
rect 24397 22760 24409 22763
rect 23891 22732 24409 22760
rect 23891 22729 23903 22732
rect 23845 22723 23903 22729
rect 24397 22729 24409 22732
rect 24443 22760 24455 22763
rect 24854 22760 24860 22772
rect 24443 22732 24860 22760
rect 24443 22729 24455 22732
rect 24397 22723 24455 22729
rect 24854 22720 24860 22732
rect 24912 22760 24918 22772
rect 25038 22760 25044 22772
rect 24912 22732 25044 22760
rect 24912 22720 24918 22732
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 26513 22763 26571 22769
rect 26513 22729 26525 22763
rect 26559 22760 26571 22763
rect 26602 22760 26608 22772
rect 26559 22732 26608 22760
rect 26559 22729 26571 22732
rect 26513 22723 26571 22729
rect 26602 22720 26608 22732
rect 26660 22720 26666 22772
rect 26418 22652 26424 22704
rect 26476 22692 26482 22704
rect 27522 22692 27528 22704
rect 26476 22664 27528 22692
rect 26476 22652 26482 22664
rect 26988 22633 27016 22664
rect 27522 22652 27528 22664
rect 27580 22652 27586 22704
rect 28718 22652 28724 22704
rect 28776 22692 28782 22704
rect 29549 22695 29607 22701
rect 29549 22692 29561 22695
rect 28776 22664 29561 22692
rect 28776 22652 28782 22664
rect 29549 22661 29561 22664
rect 29595 22661 29607 22695
rect 29549 22655 29607 22661
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22624 21051 22627
rect 21729 22627 21787 22633
rect 21729 22624 21741 22627
rect 21039 22596 21741 22624
rect 21039 22593 21051 22596
rect 20993 22587 21051 22593
rect 21729 22593 21741 22596
rect 21775 22593 21787 22627
rect 26973 22627 27031 22633
rect 21729 22587 21787 22593
rect 25700 22596 26832 22624
rect 11149 22559 11207 22565
rect 11020 22528 11065 22556
rect 11020 22516 11026 22528
rect 11149 22525 11161 22559
rect 11195 22525 11207 22559
rect 11149 22519 11207 22525
rect 11606 22516 11612 22568
rect 11664 22556 11670 22568
rect 11793 22559 11851 22565
rect 11793 22556 11805 22559
rect 11664 22528 11805 22556
rect 11664 22516 11670 22528
rect 11793 22525 11805 22528
rect 11839 22556 11851 22559
rect 11882 22556 11888 22568
rect 11839 22528 11888 22556
rect 11839 22525 11851 22528
rect 11793 22519 11851 22525
rect 11882 22516 11888 22528
rect 11940 22516 11946 22568
rect 14461 22559 14519 22565
rect 14461 22525 14473 22559
rect 14507 22556 14519 22559
rect 15286 22556 15292 22568
rect 14507 22528 15292 22556
rect 14507 22525 14519 22528
rect 14461 22519 14519 22525
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 15746 22556 15752 22568
rect 15707 22528 15752 22556
rect 15746 22516 15752 22528
rect 15804 22516 15810 22568
rect 16022 22565 16028 22568
rect 16016 22556 16028 22565
rect 15983 22528 16028 22556
rect 16016 22519 16028 22528
rect 16022 22516 16028 22519
rect 16080 22516 16086 22568
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 17589 22559 17647 22565
rect 17589 22556 17601 22559
rect 17552 22528 17601 22556
rect 17552 22516 17558 22528
rect 17589 22525 17601 22528
rect 17635 22525 17647 22559
rect 17954 22556 17960 22568
rect 17915 22528 17960 22556
rect 17589 22519 17647 22525
rect 17954 22516 17960 22528
rect 18012 22516 18018 22568
rect 18414 22556 18420 22568
rect 18375 22528 18420 22556
rect 18414 22516 18420 22528
rect 18472 22516 18478 22568
rect 18708 22556 18736 22584
rect 25700 22556 25728 22596
rect 18708 22528 25728 22556
rect 25777 22559 25835 22565
rect 25777 22525 25789 22559
rect 25823 22556 25835 22559
rect 26234 22556 26240 22568
rect 25823 22528 26240 22556
rect 25823 22525 25835 22528
rect 25777 22519 25835 22525
rect 26234 22516 26240 22528
rect 26292 22516 26298 22568
rect 26697 22559 26755 22565
rect 26697 22525 26709 22559
rect 26743 22525 26755 22559
rect 26697 22519 26755 22525
rect 7852 22460 8248 22488
rect 11333 22491 11391 22497
rect 11333 22457 11345 22491
rect 11379 22488 11391 22491
rect 12038 22491 12096 22497
rect 12038 22488 12050 22491
rect 11379 22460 12050 22488
rect 11379 22457 11391 22460
rect 11333 22451 11391 22457
rect 12038 22457 12050 22460
rect 12084 22457 12096 22491
rect 12038 22451 12096 22457
rect 15838 22448 15844 22500
rect 15896 22488 15902 22500
rect 16298 22488 16304 22500
rect 15896 22460 16304 22488
rect 15896 22448 15902 22460
rect 16298 22448 16304 22460
rect 16356 22448 16362 22500
rect 18693 22491 18751 22497
rect 18693 22457 18705 22491
rect 18739 22488 18751 22491
rect 19794 22488 19800 22500
rect 18739 22460 19800 22488
rect 18739 22457 18751 22460
rect 18693 22451 18751 22457
rect 19794 22448 19800 22460
rect 19852 22448 19858 22500
rect 20726 22491 20784 22497
rect 20726 22488 20738 22491
rect 19895 22460 20738 22488
rect 7098 22420 7104 22432
rect 5460 22392 7104 22420
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 7558 22420 7564 22432
rect 7519 22392 7564 22420
rect 7558 22380 7564 22392
rect 7616 22380 7622 22432
rect 7650 22380 7656 22432
rect 7708 22420 7714 22432
rect 8018 22420 8024 22432
rect 7708 22392 8024 22420
rect 7708 22380 7714 22392
rect 8018 22380 8024 22392
rect 8076 22380 8082 22432
rect 8294 22380 8300 22432
rect 8352 22420 8358 22432
rect 9582 22420 9588 22432
rect 8352 22392 9588 22420
rect 8352 22380 8358 22392
rect 9582 22380 9588 22392
rect 9640 22380 9646 22432
rect 13173 22423 13231 22429
rect 13173 22389 13185 22423
rect 13219 22420 13231 22423
rect 13354 22420 13360 22432
rect 13219 22392 13360 22420
rect 13219 22389 13231 22392
rect 13173 22383 13231 22389
rect 13354 22380 13360 22392
rect 13412 22380 13418 22432
rect 15286 22380 15292 22432
rect 15344 22420 15350 22432
rect 15470 22420 15476 22432
rect 15344 22392 15476 22420
rect 15344 22380 15350 22392
rect 15470 22380 15476 22392
rect 15528 22380 15534 22432
rect 17129 22423 17187 22429
rect 17129 22389 17141 22423
rect 17175 22420 17187 22423
rect 17310 22420 17316 22432
rect 17175 22392 17316 22420
rect 17175 22389 17187 22392
rect 17129 22383 17187 22389
rect 17310 22380 17316 22392
rect 17368 22380 17374 22432
rect 19426 22380 19432 22432
rect 19484 22420 19490 22432
rect 19895 22420 19923 22460
rect 20726 22457 20738 22460
rect 20772 22457 20784 22491
rect 20726 22451 20784 22457
rect 21266 22448 21272 22500
rect 21324 22488 21330 22500
rect 21974 22491 22032 22497
rect 21974 22488 21986 22491
rect 21324 22460 21986 22488
rect 21324 22448 21330 22460
rect 21974 22457 21986 22460
rect 22020 22457 22032 22491
rect 21974 22451 22032 22457
rect 25130 22448 25136 22500
rect 25188 22488 25194 22500
rect 25510 22491 25568 22497
rect 25510 22488 25522 22491
rect 25188 22460 25522 22488
rect 25188 22448 25194 22460
rect 25510 22457 25522 22460
rect 25556 22457 25568 22491
rect 25510 22451 25568 22457
rect 19484 22392 19923 22420
rect 26712 22420 26740 22519
rect 26804 22488 26832 22596
rect 26973 22593 26985 22627
rect 27019 22593 27031 22627
rect 28442 22624 28448 22636
rect 28403 22596 28448 22624
rect 26973 22587 27031 22593
rect 28442 22584 28448 22596
rect 28500 22584 28506 22636
rect 28534 22584 28540 22636
rect 28592 22624 28598 22636
rect 30926 22624 30932 22636
rect 28592 22596 28637 22624
rect 30887 22596 30932 22624
rect 28592 22584 28598 22596
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 26878 22516 26884 22568
rect 26936 22556 26942 22568
rect 26936 22528 26981 22556
rect 26936 22516 26942 22528
rect 27062 22516 27068 22568
rect 27120 22556 27126 22568
rect 27246 22556 27252 22568
rect 27120 22528 27165 22556
rect 27207 22528 27252 22556
rect 27120 22516 27126 22528
rect 27246 22516 27252 22528
rect 27304 22516 27310 22568
rect 28166 22556 28172 22568
rect 28127 22528 28172 22556
rect 28166 22516 28172 22528
rect 28224 22516 28230 22568
rect 28353 22559 28411 22565
rect 28353 22525 28365 22559
rect 28399 22525 28411 22559
rect 28718 22556 28724 22568
rect 28679 22528 28724 22556
rect 28353 22519 28411 22525
rect 28258 22488 28264 22500
rect 26804 22460 28264 22488
rect 28258 22448 28264 22460
rect 28316 22448 28322 22500
rect 28368 22488 28396 22519
rect 28718 22516 28724 22528
rect 28776 22516 28782 22568
rect 28810 22488 28816 22500
rect 28368 22460 28816 22488
rect 28810 22448 28816 22460
rect 28868 22448 28874 22500
rect 28905 22491 28963 22497
rect 28905 22457 28917 22491
rect 28951 22488 28963 22491
rect 30662 22491 30720 22497
rect 30662 22488 30674 22491
rect 28951 22460 30674 22488
rect 28951 22457 28963 22460
rect 28905 22451 28963 22457
rect 30662 22457 30674 22460
rect 30708 22457 30720 22491
rect 30662 22451 30720 22457
rect 29362 22420 29368 22432
rect 26712 22392 29368 22420
rect 19484 22380 19490 22392
rect 29362 22380 29368 22392
rect 29420 22380 29426 22432
rect 1104 22330 32016 22352
rect 1104 22278 11253 22330
rect 11305 22278 11317 22330
rect 11369 22278 11381 22330
rect 11433 22278 11445 22330
rect 11497 22278 11509 22330
rect 11561 22278 21557 22330
rect 21609 22278 21621 22330
rect 21673 22278 21685 22330
rect 21737 22278 21749 22330
rect 21801 22278 21813 22330
rect 21865 22278 32016 22330
rect 1104 22256 32016 22278
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 7650 22216 7656 22228
rect 7524 22188 7656 22216
rect 7524 22176 7530 22188
rect 7650 22176 7656 22188
rect 7708 22176 7714 22228
rect 9490 22176 9496 22228
rect 9548 22176 9554 22228
rect 11054 22216 11060 22228
rect 10520 22188 11060 22216
rect 5902 22148 5908 22160
rect 5828 22120 5908 22148
rect 1394 22080 1400 22092
rect 1355 22052 1400 22080
rect 1394 22040 1400 22052
rect 1452 22040 1458 22092
rect 1670 22089 1676 22092
rect 1664 22043 1676 22089
rect 1728 22080 1734 22092
rect 3234 22080 3240 22092
rect 1728 22052 1764 22080
rect 3195 22052 3240 22080
rect 1670 22040 1676 22043
rect 1728 22040 1734 22052
rect 3234 22040 3240 22052
rect 3292 22040 3298 22092
rect 3418 22080 3424 22092
rect 3379 22052 3424 22080
rect 3418 22040 3424 22052
rect 3476 22040 3482 22092
rect 3602 22080 3608 22092
rect 3563 22052 3608 22080
rect 3602 22040 3608 22052
rect 3660 22040 3666 22092
rect 3789 22083 3847 22089
rect 3789 22049 3801 22083
rect 3835 22049 3847 22083
rect 3789 22043 3847 22049
rect 3973 22083 4031 22089
rect 3973 22049 3985 22083
rect 4019 22080 4031 22083
rect 4062 22080 4068 22092
rect 4019 22052 4068 22080
rect 4019 22049 4031 22052
rect 3973 22043 4031 22049
rect 3697 22015 3755 22021
rect 3697 21981 3709 22015
rect 3743 21981 3755 22015
rect 3804 22012 3832 22043
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 5258 22040 5264 22092
rect 5316 22080 5322 22092
rect 5546 22083 5604 22089
rect 5546 22080 5558 22083
rect 5316 22052 5558 22080
rect 5316 22040 5322 22052
rect 5546 22049 5558 22052
rect 5592 22049 5604 22083
rect 5546 22043 5604 22049
rect 5718 22040 5724 22092
rect 5776 22040 5782 22092
rect 5828 22089 5856 22120
rect 5902 22108 5908 22120
rect 5960 22108 5966 22160
rect 9508 22148 9536 22176
rect 9048 22120 9536 22148
rect 6822 22089 6828 22092
rect 5813 22083 5871 22089
rect 5813 22049 5825 22083
rect 5859 22080 5871 22083
rect 6816 22080 6828 22089
rect 5859 22052 5961 22080
rect 6783 22052 6828 22080
rect 5859 22050 5948 22052
rect 5859 22049 5871 22050
rect 5813 22043 5871 22049
rect 4430 22012 4436 22024
rect 3804 21984 4436 22012
rect 3697 21975 3755 21981
rect 3712 21944 3740 21975
rect 4430 21972 4436 21984
rect 4488 21972 4494 22024
rect 5736 22012 5764 22040
rect 5920 22012 5948 22050
rect 6816 22043 6828 22052
rect 6822 22040 6828 22043
rect 6880 22040 6886 22092
rect 9048 22089 9076 22120
rect 9033 22083 9091 22089
rect 9033 22049 9045 22083
rect 9079 22080 9091 22083
rect 9217 22083 9275 22089
rect 9079 22052 9113 22080
rect 9079 22049 9091 22052
rect 9033 22043 9091 22049
rect 9217 22049 9229 22083
rect 9263 22049 9275 22083
rect 9217 22043 9275 22049
rect 9585 22083 9643 22089
rect 9585 22049 9597 22083
rect 9631 22080 9643 22083
rect 9950 22080 9956 22092
rect 9631 22052 9956 22080
rect 9631 22049 9643 22052
rect 9585 22043 9643 22049
rect 6546 22012 6552 22024
rect 5736 21984 5856 22012
rect 5920 21984 6552 22012
rect 5828 21944 5856 21984
rect 6546 21972 6552 21984
rect 6604 21972 6610 22024
rect 8849 22015 8907 22021
rect 8849 21981 8861 22015
rect 8895 22012 8907 22015
rect 8938 22012 8944 22024
rect 8895 21984 8944 22012
rect 8895 21981 8907 21984
rect 8849 21975 8907 21981
rect 8938 21972 8944 21984
rect 8996 21972 9002 22024
rect 5902 21944 5908 21956
rect 3712 21916 4936 21944
rect 5828 21916 5908 21944
rect 2314 21836 2320 21888
rect 2372 21876 2378 21888
rect 2777 21879 2835 21885
rect 2777 21876 2789 21879
rect 2372 21848 2789 21876
rect 2372 21836 2378 21848
rect 2777 21845 2789 21848
rect 2823 21845 2835 21879
rect 4430 21876 4436 21888
rect 4391 21848 4436 21876
rect 2777 21839 2835 21845
rect 4430 21836 4436 21848
rect 4488 21836 4494 21888
rect 4908 21876 4936 21916
rect 5902 21904 5908 21916
rect 5960 21904 5966 21956
rect 6270 21904 6276 21956
rect 6328 21904 6334 21956
rect 9122 21904 9128 21956
rect 9180 21944 9186 21956
rect 9232 21944 9260 22043
rect 9950 22040 9956 22052
rect 10008 22040 10014 22092
rect 10226 22080 10232 22092
rect 10187 22052 10232 22080
rect 10226 22040 10232 22052
rect 10284 22040 10290 22092
rect 10410 22080 10416 22092
rect 10371 22052 10416 22080
rect 10410 22040 10416 22052
rect 10468 22040 10474 22092
rect 10520 22021 10548 22188
rect 11054 22176 11060 22188
rect 11112 22176 11118 22228
rect 15838 22176 15844 22228
rect 15896 22216 15902 22228
rect 19242 22216 19248 22228
rect 15896 22188 19248 22216
rect 15896 22176 15902 22188
rect 19242 22176 19248 22188
rect 19300 22176 19306 22228
rect 20990 22216 20996 22228
rect 19536 22188 20996 22216
rect 11146 22148 11152 22160
rect 10796 22120 11152 22148
rect 10796 22089 10824 22120
rect 11146 22108 11152 22120
rect 11204 22108 11210 22160
rect 16298 22148 16304 22160
rect 11440 22120 11744 22148
rect 10781 22083 10839 22089
rect 10781 22049 10793 22083
rect 10827 22049 10839 22083
rect 10781 22043 10839 22049
rect 10965 22083 11023 22089
rect 10965 22049 10977 22083
rect 11011 22080 11023 22083
rect 11440 22080 11468 22120
rect 11011 22052 11468 22080
rect 11011 22049 11023 22052
rect 10965 22043 11023 22049
rect 11606 22040 11612 22092
rect 11664 22040 11670 22092
rect 11716 22080 11744 22120
rect 14660 22120 16304 22148
rect 11773 22083 11831 22089
rect 11773 22080 11785 22083
rect 11716 22052 11785 22080
rect 11773 22049 11785 22052
rect 11819 22049 11831 22083
rect 13354 22080 13360 22092
rect 13315 22052 13360 22080
rect 11773 22043 11831 22049
rect 13354 22040 13360 22052
rect 13412 22040 13418 22092
rect 13446 22040 13452 22092
rect 13504 22080 13510 22092
rect 14660 22089 14688 22120
rect 16298 22108 16304 22120
rect 16356 22148 16362 22160
rect 19334 22148 19340 22160
rect 16356 22120 17356 22148
rect 16356 22108 16362 22120
rect 17328 22092 17356 22120
rect 18432 22120 19340 22148
rect 14645 22083 14703 22089
rect 13504 22052 13549 22080
rect 13504 22040 13510 22052
rect 14645 22049 14657 22083
rect 14691 22049 14703 22083
rect 14645 22043 14703 22049
rect 15933 22083 15991 22089
rect 15933 22049 15945 22083
rect 15979 22080 15991 22083
rect 16206 22080 16212 22092
rect 15979 22052 16212 22080
rect 15979 22049 15991 22052
rect 15933 22043 15991 22049
rect 16206 22040 16212 22052
rect 16264 22040 16270 22092
rect 16761 22083 16819 22089
rect 16761 22049 16773 22083
rect 16807 22080 16819 22083
rect 16850 22080 16856 22092
rect 16807 22052 16856 22080
rect 16807 22049 16819 22052
rect 16761 22043 16819 22049
rect 16850 22040 16856 22052
rect 16908 22040 16914 22092
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 17037 22083 17095 22089
rect 17037 22049 17049 22083
rect 17083 22080 17095 22083
rect 17218 22080 17224 22092
rect 17083 22052 17224 22080
rect 17083 22049 17095 22052
rect 17037 22043 17095 22049
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 10505 22015 10563 22021
rect 10505 21981 10517 22015
rect 10551 21981 10563 22015
rect 10505 21975 10563 21981
rect 9180 21916 9260 21944
rect 9180 21904 9186 21916
rect 5810 21876 5816 21888
rect 4908 21848 5816 21876
rect 5810 21836 5816 21848
rect 5868 21876 5874 21888
rect 6288 21876 6316 21904
rect 5868 21848 6316 21876
rect 5868 21836 5874 21848
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 7929 21879 7987 21885
rect 7929 21876 7941 21879
rect 7800 21848 7941 21876
rect 7800 21836 7806 21848
rect 7929 21845 7941 21848
rect 7975 21845 7987 21879
rect 7929 21839 7987 21845
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 9416 21876 9444 21975
rect 8904 21848 9444 21876
rect 10520 21876 10548 21975
rect 10594 21972 10600 22024
rect 10652 22012 10658 22024
rect 10652 21984 10697 22012
rect 10652 21972 10658 21984
rect 11054 21972 11060 22024
rect 11112 22012 11118 22024
rect 11517 22015 11575 22021
rect 11517 22012 11529 22015
rect 11112 21984 11529 22012
rect 11112 21972 11118 21984
rect 11517 21981 11529 21984
rect 11563 22012 11575 22015
rect 11624 22012 11652 22040
rect 11563 21984 11652 22012
rect 11563 21981 11575 21984
rect 11517 21975 11575 21981
rect 15562 21972 15568 22024
rect 15620 22012 15626 22024
rect 15657 22015 15715 22021
rect 15657 22012 15669 22015
rect 15620 21984 15669 22012
rect 15620 21972 15626 21984
rect 15657 21981 15669 21984
rect 15703 21981 15715 22015
rect 16482 22012 16488 22024
rect 15657 21975 15715 21981
rect 15856 21984 16488 22012
rect 14553 21947 14611 21953
rect 14553 21913 14565 21947
rect 14599 21944 14611 21947
rect 15856 21944 15884 21984
rect 16482 21972 16488 21984
rect 16540 22012 16546 22024
rect 16960 22012 16988 22043
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 17494 22080 17500 22092
rect 17368 22052 17413 22080
rect 17455 22052 17500 22080
rect 17368 22040 17374 22052
rect 17494 22040 17500 22052
rect 17552 22040 17558 22092
rect 18432 22089 18460 22120
rect 19334 22108 19340 22120
rect 19392 22108 19398 22160
rect 18417 22083 18475 22089
rect 18417 22049 18429 22083
rect 18463 22080 18475 22083
rect 18598 22080 18604 22092
rect 18463 22052 18497 22080
rect 18559 22052 18604 22080
rect 18463 22049 18475 22052
rect 18417 22043 18475 22049
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 18969 22083 19027 22089
rect 18969 22049 18981 22083
rect 19015 22080 19027 22083
rect 19536 22080 19564 22188
rect 20990 22176 20996 22188
rect 21048 22176 21054 22228
rect 22094 22176 22100 22228
rect 22152 22216 22158 22228
rect 23290 22216 23296 22228
rect 22152 22188 23296 22216
rect 22152 22176 22158 22188
rect 23290 22176 23296 22188
rect 23348 22216 23354 22228
rect 23477 22219 23535 22225
rect 23477 22216 23489 22219
rect 23348 22188 23489 22216
rect 23348 22176 23354 22188
rect 23477 22185 23489 22188
rect 23523 22185 23535 22219
rect 23477 22179 23535 22185
rect 24946 22176 24952 22228
rect 25004 22176 25010 22228
rect 25130 22216 25136 22228
rect 25091 22188 25136 22216
rect 25130 22176 25136 22188
rect 25188 22176 25194 22228
rect 26418 22216 26424 22228
rect 26379 22188 26424 22216
rect 26418 22176 26424 22188
rect 26476 22176 26482 22228
rect 27065 22219 27123 22225
rect 27065 22185 27077 22219
rect 27111 22216 27123 22219
rect 27154 22216 27160 22228
rect 27111 22188 27160 22216
rect 27111 22185 27123 22188
rect 27065 22179 27123 22185
rect 27154 22176 27160 22188
rect 27212 22176 27218 22228
rect 22189 22151 22247 22157
rect 19812 22120 20116 22148
rect 19812 22080 19840 22120
rect 19886 22089 19892 22092
rect 19015 22052 19564 22080
rect 19628 22052 19840 22080
rect 19015 22049 19027 22052
rect 18969 22043 19027 22049
rect 19628 22024 19656 22052
rect 19880 22043 19892 22089
rect 19944 22080 19950 22092
rect 20088 22080 20116 22120
rect 22189 22117 22201 22151
rect 22235 22148 22247 22151
rect 23014 22148 23020 22160
rect 22235 22120 23020 22148
rect 22235 22117 22247 22120
rect 22189 22111 22247 22117
rect 23014 22108 23020 22120
rect 23072 22108 23078 22160
rect 24964 22148 24992 22176
rect 24872 22120 24992 22148
rect 22094 22080 22100 22092
rect 19944 22052 19980 22080
rect 20088 22052 22100 22080
rect 19886 22040 19892 22043
rect 19944 22040 19950 22052
rect 22066 22040 22100 22052
rect 22152 22040 22158 22092
rect 24397 22083 24455 22089
rect 24397 22082 24409 22083
rect 24320 22080 24409 22082
rect 23860 22054 24409 22080
rect 23860 22052 24348 22054
rect 16540 21984 16988 22012
rect 17129 22015 17187 22021
rect 16540 21972 16546 21984
rect 17129 21981 17141 22015
rect 17175 22012 17187 22015
rect 18046 22012 18052 22024
rect 17175 21984 18052 22012
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18693 22015 18751 22021
rect 18693 21981 18705 22015
rect 18739 21981 18751 22015
rect 18693 21975 18751 21981
rect 14599 21916 15884 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 17954 21904 17960 21956
rect 18012 21944 18018 21956
rect 18708 21944 18736 21975
rect 18782 21972 18788 22024
rect 18840 22012 18846 22024
rect 19610 22012 19616 22024
rect 18840 21984 18885 22012
rect 19571 21984 19616 22012
rect 18840 21972 18846 21984
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 22066 22012 22094 22040
rect 23860 22024 23888 22052
rect 24397 22049 24409 22054
rect 24443 22049 24455 22083
rect 24397 22043 24455 22049
rect 24581 22083 24639 22089
rect 24581 22049 24593 22083
rect 24627 22080 24639 22083
rect 24872 22080 24900 22120
rect 25958 22108 25964 22160
rect 26016 22148 26022 22160
rect 26053 22151 26111 22157
rect 26053 22148 26065 22151
rect 26016 22120 26065 22148
rect 26016 22108 26022 22120
rect 26053 22117 26065 22120
rect 26099 22117 26111 22151
rect 26053 22111 26111 22117
rect 26237 22151 26295 22157
rect 26237 22117 26249 22151
rect 26283 22148 26295 22151
rect 26326 22148 26332 22160
rect 26283 22120 26332 22148
rect 26283 22117 26295 22120
rect 26237 22111 26295 22117
rect 26326 22108 26332 22120
rect 26384 22148 26390 22160
rect 28718 22148 28724 22160
rect 26384 22120 27016 22148
rect 26384 22108 26390 22120
rect 24627 22052 24900 22080
rect 24949 22083 25007 22089
rect 24627 22049 24639 22052
rect 24581 22043 24639 22049
rect 24949 22049 24961 22083
rect 24995 22080 25007 22083
rect 25038 22080 25044 22092
rect 24995 22052 25044 22080
rect 24995 22049 25007 22052
rect 24949 22043 25007 22049
rect 25038 22040 25044 22052
rect 25096 22040 25102 22092
rect 26988 22089 27016 22120
rect 28276 22120 28724 22148
rect 26973 22083 27031 22089
rect 26973 22049 26985 22083
rect 27019 22049 27031 22083
rect 26973 22043 27031 22049
rect 27522 22040 27528 22092
rect 27580 22080 27586 22092
rect 28077 22083 28135 22089
rect 28077 22080 28089 22083
rect 27580 22052 28089 22080
rect 27580 22040 27586 22052
rect 28077 22049 28089 22052
rect 28123 22080 28135 22083
rect 28166 22080 28172 22092
rect 28123 22052 28172 22080
rect 28123 22049 28135 22052
rect 28077 22043 28135 22049
rect 28166 22040 28172 22052
rect 28224 22040 28230 22092
rect 28276 22087 28304 22120
rect 28718 22108 28724 22120
rect 28776 22108 28782 22160
rect 28261 22081 28319 22087
rect 28261 22047 28273 22081
rect 28307 22047 28319 22081
rect 28261 22041 28319 22047
rect 28445 22083 28503 22089
rect 28445 22049 28457 22083
rect 28491 22049 28503 22083
rect 28626 22080 28632 22092
rect 28587 22052 28632 22080
rect 28445 22043 28503 22049
rect 22278 22012 22284 22024
rect 22066 21984 22284 22012
rect 22278 21972 22284 21984
rect 22336 21972 22342 22024
rect 23842 21972 23848 22024
rect 23900 21972 23906 22024
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 18012 21916 18736 21944
rect 24688 21944 24716 21975
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 28350 22012 28356 22024
rect 24820 21984 24865 22012
rect 28311 21984 28356 22012
rect 24820 21972 24826 21984
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 28460 22012 28488 22043
rect 28626 22040 28632 22052
rect 28684 22040 28690 22092
rect 29273 22083 29331 22089
rect 29273 22049 29285 22083
rect 29319 22049 29331 22083
rect 29273 22043 29331 22049
rect 28534 22012 28540 22024
rect 28460 21984 28540 22012
rect 28534 21972 28540 21984
rect 28592 21972 28598 22024
rect 24854 21944 24860 21956
rect 24688 21916 24860 21944
rect 18012 21904 18018 21916
rect 24854 21904 24860 21916
rect 24912 21944 24918 21956
rect 26050 21944 26056 21956
rect 24912 21916 26056 21944
rect 24912 21904 24918 21916
rect 26050 21904 26056 21916
rect 26108 21904 26114 21956
rect 28166 21904 28172 21956
rect 28224 21944 28230 21956
rect 28718 21944 28724 21956
rect 28224 21916 28724 21944
rect 28224 21904 28230 21916
rect 28718 21904 28724 21916
rect 28776 21944 28782 21956
rect 29288 21944 29316 22043
rect 29362 22040 29368 22092
rect 29420 22080 29426 22092
rect 30469 22083 30527 22089
rect 29420 22052 29465 22080
rect 29420 22040 29426 22052
rect 30469 22049 30481 22083
rect 30515 22049 30527 22083
rect 31294 22080 31300 22092
rect 31255 22052 31300 22080
rect 30469 22043 30527 22049
rect 28776 21916 29316 21944
rect 28776 21904 28782 21916
rect 11882 21876 11888 21888
rect 10520 21848 11888 21876
rect 8904 21836 8910 21848
rect 11882 21836 11888 21848
rect 11940 21836 11946 21888
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 12897 21879 12955 21885
rect 12897 21876 12909 21879
rect 12492 21848 12909 21876
rect 12492 21836 12498 21848
rect 12897 21845 12909 21848
rect 12943 21845 12955 21879
rect 12897 21839 12955 21845
rect 19153 21879 19211 21885
rect 19153 21845 19165 21879
rect 19199 21876 19211 21879
rect 19886 21876 19892 21888
rect 19199 21848 19892 21876
rect 19199 21845 19211 21848
rect 19153 21839 19211 21845
rect 19886 21836 19892 21848
rect 19944 21836 19950 21888
rect 20346 21836 20352 21888
rect 20404 21876 20410 21888
rect 23658 21876 23664 21888
rect 20404 21848 23664 21876
rect 20404 21836 20410 21848
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 23934 21836 23940 21888
rect 23992 21876 23998 21888
rect 27062 21876 27068 21888
rect 23992 21848 27068 21876
rect 23992 21836 23998 21848
rect 27062 21836 27068 21848
rect 27120 21836 27126 21888
rect 28810 21876 28816 21888
rect 28771 21848 28816 21876
rect 28810 21836 28816 21848
rect 28868 21836 28874 21888
rect 28902 21836 28908 21888
rect 28960 21876 28966 21888
rect 29917 21879 29975 21885
rect 29917 21876 29929 21879
rect 28960 21848 29929 21876
rect 28960 21836 28966 21848
rect 29917 21845 29929 21848
rect 29963 21845 29975 21879
rect 30484 21876 30512 22043
rect 31294 22040 31300 22052
rect 31352 22040 31358 22092
rect 30653 21947 30711 21953
rect 30653 21913 30665 21947
rect 30699 21944 30711 21947
rect 30699 21916 31754 21944
rect 30699 21913 30711 21916
rect 30653 21907 30711 21913
rect 31113 21879 31171 21885
rect 31113 21876 31125 21879
rect 30484 21848 31125 21876
rect 29917 21839 29975 21845
rect 31113 21845 31125 21848
rect 31159 21845 31171 21879
rect 31726 21876 31754 21916
rect 31726 21848 32352 21876
rect 31113 21839 31171 21845
rect 1104 21786 32016 21808
rect 1104 21734 6102 21786
rect 6154 21734 6166 21786
rect 6218 21734 6230 21786
rect 6282 21734 6294 21786
rect 6346 21734 6358 21786
rect 6410 21734 16405 21786
rect 16457 21734 16469 21786
rect 16521 21734 16533 21786
rect 16585 21734 16597 21786
rect 16649 21734 16661 21786
rect 16713 21734 26709 21786
rect 26761 21734 26773 21786
rect 26825 21734 26837 21786
rect 26889 21734 26901 21786
rect 26953 21734 26965 21786
rect 27017 21734 32016 21786
rect 1104 21712 32016 21734
rect 1581 21675 1639 21681
rect 1581 21641 1593 21675
rect 1627 21672 1639 21675
rect 1670 21672 1676 21684
rect 1627 21644 1676 21672
rect 1627 21641 1639 21644
rect 1581 21635 1639 21641
rect 1670 21632 1676 21644
rect 1728 21632 1734 21684
rect 2406 21632 2412 21684
rect 2464 21672 2470 21684
rect 4614 21672 4620 21684
rect 2464 21644 4620 21672
rect 2464 21632 2470 21644
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 4706 21632 4712 21684
rect 4764 21672 4770 21684
rect 5258 21672 5264 21684
rect 4764 21644 4809 21672
rect 5219 21644 5264 21672
rect 4764 21632 4770 21644
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 8570 21632 8576 21684
rect 8628 21672 8634 21684
rect 9217 21675 9275 21681
rect 9217 21672 9229 21675
rect 8628 21644 9229 21672
rect 8628 21632 8634 21644
rect 9217 21641 9229 21644
rect 9263 21641 9275 21675
rect 9217 21635 9275 21641
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 13630 21672 13636 21684
rect 13228 21644 13636 21672
rect 13228 21632 13234 21644
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 14458 21672 14464 21684
rect 14419 21644 14464 21672
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 17773 21675 17831 21681
rect 14559 21644 16712 21672
rect 5810 21564 5816 21616
rect 5868 21564 5874 21616
rect 8938 21564 8944 21616
rect 8996 21604 9002 21616
rect 9401 21607 9459 21613
rect 9401 21604 9413 21607
rect 8996 21576 9413 21604
rect 8996 21564 9002 21576
rect 9401 21573 9413 21576
rect 9447 21573 9459 21607
rect 9401 21567 9459 21573
rect 11974 21564 11980 21616
rect 12032 21604 12038 21616
rect 14559 21604 14587 21644
rect 16684 21604 16712 21644
rect 17773 21641 17785 21675
rect 17819 21672 17831 21675
rect 18138 21672 18144 21684
rect 17819 21644 18144 21672
rect 17819 21641 17831 21644
rect 17773 21635 17831 21641
rect 18138 21632 18144 21644
rect 18196 21632 18202 21684
rect 18322 21632 18328 21684
rect 18380 21672 18386 21684
rect 18417 21675 18475 21681
rect 18417 21672 18429 21675
rect 18380 21644 18429 21672
rect 18380 21632 18386 21644
rect 18417 21641 18429 21644
rect 18463 21641 18475 21675
rect 19426 21672 19432 21684
rect 19387 21644 19432 21672
rect 18417 21635 18475 21641
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 21269 21675 21327 21681
rect 19536 21644 20116 21672
rect 19536 21604 19564 21644
rect 19978 21604 19984 21616
rect 12032 21576 14587 21604
rect 14660 21576 15700 21604
rect 16684 21576 19564 21604
rect 19904 21576 19984 21604
rect 12032 21564 12038 21576
rect 1946 21536 1952 21548
rect 1907 21508 1952 21536
rect 1946 21496 1952 21508
rect 2004 21496 2010 21548
rect 2498 21536 2504 21548
rect 2148 21508 2504 21536
rect 0 21468 800 21482
rect 1765 21471 1823 21477
rect 0 21440 1072 21468
rect 0 21426 800 21440
rect 1044 20992 1072 21440
rect 1765 21437 1777 21471
rect 1811 21437 1823 21471
rect 2038 21468 2044 21480
rect 1999 21440 2044 21468
rect 1765 21431 1823 21437
rect 1780 21400 1808 21431
rect 2038 21428 2044 21440
rect 2096 21428 2102 21480
rect 2148 21477 2176 21508
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 4798 21496 4804 21548
rect 4856 21536 4862 21548
rect 5074 21536 5080 21548
rect 4856 21508 5080 21536
rect 4856 21496 4862 21508
rect 5074 21496 5080 21508
rect 5132 21496 5138 21548
rect 5626 21536 5632 21548
rect 5587 21508 5632 21536
rect 5626 21496 5632 21508
rect 5684 21496 5690 21548
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21536 5779 21539
rect 5828 21536 5856 21564
rect 5767 21508 5856 21536
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 6546 21496 6552 21548
rect 6604 21536 6610 21548
rect 7009 21539 7067 21545
rect 7009 21536 7021 21539
rect 6604 21508 7021 21536
rect 6604 21496 6610 21508
rect 7009 21505 7021 21508
rect 7055 21505 7067 21539
rect 7009 21499 7067 21505
rect 9122 21496 9128 21548
rect 9180 21536 9186 21548
rect 9306 21536 9312 21548
rect 9180 21508 9312 21536
rect 9180 21496 9186 21508
rect 9306 21496 9312 21508
rect 9364 21496 9370 21548
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 9953 21539 10011 21545
rect 9953 21536 9965 21539
rect 9640 21508 9965 21536
rect 9640 21496 9646 21508
rect 9953 21505 9965 21508
rect 9999 21536 10011 21539
rect 10134 21536 10140 21548
rect 9999 21508 10140 21536
rect 9999 21505 10011 21508
rect 9953 21499 10011 21505
rect 10134 21496 10140 21508
rect 10192 21496 10198 21548
rect 10594 21496 10600 21548
rect 10652 21536 10658 21548
rect 10962 21536 10968 21548
rect 10652 21508 10968 21536
rect 10652 21496 10658 21508
rect 10962 21496 10968 21508
rect 11020 21536 11026 21548
rect 11020 21508 11560 21536
rect 11020 21496 11026 21508
rect 2133 21471 2191 21477
rect 2133 21437 2145 21471
rect 2179 21437 2191 21471
rect 2133 21431 2191 21437
rect 2222 21428 2228 21480
rect 2280 21468 2286 21480
rect 2317 21471 2375 21477
rect 2317 21468 2329 21471
rect 2280 21440 2329 21468
rect 2280 21428 2286 21440
rect 2317 21437 2329 21440
rect 2363 21437 2375 21471
rect 2317 21431 2375 21437
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 3786 21468 3792 21480
rect 3660 21440 3792 21468
rect 3660 21428 3666 21440
rect 3786 21428 3792 21440
rect 3844 21428 3850 21480
rect 4430 21428 4436 21480
rect 4488 21468 4494 21480
rect 5442 21468 5448 21480
rect 4488 21440 5448 21468
rect 4488 21428 4494 21440
rect 5442 21428 5448 21440
rect 5500 21428 5506 21480
rect 5810 21468 5816 21480
rect 5771 21440 5816 21468
rect 5810 21428 5816 21440
rect 5868 21428 5874 21480
rect 5994 21468 6000 21480
rect 5955 21440 6000 21468
rect 5994 21428 6000 21440
rect 6052 21468 6058 21480
rect 6454 21468 6460 21480
rect 6052 21440 6460 21468
rect 6052 21428 6058 21440
rect 6454 21428 6460 21440
rect 6512 21428 6518 21480
rect 7276 21471 7334 21477
rect 7276 21437 7288 21471
rect 7322 21468 7334 21471
rect 7558 21468 7564 21480
rect 7322 21440 7564 21468
rect 7322 21437 7334 21440
rect 7276 21431 7334 21437
rect 7558 21428 7564 21440
rect 7616 21428 7622 21480
rect 10226 21468 10232 21480
rect 10139 21440 10232 21468
rect 10226 21428 10232 21440
rect 10284 21428 10290 21480
rect 10870 21428 10876 21480
rect 10928 21468 10934 21480
rect 11532 21477 11560 21508
rect 13262 21496 13268 21548
rect 13320 21536 13326 21548
rect 14660 21536 14688 21576
rect 14918 21536 14924 21548
rect 13320 21508 13584 21536
rect 13320 21496 13326 21508
rect 11241 21471 11299 21477
rect 11241 21468 11253 21471
rect 10928 21440 11253 21468
rect 10928 21428 10934 21440
rect 11241 21437 11253 21440
rect 11287 21437 11299 21471
rect 11241 21431 11299 21437
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21468 11575 21471
rect 11698 21468 11704 21480
rect 11563 21440 11704 21468
rect 11563 21437 11575 21440
rect 11517 21431 11575 21437
rect 11698 21428 11704 21440
rect 11756 21428 11762 21480
rect 12894 21428 12900 21480
rect 12952 21468 12958 21480
rect 12989 21471 13047 21477
rect 12989 21468 13001 21471
rect 12952 21440 13001 21468
rect 12952 21428 12958 21440
rect 12989 21437 13001 21440
rect 13035 21437 13047 21471
rect 12989 21431 13047 21437
rect 13173 21471 13231 21477
rect 13173 21437 13185 21471
rect 13219 21468 13231 21471
rect 13354 21468 13360 21480
rect 13219 21440 13360 21468
rect 13219 21437 13231 21440
rect 13173 21431 13231 21437
rect 13354 21428 13360 21440
rect 13412 21428 13418 21480
rect 13556 21477 13584 21508
rect 13740 21508 14688 21536
rect 14879 21508 14924 21536
rect 13541 21471 13599 21477
rect 13541 21437 13553 21471
rect 13587 21437 13599 21471
rect 13541 21431 13599 21437
rect 2406 21400 2412 21412
rect 1780 21372 2412 21400
rect 2406 21360 2412 21372
rect 2464 21360 2470 21412
rect 4890 21400 4896 21412
rect 3160 21372 4896 21400
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 3160 21341 3188 21372
rect 4890 21360 4896 21372
rect 4948 21360 4954 21412
rect 9033 21403 9091 21409
rect 9033 21369 9045 21403
rect 9079 21400 9091 21403
rect 9122 21400 9128 21412
rect 9079 21372 9128 21400
rect 9079 21369 9091 21372
rect 9033 21363 9091 21369
rect 9122 21360 9128 21372
rect 9180 21360 9186 21412
rect 9249 21403 9307 21409
rect 9249 21369 9261 21403
rect 9295 21400 9307 21403
rect 9858 21400 9864 21412
rect 9295 21372 9864 21400
rect 9295 21369 9307 21372
rect 9249 21363 9307 21369
rect 9858 21360 9864 21372
rect 9916 21360 9922 21412
rect 10244 21400 10272 21428
rect 12158 21400 12164 21412
rect 10244 21372 12164 21400
rect 12158 21360 12164 21372
rect 12216 21360 12222 21412
rect 13449 21403 13507 21409
rect 13449 21369 13461 21403
rect 13495 21400 13507 21403
rect 13630 21400 13636 21412
rect 13495 21372 13636 21400
rect 13495 21369 13507 21372
rect 13449 21363 13507 21369
rect 13630 21360 13636 21372
rect 13688 21360 13694 21412
rect 3145 21335 3203 21341
rect 3145 21332 3157 21335
rect 3108 21304 3157 21332
rect 3108 21292 3114 21304
rect 3145 21301 3157 21304
rect 3191 21301 3203 21335
rect 3145 21295 3203 21301
rect 3326 21292 3332 21344
rect 3384 21332 3390 21344
rect 3878 21332 3884 21344
rect 3384 21304 3884 21332
rect 3384 21292 3390 21304
rect 3878 21292 3884 21304
rect 3936 21292 3942 21344
rect 4249 21335 4307 21341
rect 4249 21301 4261 21335
rect 4295 21332 4307 21335
rect 4614 21332 4620 21344
rect 4295 21304 4620 21332
rect 4295 21301 4307 21304
rect 4249 21295 4307 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 6549 21335 6607 21341
rect 6549 21301 6561 21335
rect 6595 21332 6607 21335
rect 7190 21332 7196 21344
rect 6595 21304 7196 21332
rect 6595 21301 6607 21304
rect 6549 21295 6607 21301
rect 7190 21292 7196 21304
rect 7248 21332 7254 21344
rect 7650 21332 7656 21344
rect 7248 21304 7656 21332
rect 7248 21292 7254 21304
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 8386 21332 8392 21344
rect 8347 21304 8392 21332
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 13078 21292 13084 21344
rect 13136 21332 13142 21344
rect 13262 21332 13268 21344
rect 13136 21304 13268 21332
rect 13136 21292 13142 21304
rect 13262 21292 13268 21304
rect 13320 21332 13326 21344
rect 13740 21332 13768 21508
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 15378 21536 15384 21548
rect 15212 21508 15384 21536
rect 14366 21428 14372 21480
rect 14424 21468 14430 21480
rect 15010 21477 15016 21480
rect 14645 21471 14703 21477
rect 14645 21468 14657 21471
rect 14424 21440 14657 21468
rect 14424 21428 14430 21440
rect 14645 21437 14657 21440
rect 14691 21437 14703 21471
rect 14645 21431 14703 21437
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21437 14887 21471
rect 15009 21468 15016 21477
rect 14971 21440 15016 21468
rect 14829 21431 14887 21437
rect 15009 21431 15016 21440
rect 14844 21400 14872 21431
rect 15010 21428 15016 21431
rect 15068 21428 15074 21480
rect 15212 21479 15240 21508
rect 15378 21496 15384 21508
rect 15436 21536 15442 21548
rect 15562 21536 15568 21548
rect 15436 21508 15568 21536
rect 15436 21496 15442 21508
rect 15562 21496 15568 21508
rect 15620 21496 15626 21548
rect 15672 21536 15700 21576
rect 15672 21508 15884 21536
rect 15197 21473 15255 21479
rect 15197 21439 15209 21473
rect 15243 21439 15255 21473
rect 15197 21433 15255 21439
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 15746 21468 15752 21480
rect 15528 21440 15752 21468
rect 15528 21428 15534 21440
rect 15746 21428 15752 21440
rect 15804 21428 15810 21480
rect 15856 21468 15884 21508
rect 17678 21496 17684 21548
rect 17736 21536 17742 21548
rect 18322 21536 18328 21548
rect 17736 21508 18328 21536
rect 17736 21496 17742 21508
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 18782 21496 18788 21548
rect 18840 21536 18846 21548
rect 19904 21545 19932 21576
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 20088 21604 20116 21644
rect 21269 21641 21281 21675
rect 21315 21672 21327 21675
rect 21450 21672 21456 21684
rect 21315 21644 21456 21672
rect 21315 21641 21327 21644
rect 21269 21635 21327 21641
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22281 21675 22339 21681
rect 22281 21672 22293 21675
rect 22244 21644 22293 21672
rect 22244 21632 22250 21644
rect 22281 21641 22293 21644
rect 22327 21672 22339 21675
rect 22462 21672 22468 21684
rect 22327 21644 22468 21672
rect 22327 21641 22339 21644
rect 22281 21635 22339 21641
rect 22462 21632 22468 21644
rect 22520 21632 22526 21684
rect 23109 21675 23167 21681
rect 23109 21641 23121 21675
rect 23155 21672 23167 21675
rect 23934 21672 23940 21684
rect 23155 21644 23940 21672
rect 23155 21641 23167 21644
rect 23109 21635 23167 21641
rect 23934 21632 23940 21644
rect 23992 21632 23998 21684
rect 24394 21672 24400 21684
rect 24355 21644 24400 21672
rect 24394 21632 24400 21644
rect 24452 21632 24458 21684
rect 25314 21672 25320 21684
rect 24504 21644 25320 21672
rect 23753 21607 23811 21613
rect 20088 21576 22094 21604
rect 22066 21548 22094 21576
rect 23753 21573 23765 21607
rect 23799 21604 23811 21607
rect 24504 21604 24532 21644
rect 25314 21632 25320 21644
rect 25372 21632 25378 21684
rect 27522 21632 27528 21684
rect 27580 21672 27586 21684
rect 27580 21644 28764 21672
rect 27580 21632 27586 21644
rect 24946 21604 24952 21616
rect 23799 21576 24532 21604
rect 24596 21576 24952 21604
rect 23799 21573 23811 21576
rect 23753 21567 23811 21573
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 18840 21508 19809 21536
rect 18840 21496 18846 21508
rect 19797 21505 19809 21508
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21505 19947 21539
rect 21082 21536 21088 21548
rect 19889 21499 19947 21505
rect 20088 21508 21088 21536
rect 16390 21468 16396 21480
rect 15856 21440 16396 21468
rect 16390 21428 16396 21440
rect 16448 21428 16454 21480
rect 16574 21428 16580 21480
rect 16632 21468 16638 21480
rect 17865 21471 17923 21477
rect 16632 21440 17816 21468
rect 16632 21428 16638 21440
rect 16016 21403 16074 21409
rect 14844 21372 14918 21400
rect 13320 21304 13768 21332
rect 13320 21292 13326 21304
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 14890 21332 14918 21372
rect 16016 21369 16028 21403
rect 16062 21400 16074 21403
rect 16850 21400 16856 21412
rect 16062 21372 16856 21400
rect 16062 21369 16074 21372
rect 16016 21363 16074 21369
rect 16850 21360 16856 21372
rect 16908 21360 16914 21412
rect 15654 21332 15660 21344
rect 14516 21304 15660 21332
rect 14516 21292 14522 21304
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 17126 21332 17132 21344
rect 17000 21304 17132 21332
rect 17000 21292 17006 21304
rect 17126 21292 17132 21304
rect 17184 21292 17190 21344
rect 17788 21332 17816 21440
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 18598 21468 18604 21480
rect 17911 21440 18604 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 18598 21428 18604 21440
rect 18656 21468 18662 21480
rect 19613 21471 19671 21477
rect 19613 21468 19625 21471
rect 18656 21440 19625 21468
rect 18656 21428 18662 21440
rect 19613 21437 19625 21440
rect 19659 21468 19671 21471
rect 19702 21468 19708 21480
rect 19659 21440 19708 21468
rect 19659 21437 19671 21440
rect 19613 21431 19671 21437
rect 19702 21428 19708 21440
rect 19760 21428 19766 21480
rect 19981 21471 20039 21477
rect 19981 21437 19993 21471
rect 20027 21468 20039 21471
rect 20088 21468 20116 21508
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 22066 21508 22100 21548
rect 22094 21496 22100 21508
rect 22152 21536 22158 21548
rect 24394 21536 24400 21548
rect 22152 21508 24400 21536
rect 22152 21496 22158 21508
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 20027 21440 20116 21468
rect 23201 21471 23259 21477
rect 20165 21449 20223 21455
rect 20027 21437 20039 21440
rect 19981 21431 20039 21437
rect 20165 21415 20177 21449
rect 20211 21415 20223 21449
rect 23201 21437 23213 21471
rect 23247 21437 23259 21471
rect 23658 21468 23664 21480
rect 23619 21440 23664 21468
rect 23201 21431 23259 21437
rect 20165 21412 20223 21415
rect 18506 21400 18512 21412
rect 18467 21372 18512 21400
rect 18506 21360 18512 21372
rect 18564 21360 18570 21412
rect 19334 21360 19340 21412
rect 19392 21400 19398 21412
rect 20162 21400 20168 21412
rect 19392 21372 20168 21400
rect 19392 21360 19398 21372
rect 20162 21360 20168 21372
rect 20220 21360 20226 21412
rect 20254 21332 20260 21344
rect 17788 21304 20260 21332
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 20717 21335 20775 21341
rect 20717 21301 20729 21335
rect 20763 21332 20775 21335
rect 20806 21332 20812 21344
rect 20763 21304 20812 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 23216 21332 23244 21431
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 24596 21477 24624 21576
rect 24946 21564 24952 21576
rect 25004 21564 25010 21616
rect 25774 21564 25780 21616
rect 25832 21564 25838 21616
rect 28442 21604 28448 21616
rect 28368 21576 28448 21604
rect 24765 21539 24823 21545
rect 24765 21505 24777 21539
rect 24811 21536 24823 21539
rect 25792 21536 25820 21564
rect 28368 21545 28396 21576
rect 28442 21564 28448 21576
rect 28500 21564 28506 21616
rect 25961 21539 26019 21545
rect 25961 21536 25973 21539
rect 24811 21508 25973 21536
rect 24811 21505 24823 21508
rect 24765 21499 24823 21505
rect 25961 21505 25973 21508
rect 26007 21536 26019 21539
rect 27157 21539 27215 21545
rect 27157 21536 27169 21539
rect 26007 21508 27169 21536
rect 26007 21505 26019 21508
rect 25961 21499 26019 21505
rect 27157 21505 27169 21508
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21536 27307 21539
rect 28353 21539 28411 21545
rect 27295 21508 28304 21536
rect 27295 21505 27307 21508
rect 27249 21499 27307 21505
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21437 24639 21471
rect 24854 21468 24860 21480
rect 24767 21440 24860 21468
rect 24581 21431 24639 21437
rect 24854 21428 24860 21440
rect 24912 21428 24918 21480
rect 24946 21428 24952 21480
rect 25004 21468 25010 21480
rect 25004 21440 25049 21468
rect 25004 21428 25010 21440
rect 25130 21428 25136 21480
rect 25188 21468 25194 21480
rect 25593 21471 25651 21477
rect 25869 21471 25927 21477
rect 25593 21468 25605 21471
rect 25188 21440 25605 21468
rect 25188 21428 25194 21440
rect 25593 21437 25605 21440
rect 25639 21437 25651 21471
rect 25777 21465 25835 21471
rect 25777 21462 25789 21465
rect 25593 21431 25651 21437
rect 25720 21434 25789 21462
rect 23566 21360 23572 21412
rect 23624 21400 23630 21412
rect 24872 21400 24900 21428
rect 23624 21372 24900 21400
rect 23624 21360 23630 21372
rect 25498 21332 25504 21344
rect 23216 21304 25504 21332
rect 25498 21292 25504 21304
rect 25556 21332 25562 21344
rect 25720 21332 25748 21434
rect 25777 21431 25789 21434
rect 25823 21431 25835 21465
rect 25869 21437 25881 21471
rect 25915 21468 25927 21471
rect 26142 21468 26148 21480
rect 25915 21440 26004 21468
rect 26103 21440 26148 21468
rect 25915 21437 25927 21440
rect 25869 21431 25927 21437
rect 25777 21425 25835 21431
rect 25976 21400 26004 21440
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 26973 21471 27031 21477
rect 26973 21437 26985 21471
rect 27019 21437 27031 21471
rect 26973 21431 27031 21437
rect 27341 21471 27399 21477
rect 27341 21437 27353 21471
rect 27387 21437 27399 21471
rect 27522 21468 27528 21480
rect 27483 21440 27528 21468
rect 27341 21431 27399 21437
rect 26050 21400 26056 21412
rect 25976 21372 26056 21400
rect 26050 21360 26056 21372
rect 26108 21360 26114 21412
rect 26988 21400 27016 21431
rect 26226 21372 27016 21400
rect 27356 21400 27384 21431
rect 27522 21428 27528 21440
rect 27580 21428 27586 21480
rect 28166 21468 28172 21480
rect 28127 21440 28172 21468
rect 28166 21428 28172 21440
rect 28224 21428 28230 21480
rect 28276 21468 28304 21508
rect 28353 21505 28365 21539
rect 28399 21505 28411 21539
rect 28353 21499 28411 21505
rect 28442 21468 28448 21480
rect 28276 21440 28448 21468
rect 28442 21428 28448 21440
rect 28500 21428 28506 21480
rect 28534 21428 28540 21480
rect 28592 21468 28598 21480
rect 28736 21477 28764 21644
rect 29454 21632 29460 21684
rect 29512 21672 29518 21684
rect 31294 21672 31300 21684
rect 29512 21644 31300 21672
rect 29512 21632 29518 21644
rect 31294 21632 31300 21644
rect 31352 21632 31358 21684
rect 31018 21564 31024 21616
rect 31076 21604 31082 21616
rect 31113 21607 31171 21613
rect 31113 21604 31125 21607
rect 31076 21576 31125 21604
rect 31076 21564 31082 21576
rect 31113 21573 31125 21576
rect 31159 21573 31171 21607
rect 32324 21604 32352 21848
rect 31113 21567 31171 21573
rect 32232 21576 32352 21604
rect 30469 21539 30527 21545
rect 30469 21505 30481 21539
rect 30515 21536 30527 21539
rect 30650 21536 30656 21548
rect 30515 21508 30656 21536
rect 30515 21505 30527 21508
rect 30469 21499 30527 21505
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 31386 21496 31392 21548
rect 31444 21536 31450 21548
rect 31570 21536 31576 21548
rect 31444 21508 31576 21536
rect 31444 21496 31450 21508
rect 31570 21496 31576 21508
rect 31628 21496 31634 21548
rect 28721 21471 28779 21477
rect 28592 21440 28637 21468
rect 28592 21428 28598 21440
rect 28721 21437 28733 21471
rect 28767 21437 28779 21471
rect 28721 21431 28779 21437
rect 30561 21471 30619 21477
rect 30561 21437 30573 21471
rect 30607 21468 30619 21471
rect 30834 21468 30840 21480
rect 30607 21440 30840 21468
rect 30607 21437 30619 21440
rect 30561 21431 30619 21437
rect 30834 21428 30840 21440
rect 30892 21468 30898 21480
rect 31021 21471 31079 21477
rect 31021 21468 31033 21471
rect 30892 21440 31033 21468
rect 30892 21428 30898 21440
rect 31021 21437 31033 21440
rect 31067 21437 31079 21471
rect 31021 21431 31079 21437
rect 28184 21400 28212 21428
rect 30282 21400 30288 21412
rect 27356 21372 28212 21400
rect 30243 21372 30288 21400
rect 26226 21332 26254 21372
rect 30282 21360 30288 21372
rect 30340 21360 30346 21412
rect 31036 21400 31064 21431
rect 31202 21428 31208 21480
rect 31260 21468 31266 21480
rect 31297 21471 31355 21477
rect 31297 21468 31309 21471
rect 31260 21440 31309 21468
rect 31260 21428 31266 21440
rect 31297 21437 31309 21440
rect 31343 21437 31355 21471
rect 32232 21468 32260 21576
rect 32320 21468 33120 21482
rect 32232 21440 33120 21468
rect 31297 21431 31355 21437
rect 32320 21426 33120 21440
rect 31570 21400 31576 21412
rect 31036 21372 31576 21400
rect 31570 21360 31576 21372
rect 31628 21360 31634 21412
rect 26326 21332 26332 21344
rect 25556 21304 26254 21332
rect 26287 21304 26332 21332
rect 25556 21292 25562 21304
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 26602 21292 26608 21344
rect 26660 21332 26666 21344
rect 26789 21335 26847 21341
rect 26789 21332 26801 21335
rect 26660 21304 26801 21332
rect 26660 21292 26666 21304
rect 26789 21301 26801 21304
rect 26835 21301 26847 21335
rect 27982 21332 27988 21344
rect 27943 21304 27988 21332
rect 26789 21295 26847 21301
rect 27982 21292 27988 21304
rect 28040 21292 28046 21344
rect 28074 21292 28080 21344
rect 28132 21332 28138 21344
rect 29549 21335 29607 21341
rect 29549 21332 29561 21335
rect 28132 21304 29561 21332
rect 28132 21292 28138 21304
rect 29549 21301 29561 21304
rect 29595 21301 29607 21335
rect 29549 21295 29607 21301
rect 30466 21292 30472 21344
rect 30524 21332 30530 21344
rect 30561 21335 30619 21341
rect 30561 21332 30573 21335
rect 30524 21304 30573 21332
rect 30524 21292 30530 21304
rect 30561 21301 30573 21304
rect 30607 21301 30619 21335
rect 30561 21295 30619 21301
rect 31021 21335 31079 21341
rect 31021 21301 31033 21335
rect 31067 21332 31079 21335
rect 31202 21332 31208 21344
rect 31067 21304 31208 21332
rect 31067 21301 31079 21304
rect 31021 21295 31079 21301
rect 31202 21292 31208 21304
rect 31260 21292 31266 21344
rect 1104 21242 32016 21264
rect 1104 21190 11253 21242
rect 11305 21190 11317 21242
rect 11369 21190 11381 21242
rect 11433 21190 11445 21242
rect 11497 21190 11509 21242
rect 11561 21190 21557 21242
rect 21609 21190 21621 21242
rect 21673 21190 21685 21242
rect 21737 21190 21749 21242
rect 21801 21190 21813 21242
rect 21865 21190 32016 21242
rect 1104 21168 32016 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 5629 21131 5687 21137
rect 5629 21128 5641 21131
rect 3476 21100 5641 21128
rect 3476 21088 3482 21100
rect 5629 21097 5641 21100
rect 5675 21128 5687 21131
rect 6730 21128 6736 21140
rect 5675 21100 6736 21128
rect 5675 21097 5687 21100
rect 5629 21091 5687 21097
rect 6730 21088 6736 21100
rect 6788 21128 6794 21140
rect 7282 21128 7288 21140
rect 6788 21100 7288 21128
rect 6788 21088 6794 21100
rect 7282 21088 7288 21100
rect 7340 21088 7346 21140
rect 8294 21088 8300 21140
rect 8352 21128 8358 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8352 21100 8953 21128
rect 8352 21088 8358 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 9122 21088 9128 21140
rect 9180 21128 9186 21140
rect 9585 21131 9643 21137
rect 9585 21128 9597 21131
rect 9180 21100 9597 21128
rect 9180 21088 9186 21100
rect 9585 21097 9597 21100
rect 9631 21097 9643 21131
rect 12894 21128 12900 21140
rect 12855 21100 12900 21128
rect 9585 21091 9643 21097
rect 12894 21088 12900 21100
rect 12952 21088 12958 21140
rect 16574 21128 16580 21140
rect 14200 21100 16580 21128
rect 1854 21020 1860 21072
rect 1912 21060 1918 21072
rect 2682 21060 2688 21072
rect 1912 21032 2688 21060
rect 1912 21020 1918 21032
rect 2682 21020 2688 21032
rect 2740 21020 2746 21072
rect 3234 21060 3240 21072
rect 2884 21032 3240 21060
rect 1397 20995 1455 21001
rect 1397 20992 1409 20995
rect 1044 20964 1409 20992
rect 1397 20961 1409 20964
rect 1443 20961 1455 20995
rect 1397 20955 1455 20961
rect 2225 20995 2283 21001
rect 2225 20961 2237 20995
rect 2271 20992 2283 20995
rect 2406 20992 2412 21004
rect 2271 20964 2412 20992
rect 2271 20961 2283 20964
rect 2225 20955 2283 20961
rect 1412 20924 1440 20955
rect 2406 20952 2412 20964
rect 2464 20952 2470 21004
rect 2884 21001 2912 21032
rect 3234 21020 3240 21032
rect 3292 21060 3298 21072
rect 3605 21063 3663 21069
rect 3605 21060 3617 21063
rect 3292 21032 3617 21060
rect 3292 21020 3298 21032
rect 3605 21029 3617 21032
rect 3651 21029 3663 21063
rect 3605 21023 3663 21029
rect 3786 21020 3792 21072
rect 3844 21069 3850 21072
rect 3844 21063 3863 21069
rect 3851 21029 3863 21063
rect 3844 21023 3863 21029
rect 5721 21063 5779 21069
rect 5721 21029 5733 21063
rect 5767 21060 5779 21063
rect 5902 21060 5908 21072
rect 5767 21032 5908 21060
rect 5767 21029 5779 21032
rect 5721 21023 5779 21029
rect 3844 21020 3850 21023
rect 5902 21020 5908 21032
rect 5960 21060 5966 21072
rect 7006 21060 7012 21072
rect 5960 21032 7012 21060
rect 5960 21020 5966 21032
rect 7006 21020 7012 21032
rect 7064 21020 7070 21072
rect 10873 21063 10931 21069
rect 10873 21029 10885 21063
rect 10919 21060 10931 21063
rect 14200 21060 14228 21100
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 16758 21128 16764 21140
rect 16719 21100 16764 21128
rect 16758 21088 16764 21100
rect 16816 21088 16822 21140
rect 18138 21088 18144 21140
rect 18196 21128 18202 21140
rect 21910 21128 21916 21140
rect 18196 21100 21916 21128
rect 18196 21088 18202 21100
rect 21910 21088 21916 21100
rect 21968 21088 21974 21140
rect 22112 21100 23520 21128
rect 14918 21060 14924 21072
rect 10919 21032 11744 21060
rect 10919 21029 10931 21032
rect 10873 21023 10931 21029
rect 2869 20995 2927 21001
rect 2869 20961 2881 20995
rect 2915 20961 2927 20995
rect 3510 20992 3516 21004
rect 2869 20955 2927 20961
rect 2976 20964 3516 20992
rect 2976 20924 3004 20964
rect 3510 20952 3516 20964
rect 3568 20952 3574 21004
rect 3620 20964 4476 20992
rect 3142 20924 3148 20936
rect 1412 20896 3004 20924
rect 3103 20896 3148 20924
rect 3142 20884 3148 20896
rect 3200 20884 3206 20936
rect 3326 20884 3332 20936
rect 3384 20924 3390 20936
rect 3620 20924 3648 20964
rect 3384 20896 3648 20924
rect 3384 20884 3390 20896
rect 3878 20884 3884 20936
rect 3936 20924 3942 20936
rect 4062 20924 4068 20936
rect 3936 20896 4068 20924
rect 3936 20884 3942 20896
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4448 20924 4476 20964
rect 4522 20952 4528 21004
rect 4580 20992 4586 21004
rect 4617 20995 4675 21001
rect 4617 20992 4629 20995
rect 4580 20964 4629 20992
rect 4580 20952 4586 20964
rect 4617 20961 4629 20964
rect 4663 20961 4675 20995
rect 4617 20955 4675 20961
rect 5994 20952 6000 21004
rect 6052 20992 6058 21004
rect 7193 20995 7251 21001
rect 7193 20992 7205 20995
rect 6052 20964 7205 20992
rect 6052 20952 6058 20964
rect 7193 20961 7205 20964
rect 7239 20961 7251 20995
rect 7193 20955 7251 20961
rect 8018 20952 8024 21004
rect 8076 20992 8082 21004
rect 8205 20995 8263 21001
rect 8205 20992 8217 20995
rect 8076 20964 8217 20992
rect 8076 20952 8082 20964
rect 8205 20961 8217 20964
rect 8251 20961 8263 20995
rect 8386 20992 8392 21004
rect 8299 20964 8392 20992
rect 8205 20955 8263 20961
rect 8386 20952 8392 20964
rect 8444 20992 8450 21004
rect 8938 20992 8944 21004
rect 8444 20964 8944 20992
rect 8444 20952 8450 20964
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9766 20992 9772 21004
rect 9723 20964 9772 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 10789 20995 10847 21001
rect 10789 20961 10801 20995
rect 10835 20992 10847 20995
rect 10962 20992 10968 21004
rect 10835 20964 10968 20992
rect 10835 20961 10847 20964
rect 10789 20955 10847 20961
rect 10962 20952 10968 20964
rect 11020 20992 11026 21004
rect 11146 20992 11152 21004
rect 11020 20964 11152 20992
rect 11020 20952 11026 20964
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 11514 20992 11520 21004
rect 11475 20964 11520 20992
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 11716 21001 11744 21032
rect 11808 21032 14228 21060
rect 14568 21032 14924 21060
rect 11808 21001 11836 21032
rect 11701 20995 11759 21001
rect 11701 20961 11713 20995
rect 11747 20961 11759 20995
rect 11701 20955 11759 20961
rect 11793 20995 11851 21001
rect 11793 20961 11805 20995
rect 11839 20961 11851 20995
rect 11793 20955 11851 20961
rect 12069 20995 12127 21001
rect 12069 20961 12081 20995
rect 12115 20992 12127 20995
rect 12434 20992 12440 21004
rect 12115 20964 12440 20992
rect 12115 20961 12127 20964
rect 12069 20955 12127 20961
rect 12434 20952 12440 20964
rect 12492 20952 12498 21004
rect 13078 20992 13084 21004
rect 13039 20964 13084 20992
rect 13078 20952 13084 20964
rect 13136 20952 13142 21004
rect 13262 20992 13268 21004
rect 13223 20964 13268 20992
rect 13262 20952 13268 20964
rect 13320 20952 13326 21004
rect 13446 20992 13452 21004
rect 13407 20964 13452 20992
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 13633 20995 13691 21001
rect 13633 20961 13645 20995
rect 13679 20961 13691 20995
rect 14274 20992 14280 21004
rect 14235 20964 14280 20992
rect 13633 20955 13691 20961
rect 4706 20924 4712 20936
rect 4448 20896 4712 20924
rect 4706 20884 4712 20896
rect 4764 20884 4770 20936
rect 5166 20884 5172 20936
rect 5224 20924 5230 20936
rect 5902 20924 5908 20936
rect 5224 20896 5908 20924
rect 5224 20884 5230 20896
rect 5902 20884 5908 20896
rect 5960 20884 5966 20936
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20924 6515 20927
rect 6917 20927 6975 20933
rect 6917 20924 6929 20927
rect 6503 20896 6929 20924
rect 6503 20893 6515 20896
rect 6457 20887 6515 20893
rect 6917 20893 6929 20896
rect 6963 20924 6975 20927
rect 9214 20924 9220 20936
rect 6963 20896 9220 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 9214 20884 9220 20896
rect 9272 20884 9278 20936
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20924 11943 20927
rect 11974 20924 11980 20936
rect 11931 20896 11980 20924
rect 11931 20893 11943 20896
rect 11885 20887 11943 20893
rect 1394 20816 1400 20868
rect 1452 20856 1458 20868
rect 1581 20859 1639 20865
rect 1581 20856 1593 20859
rect 1452 20828 1593 20856
rect 1452 20816 1458 20828
rect 1581 20825 1593 20828
rect 1627 20856 1639 20859
rect 2774 20856 2780 20868
rect 1627 20828 2780 20856
rect 1627 20825 1639 20828
rect 1581 20819 1639 20825
rect 2774 20816 2780 20828
rect 2832 20816 2838 20868
rect 3053 20859 3111 20865
rect 3053 20825 3065 20859
rect 3099 20856 3111 20859
rect 4890 20856 4896 20868
rect 3099 20828 4896 20856
rect 3099 20825 3111 20828
rect 3053 20819 3111 20825
rect 4890 20816 4896 20828
rect 4948 20816 4954 20868
rect 9950 20816 9956 20868
rect 10008 20856 10014 20868
rect 11900 20856 11928 20887
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 13357 20927 13415 20933
rect 13357 20893 13369 20927
rect 13403 20924 13415 20927
rect 13538 20924 13544 20936
rect 13403 20896 13544 20924
rect 13403 20893 13415 20896
rect 13357 20887 13415 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 10008 20828 11928 20856
rect 10008 20816 10014 20828
rect 12986 20816 12992 20868
rect 13044 20856 13050 20868
rect 13648 20856 13676 20955
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 14458 20992 14464 21004
rect 14419 20964 14464 20992
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 14568 21001 14596 21032
rect 14918 21020 14924 21032
rect 14976 21020 14982 21072
rect 15010 21020 15016 21072
rect 15068 21060 15074 21072
rect 15068 21032 16712 21060
rect 15068 21020 15074 21032
rect 14553 20995 14611 21001
rect 14553 20961 14565 20995
rect 14599 20961 14611 20995
rect 14553 20955 14611 20961
rect 14645 20995 14703 21001
rect 14645 20961 14657 20995
rect 14691 20961 14703 20995
rect 14645 20955 14703 20961
rect 14829 20995 14887 21001
rect 14829 20961 14841 20995
rect 14875 20992 14887 20995
rect 15378 20992 15384 21004
rect 14875 20964 15384 20992
rect 14875 20961 14887 20964
rect 14829 20955 14887 20961
rect 14660 20924 14688 20955
rect 15378 20952 15384 20964
rect 15436 20992 15442 21004
rect 15930 20992 15936 21004
rect 15436 20964 15936 20992
rect 15436 20952 15442 20964
rect 15930 20952 15936 20964
rect 15988 20952 15994 21004
rect 16684 21001 16712 21032
rect 17310 21020 17316 21072
rect 17368 21060 17374 21072
rect 17368 21032 21036 21060
rect 17368 21020 17374 21032
rect 16669 20995 16727 21001
rect 16669 20961 16681 20995
rect 16715 20961 16727 20995
rect 16669 20955 16727 20961
rect 16758 20952 16764 21004
rect 16816 20992 16822 21004
rect 17402 20992 17408 21004
rect 16816 20964 17408 20992
rect 16816 20952 16822 20964
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 17957 20995 18015 21001
rect 17957 20961 17969 20995
rect 18003 20992 18015 20995
rect 18598 20992 18604 21004
rect 18003 20964 18604 20992
rect 18003 20961 18015 20964
rect 17957 20955 18015 20961
rect 18598 20952 18604 20964
rect 18656 20952 18662 21004
rect 18782 20952 18788 21004
rect 18840 20992 18846 21004
rect 18969 20995 19027 21001
rect 18969 20992 18981 20995
rect 18840 20964 18981 20992
rect 18840 20952 18846 20964
rect 18969 20961 18981 20964
rect 19015 20992 19027 20995
rect 20898 20992 20904 21004
rect 19015 20964 20904 20992
rect 19015 20961 19027 20964
rect 18969 20955 19027 20961
rect 20898 20952 20904 20964
rect 20956 20952 20962 21004
rect 15562 20924 15568 20936
rect 14660 20896 15568 20924
rect 15562 20884 15568 20896
rect 15620 20884 15626 20936
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 15838 20924 15844 20936
rect 15712 20896 15844 20924
rect 15712 20884 15718 20896
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 16114 20924 16120 20936
rect 16075 20896 16120 20924
rect 16114 20884 16120 20896
rect 16172 20884 16178 20936
rect 16206 20884 16212 20936
rect 16264 20924 16270 20936
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 16264 20896 18245 20924
rect 16264 20884 16270 20896
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 13044 20828 13676 20856
rect 13740 20828 15792 20856
rect 13044 20816 13050 20828
rect 2314 20788 2320 20800
rect 2275 20760 2320 20788
rect 2314 20748 2320 20760
rect 2372 20748 2378 20800
rect 2958 20788 2964 20800
rect 2871 20760 2964 20788
rect 2958 20748 2964 20760
rect 3016 20788 3022 20800
rect 3326 20788 3332 20800
rect 3016 20760 3332 20788
rect 3016 20748 3022 20760
rect 3326 20748 3332 20760
rect 3384 20748 3390 20800
rect 3789 20791 3847 20797
rect 3789 20757 3801 20791
rect 3835 20788 3847 20791
rect 3878 20788 3884 20800
rect 3835 20760 3884 20788
rect 3835 20757 3847 20760
rect 3789 20751 3847 20757
rect 3878 20748 3884 20760
rect 3936 20748 3942 20800
rect 3973 20791 4031 20797
rect 3973 20757 3985 20791
rect 4019 20788 4031 20791
rect 4154 20788 4160 20800
rect 4019 20760 4160 20788
rect 4019 20757 4031 20760
rect 3973 20751 4031 20757
rect 4154 20748 4160 20760
rect 4212 20748 4218 20800
rect 4430 20748 4436 20800
rect 4488 20788 4494 20800
rect 4525 20791 4583 20797
rect 4525 20788 4537 20791
rect 4488 20760 4537 20788
rect 4488 20748 4494 20760
rect 4525 20757 4537 20760
rect 4571 20757 4583 20791
rect 4525 20751 4583 20757
rect 10321 20791 10379 20797
rect 10321 20757 10333 20791
rect 10367 20788 10379 20791
rect 10870 20788 10876 20800
rect 10367 20760 10876 20788
rect 10367 20757 10379 20760
rect 10321 20751 10379 20757
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 11974 20748 11980 20800
rect 12032 20788 12038 20800
rect 12253 20791 12311 20797
rect 12253 20788 12265 20791
rect 12032 20760 12265 20788
rect 12032 20748 12038 20760
rect 12253 20757 12265 20760
rect 12299 20757 12311 20791
rect 12253 20751 12311 20757
rect 13538 20748 13544 20800
rect 13596 20788 13602 20800
rect 13740 20788 13768 20828
rect 13596 20760 13768 20788
rect 14093 20791 14151 20797
rect 13596 20748 13602 20760
rect 14093 20757 14105 20791
rect 14139 20788 14151 20791
rect 14366 20788 14372 20800
rect 14139 20760 14372 20788
rect 14139 20757 14151 20760
rect 14093 20751 14151 20757
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 15102 20748 15108 20800
rect 15160 20788 15166 20800
rect 15654 20788 15660 20800
rect 15160 20760 15660 20788
rect 15160 20748 15166 20760
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 15764 20788 15792 20828
rect 16390 20816 16396 20868
rect 16448 20856 16454 20868
rect 18248 20856 18276 20887
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18564 20896 18705 20924
rect 18564 20884 18570 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20070 20924 20076 20936
rect 20027 20896 20076 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 19996 20856 20024 20887
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 20162 20884 20168 20936
rect 20220 20924 20226 20936
rect 20257 20927 20315 20933
rect 20257 20924 20269 20927
rect 20220 20896 20269 20924
rect 20220 20884 20226 20896
rect 20257 20893 20269 20896
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 16448 20828 17632 20856
rect 18248 20828 20024 20856
rect 21008 20856 21036 21032
rect 21358 21020 21364 21072
rect 21416 21060 21422 21072
rect 22112 21069 22140 21100
rect 22005 21063 22063 21069
rect 22005 21060 22017 21063
rect 21416 21032 22017 21060
rect 21416 21020 21422 21032
rect 22005 21029 22017 21032
rect 22051 21029 22063 21063
rect 22005 21023 22063 21029
rect 22097 21063 22155 21069
rect 22097 21029 22109 21063
rect 22143 21029 22155 21063
rect 22097 21023 22155 21029
rect 23106 21020 23112 21072
rect 23164 21060 23170 21072
rect 23492 21060 23520 21100
rect 23842 21088 23848 21140
rect 23900 21128 23906 21140
rect 25130 21128 25136 21140
rect 23900 21100 25136 21128
rect 23900 21088 23906 21100
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 25866 21088 25872 21140
rect 25924 21128 25930 21140
rect 25924 21100 26096 21128
rect 25924 21088 25930 21100
rect 23658 21060 23664 21072
rect 23164 21032 23428 21060
rect 23492 21032 23664 21060
rect 23164 21020 23170 21032
rect 22373 20995 22431 21001
rect 22373 20961 22385 20995
rect 22419 20992 22431 20995
rect 22554 20992 22560 21004
rect 22419 20964 22560 20992
rect 22419 20961 22431 20964
rect 22373 20955 22431 20961
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 23290 20992 23296 21004
rect 23247 20964 23296 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 23290 20952 23296 20964
rect 23348 20952 23354 21004
rect 23400 20992 23428 21032
rect 23658 21020 23664 21032
rect 23716 21060 23722 21072
rect 25958 21060 25964 21072
rect 23716 21032 25964 21060
rect 23716 21020 23722 21032
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 26068 21060 26096 21100
rect 28534 21088 28540 21140
rect 28592 21128 28598 21140
rect 28629 21131 28687 21137
rect 28629 21128 28641 21131
rect 28592 21100 28641 21128
rect 28592 21088 28598 21100
rect 28629 21097 28641 21100
rect 28675 21097 28687 21131
rect 29546 21128 29552 21140
rect 28629 21091 28687 21097
rect 28736 21100 29552 21128
rect 28736 21060 28764 21100
rect 29546 21088 29552 21100
rect 29604 21088 29610 21140
rect 30742 21128 30748 21140
rect 30703 21100 30748 21128
rect 30742 21088 30748 21100
rect 30800 21088 30806 21140
rect 26068 21032 28764 21060
rect 28810 21020 28816 21072
rect 28868 21060 28874 21072
rect 29742 21063 29800 21069
rect 29742 21060 29754 21063
rect 28868 21032 29754 21060
rect 28868 21020 28874 21032
rect 29742 21029 29754 21032
rect 29788 21029 29800 21063
rect 29742 21023 29800 21029
rect 23457 20995 23515 21001
rect 23457 20992 23469 20995
rect 23400 20964 23469 20992
rect 23457 20961 23469 20964
rect 23503 20961 23515 20995
rect 23457 20955 23515 20961
rect 24026 20952 24032 21004
rect 24084 20992 24090 21004
rect 24302 20992 24308 21004
rect 24084 20964 24308 20992
rect 24084 20952 24090 20964
rect 24302 20952 24308 20964
rect 24360 20952 24366 21004
rect 24762 20952 24768 21004
rect 24820 20992 24826 21004
rect 25774 20992 25780 21004
rect 24820 20964 25780 20992
rect 24820 20952 24826 20964
rect 25774 20952 25780 20964
rect 25832 20992 25838 21004
rect 25869 20995 25927 21001
rect 25869 20992 25881 20995
rect 25832 20964 25881 20992
rect 25832 20952 25838 20964
rect 25869 20961 25881 20964
rect 25915 20961 25927 20995
rect 25869 20955 25927 20961
rect 27893 20995 27951 21001
rect 27893 20961 27905 20995
rect 27939 20992 27951 20995
rect 28350 20992 28356 21004
rect 27939 20964 28356 20992
rect 27939 20961 27951 20964
rect 27893 20955 27951 20961
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 31018 20992 31024 21004
rect 30979 20964 31024 20992
rect 31018 20952 31024 20964
rect 31076 20952 31082 21004
rect 31202 20992 31208 21004
rect 31163 20964 31208 20992
rect 31202 20952 31208 20964
rect 31260 20952 31266 21004
rect 22462 20924 22468 20936
rect 22423 20896 22468 20924
rect 22462 20884 22468 20896
rect 22520 20884 22526 20936
rect 25590 20924 25596 20936
rect 25551 20896 25596 20924
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 28074 20884 28080 20936
rect 28132 20924 28138 20936
rect 28169 20927 28227 20933
rect 28169 20924 28181 20927
rect 28132 20896 28181 20924
rect 28132 20884 28138 20896
rect 28169 20893 28181 20896
rect 28215 20893 28227 20927
rect 28169 20887 28227 20893
rect 30009 20927 30067 20933
rect 30009 20893 30021 20927
rect 30055 20924 30067 20927
rect 30374 20924 30380 20936
rect 30055 20896 30380 20924
rect 30055 20893 30067 20896
rect 30009 20887 30067 20893
rect 30374 20884 30380 20896
rect 30432 20924 30438 20936
rect 30834 20924 30840 20936
rect 30432 20896 30840 20924
rect 30432 20884 30438 20896
rect 30834 20884 30840 20896
rect 30892 20884 30898 20936
rect 30926 20884 30932 20936
rect 30984 20924 30990 20936
rect 30984 20896 31029 20924
rect 30984 20884 30990 20896
rect 31110 20884 31116 20936
rect 31168 20924 31174 20936
rect 31168 20896 31213 20924
rect 31168 20884 31174 20896
rect 22922 20856 22928 20868
rect 21008 20828 22928 20856
rect 16448 20816 16454 20828
rect 17310 20788 17316 20800
rect 15764 20760 17316 20788
rect 17310 20748 17316 20760
rect 17368 20748 17374 20800
rect 17604 20788 17632 20828
rect 22922 20816 22928 20828
rect 22980 20816 22986 20868
rect 19150 20788 19156 20800
rect 17604 20760 19156 20788
rect 19150 20748 19156 20760
rect 19208 20748 19214 20800
rect 19794 20748 19800 20800
rect 19852 20788 19858 20800
rect 24118 20788 24124 20800
rect 19852 20760 24124 20788
rect 19852 20748 19858 20760
rect 24118 20748 24124 20760
rect 24176 20748 24182 20800
rect 24578 20788 24584 20800
rect 24539 20760 24584 20788
rect 24578 20748 24584 20760
rect 24636 20788 24642 20800
rect 24946 20788 24952 20800
rect 24636 20760 24952 20788
rect 24636 20748 24642 20760
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 25130 20748 25136 20800
rect 25188 20788 25194 20800
rect 27154 20788 27160 20800
rect 25188 20760 27160 20788
rect 25188 20748 25194 20760
rect 27154 20748 27160 20760
rect 27212 20748 27218 20800
rect 1104 20698 32016 20720
rect 1104 20646 6102 20698
rect 6154 20646 6166 20698
rect 6218 20646 6230 20698
rect 6282 20646 6294 20698
rect 6346 20646 6358 20698
rect 6410 20646 16405 20698
rect 16457 20646 16469 20698
rect 16521 20646 16533 20698
rect 16585 20646 16597 20698
rect 16649 20646 16661 20698
rect 16713 20646 26709 20698
rect 26761 20646 26773 20698
rect 26825 20646 26837 20698
rect 26889 20646 26901 20698
rect 26953 20646 26965 20698
rect 27017 20646 32016 20698
rect 1104 20624 32016 20646
rect 7650 20584 7656 20596
rect 2746 20556 7656 20584
rect 2746 20528 2774 20556
rect 7650 20544 7656 20556
rect 7708 20584 7714 20596
rect 8846 20584 8852 20596
rect 7708 20556 8852 20584
rect 7708 20544 7714 20556
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13173 20587 13231 20593
rect 13173 20584 13185 20587
rect 13136 20556 13185 20584
rect 13136 20544 13142 20556
rect 13173 20553 13185 20556
rect 13219 20553 13231 20587
rect 13354 20584 13360 20596
rect 13315 20556 13360 20584
rect 13173 20547 13231 20553
rect 2682 20476 2688 20528
rect 2740 20488 2774 20528
rect 3145 20519 3203 20525
rect 2740 20476 2746 20488
rect 3145 20485 3157 20519
rect 3191 20516 3203 20519
rect 5166 20516 5172 20528
rect 3191 20488 5172 20516
rect 3191 20485 3203 20488
rect 3145 20479 3203 20485
rect 5166 20476 5172 20488
rect 5224 20476 5230 20528
rect 5261 20519 5319 20525
rect 5261 20485 5273 20519
rect 5307 20516 5319 20519
rect 9950 20516 9956 20528
rect 5307 20488 9956 20516
rect 5307 20485 5319 20488
rect 5261 20479 5319 20485
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 10962 20476 10968 20528
rect 11020 20516 11026 20528
rect 11146 20516 11152 20528
rect 11020 20488 11152 20516
rect 11020 20476 11026 20488
rect 11146 20476 11152 20488
rect 11204 20516 11210 20528
rect 13188 20516 13216 20547
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 15010 20544 15016 20596
rect 15068 20584 15074 20596
rect 16669 20587 16727 20593
rect 15068 20556 16436 20584
rect 15068 20544 15074 20556
rect 16298 20516 16304 20528
rect 11204 20488 12020 20516
rect 13188 20488 13400 20516
rect 11204 20476 11210 20488
rect 2958 20448 2964 20460
rect 2919 20420 2964 20448
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 4430 20448 4436 20460
rect 4391 20420 4436 20448
rect 4430 20408 4436 20420
rect 4488 20408 4494 20460
rect 5810 20408 5816 20460
rect 5868 20448 5874 20460
rect 5868 20420 6408 20448
rect 5868 20408 5874 20420
rect 2038 20340 2044 20392
rect 2096 20380 2102 20392
rect 2317 20383 2375 20389
rect 2317 20380 2329 20383
rect 2096 20352 2329 20380
rect 2096 20340 2102 20352
rect 2317 20349 2329 20352
rect 2363 20349 2375 20383
rect 2317 20343 2375 20349
rect 2406 20340 2412 20392
rect 2464 20380 2470 20392
rect 2501 20383 2559 20389
rect 2501 20380 2513 20383
rect 2464 20352 2513 20380
rect 2464 20340 2470 20352
rect 2501 20349 2513 20352
rect 2547 20349 2559 20383
rect 2501 20343 2559 20349
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 4246 20380 4252 20392
rect 3292 20352 3337 20380
rect 4207 20352 4252 20380
rect 3292 20340 3298 20352
rect 4246 20340 4252 20352
rect 4304 20340 4310 20392
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20349 4583 20383
rect 4890 20380 4896 20392
rect 4851 20352 4896 20380
rect 4525 20343 4583 20349
rect 2961 20315 3019 20321
rect 2961 20281 2973 20315
rect 3007 20312 3019 20315
rect 4540 20312 4568 20343
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 6380 20389 6408 20420
rect 7558 20408 7564 20460
rect 7616 20448 7622 20460
rect 8202 20448 8208 20460
rect 7616 20420 8064 20448
rect 8163 20420 8208 20448
rect 7616 20408 7622 20420
rect 5905 20383 5963 20389
rect 5905 20380 5917 20383
rect 5500 20352 5917 20380
rect 5500 20340 5506 20352
rect 5905 20349 5917 20352
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 6365 20383 6423 20389
rect 6365 20349 6377 20383
rect 6411 20380 6423 20383
rect 6546 20380 6552 20392
rect 6411 20352 6552 20380
rect 6411 20349 6423 20352
rect 6365 20343 6423 20349
rect 6546 20340 6552 20352
rect 6604 20340 6610 20392
rect 7006 20380 7012 20392
rect 6967 20352 7012 20380
rect 7006 20340 7012 20352
rect 7064 20340 7070 20392
rect 7926 20380 7932 20392
rect 7887 20352 7932 20380
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8036 20389 8064 20420
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 11882 20448 11888 20460
rect 11843 20420 11888 20448
rect 11882 20408 11888 20420
rect 11940 20408 11946 20460
rect 11992 20448 12020 20488
rect 13372 20460 13400 20488
rect 16132 20488 16304 20516
rect 12434 20448 12440 20460
rect 11992 20420 12440 20448
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 8478 20380 8484 20392
rect 8067 20352 8484 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8478 20340 8484 20352
rect 8536 20340 8542 20392
rect 8938 20380 8944 20392
rect 8899 20352 8944 20380
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11054 20380 11060 20392
rect 11011 20352 11060 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11514 20340 11520 20392
rect 11572 20380 11578 20392
rect 11609 20383 11667 20389
rect 11609 20380 11621 20383
rect 11572 20352 11621 20380
rect 11572 20340 11578 20352
rect 11609 20349 11621 20352
rect 11655 20349 11667 20383
rect 11609 20343 11667 20349
rect 3007 20284 4568 20312
rect 3007 20281 3019 20284
rect 2961 20275 3019 20281
rect 5166 20272 5172 20324
rect 5224 20312 5230 20324
rect 6457 20315 6515 20321
rect 6457 20312 6469 20315
rect 5224 20284 6469 20312
rect 5224 20272 5230 20284
rect 6457 20281 6469 20284
rect 6503 20281 6515 20315
rect 9033 20315 9091 20321
rect 9033 20312 9045 20315
rect 6457 20275 6515 20281
rect 8036 20284 9045 20312
rect 1578 20204 1584 20256
rect 1636 20244 1642 20256
rect 1762 20244 1768 20256
rect 1636 20216 1768 20244
rect 1636 20204 1642 20216
rect 1762 20204 1768 20216
rect 1820 20204 1826 20256
rect 2409 20247 2467 20253
rect 2409 20213 2421 20247
rect 2455 20244 2467 20247
rect 3418 20244 3424 20256
rect 2455 20216 3424 20244
rect 2455 20213 2467 20216
rect 2409 20207 2467 20213
rect 3418 20204 3424 20216
rect 3476 20204 3482 20256
rect 5442 20204 5448 20256
rect 5500 20244 5506 20256
rect 5813 20247 5871 20253
rect 5813 20244 5825 20247
rect 5500 20216 5825 20244
rect 5500 20204 5506 20216
rect 5813 20213 5825 20216
rect 5859 20213 5871 20247
rect 5813 20207 5871 20213
rect 5994 20204 6000 20256
rect 6052 20244 6058 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 6052 20216 7113 20244
rect 6052 20204 6058 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7101 20207 7159 20213
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 8036 20244 8064 20284
rect 9033 20281 9045 20284
rect 9079 20281 9091 20315
rect 9033 20275 9091 20281
rect 10720 20315 10778 20321
rect 10720 20281 10732 20315
rect 10766 20312 10778 20315
rect 11425 20315 11483 20321
rect 11425 20312 11437 20315
rect 10766 20284 11437 20312
rect 10766 20281 10778 20284
rect 10720 20275 10778 20281
rect 11425 20281 11437 20284
rect 11471 20281 11483 20315
rect 11425 20275 11483 20281
rect 11624 20256 11652 20343
rect 11698 20340 11704 20392
rect 11756 20380 11762 20392
rect 11992 20389 12020 20420
rect 12434 20408 12440 20420
rect 12492 20408 12498 20460
rect 13354 20408 13360 20460
rect 13412 20408 13418 20460
rect 11793 20383 11851 20389
rect 11793 20380 11805 20383
rect 11756 20352 11805 20380
rect 11756 20340 11762 20352
rect 11793 20349 11805 20352
rect 11839 20349 11851 20383
rect 11793 20343 11851 20349
rect 11973 20383 12031 20389
rect 11973 20349 11985 20383
rect 12019 20349 12031 20383
rect 11973 20343 12031 20349
rect 12066 20340 12072 20392
rect 12124 20380 12130 20392
rect 12161 20383 12219 20389
rect 12161 20380 12173 20383
rect 12124 20352 12173 20380
rect 12124 20340 12130 20352
rect 12161 20349 12173 20352
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20380 12863 20383
rect 12986 20380 12992 20392
rect 12851 20352 12992 20380
rect 12851 20349 12863 20352
rect 12805 20343 12863 20349
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 14093 20383 14151 20389
rect 14093 20349 14105 20383
rect 14139 20380 14151 20383
rect 15470 20380 15476 20392
rect 14139 20352 15476 20380
rect 14139 20349 14151 20352
rect 14093 20343 14151 20349
rect 14476 20324 14504 20352
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 15930 20380 15936 20392
rect 15891 20352 15936 20380
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 16132 20389 16160 20488
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20448 16267 20451
rect 16408 20448 16436 20556
rect 16669 20553 16681 20587
rect 16715 20584 16727 20587
rect 16850 20584 16856 20596
rect 16715 20556 16856 20584
rect 16715 20553 16727 20556
rect 16669 20547 16727 20553
rect 16850 20544 16856 20556
rect 16908 20544 16914 20596
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 21450 20584 21456 20596
rect 20312 20556 21456 20584
rect 20312 20544 20318 20556
rect 21450 20544 21456 20556
rect 21508 20584 21514 20596
rect 22462 20584 22468 20596
rect 21508 20556 22324 20584
rect 22423 20556 22468 20584
rect 21508 20544 21514 20556
rect 16482 20476 16488 20528
rect 16540 20516 16546 20528
rect 17218 20516 17224 20528
rect 16540 20488 17224 20516
rect 16540 20476 16546 20488
rect 17218 20476 17224 20488
rect 17276 20476 17282 20528
rect 17678 20476 17684 20528
rect 17736 20516 17742 20528
rect 18506 20516 18512 20528
rect 17736 20488 18512 20516
rect 17736 20476 17742 20488
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 18874 20476 18880 20528
rect 18932 20516 18938 20528
rect 21358 20516 21364 20528
rect 18932 20488 21364 20516
rect 18932 20476 18938 20488
rect 21358 20476 21364 20488
rect 21416 20476 21422 20528
rect 22296 20516 22324 20556
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 23106 20584 23112 20596
rect 23067 20556 23112 20584
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 25498 20584 25504 20596
rect 23216 20556 24808 20584
rect 25459 20556 25504 20584
rect 23216 20516 23244 20556
rect 24578 20516 24584 20528
rect 22020 20488 23244 20516
rect 23308 20488 24584 20516
rect 17954 20448 17960 20460
rect 16255 20420 16436 20448
rect 17236 20420 17960 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 17236 20392 17264 20420
rect 17954 20408 17960 20420
rect 18012 20448 18018 20460
rect 19521 20451 19579 20457
rect 19521 20448 19533 20451
rect 18012 20420 19533 20448
rect 18012 20408 18018 20420
rect 19521 20417 19533 20420
rect 19567 20448 19579 20451
rect 19702 20448 19708 20460
rect 19567 20420 19708 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19702 20408 19708 20420
rect 19760 20448 19766 20460
rect 22020 20457 22048 20488
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 19760 20420 20821 20448
rect 19760 20408 19766 20420
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22152 20420 22197 20448
rect 22152 20408 22158 20420
rect 16117 20383 16175 20389
rect 16117 20349 16129 20383
rect 16163 20349 16175 20383
rect 16117 20343 16175 20349
rect 16301 20383 16359 20389
rect 16301 20349 16313 20383
rect 16347 20349 16359 20383
rect 16301 20343 16359 20349
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20380 16543 20383
rect 16574 20380 16580 20392
rect 16531 20352 16580 20380
rect 16531 20349 16543 20352
rect 16485 20343 16543 20349
rect 14366 20321 14372 20324
rect 14360 20312 14372 20321
rect 14327 20284 14372 20312
rect 14360 20275 14372 20284
rect 14366 20272 14372 20275
rect 14424 20272 14430 20324
rect 14458 20272 14464 20324
rect 14516 20272 14522 20324
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 15378 20312 15384 20324
rect 14884 20284 15384 20312
rect 14884 20272 14890 20284
rect 15378 20272 15384 20284
rect 15436 20272 15442 20324
rect 15838 20272 15844 20324
rect 15896 20312 15902 20324
rect 16316 20312 16344 20343
rect 16574 20340 16580 20352
rect 16632 20340 16638 20392
rect 17218 20340 17224 20392
rect 17276 20340 17282 20392
rect 18233 20383 18291 20389
rect 18233 20349 18245 20383
rect 18279 20349 18291 20383
rect 18506 20380 18512 20392
rect 18467 20352 18512 20380
rect 18233 20343 18291 20349
rect 15896 20284 16344 20312
rect 15896 20272 15902 20284
rect 17586 20272 17592 20324
rect 17644 20312 17650 20324
rect 18248 20312 18276 20343
rect 18506 20340 18512 20352
rect 18564 20340 18570 20392
rect 19245 20383 19303 20389
rect 19245 20380 19257 20383
rect 19168 20352 19257 20380
rect 18874 20312 18880 20324
rect 17644 20284 18880 20312
rect 17644 20272 17650 20284
rect 18874 20272 18880 20284
rect 18932 20272 18938 20324
rect 7984 20216 8064 20244
rect 8205 20247 8263 20253
rect 7984 20204 7990 20216
rect 8205 20213 8217 20247
rect 8251 20244 8263 20247
rect 8846 20244 8852 20256
rect 8251 20216 8852 20244
rect 8251 20213 8263 20216
rect 8205 20207 8263 20213
rect 8846 20204 8852 20216
rect 8904 20204 8910 20256
rect 9585 20247 9643 20253
rect 9585 20213 9597 20247
rect 9631 20244 9643 20247
rect 10410 20244 10416 20256
rect 9631 20216 10416 20244
rect 9631 20213 9643 20216
rect 9585 20207 9643 20213
rect 10410 20204 10416 20216
rect 10468 20244 10474 20256
rect 11606 20244 11612 20256
rect 10468 20216 11612 20244
rect 10468 20204 10474 20216
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 12710 20204 12716 20256
rect 12768 20244 12774 20256
rect 13173 20247 13231 20253
rect 13173 20244 13185 20247
rect 12768 20216 13185 20244
rect 12768 20204 12774 20216
rect 13173 20213 13185 20216
rect 13219 20244 13231 20247
rect 13262 20244 13268 20256
rect 13219 20216 13268 20244
rect 13219 20213 13231 20216
rect 13173 20207 13231 20213
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 15102 20204 15108 20256
rect 15160 20244 15166 20256
rect 15473 20247 15531 20253
rect 15473 20244 15485 20247
rect 15160 20216 15485 20244
rect 15160 20204 15166 20216
rect 15473 20213 15485 20216
rect 15519 20213 15531 20247
rect 15473 20207 15531 20213
rect 16666 20204 16672 20256
rect 16724 20244 16730 20256
rect 17129 20247 17187 20253
rect 17129 20244 17141 20247
rect 16724 20216 17141 20244
rect 16724 20204 16730 20216
rect 17129 20213 17141 20216
rect 17175 20244 17187 20247
rect 19168 20244 19196 20352
rect 19245 20349 19257 20352
rect 19291 20349 19303 20383
rect 19245 20343 19303 20349
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 20533 20383 20591 20389
rect 20533 20380 20545 20383
rect 20220 20352 20545 20380
rect 20220 20340 20226 20352
rect 20533 20349 20545 20352
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20378 20775 20383
rect 20763 20350 20852 20378
rect 20763 20349 20775 20350
rect 20717 20343 20775 20349
rect 20824 20312 20852 20350
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 20956 20352 21001 20380
rect 20956 20340 20962 20352
rect 21082 20340 21088 20392
rect 21140 20380 21146 20392
rect 21729 20383 21787 20389
rect 21729 20380 21741 20383
rect 21140 20352 21741 20380
rect 21140 20340 21146 20352
rect 21729 20349 21741 20352
rect 21775 20349 21787 20383
rect 21910 20380 21916 20392
rect 21871 20352 21916 20380
rect 21729 20343 21787 20349
rect 21910 20340 21916 20352
rect 21968 20340 21974 20392
rect 23308 20389 23336 20488
rect 24578 20476 24584 20488
rect 24636 20476 24642 20528
rect 24780 20516 24808 20556
rect 25498 20544 25504 20556
rect 25556 20544 25562 20596
rect 28718 20584 28724 20596
rect 25608 20556 28304 20584
rect 28679 20556 28724 20584
rect 25608 20516 25636 20556
rect 24780 20488 25636 20516
rect 28276 20516 28304 20556
rect 28718 20544 28724 20556
rect 28776 20544 28782 20596
rect 30929 20587 30987 20593
rect 30929 20553 30941 20587
rect 30975 20584 30987 20587
rect 31662 20584 31668 20596
rect 30975 20556 31668 20584
rect 30975 20553 30987 20556
rect 30929 20547 30987 20553
rect 31662 20544 31668 20556
rect 31720 20544 31726 20596
rect 30190 20516 30196 20528
rect 28276 20488 30196 20516
rect 30190 20476 30196 20488
rect 30248 20476 30254 20528
rect 23382 20408 23388 20460
rect 23440 20448 23446 20460
rect 23560 20451 23618 20457
rect 23560 20448 23572 20451
rect 23440 20420 23572 20448
rect 23440 20408 23446 20420
rect 23560 20417 23572 20420
rect 23606 20417 23618 20451
rect 30466 20448 30472 20460
rect 30427 20420 30472 20448
rect 23560 20411 23618 20417
rect 30466 20408 30472 20420
rect 30524 20408 30530 20460
rect 30650 20448 30656 20460
rect 30611 20420 30656 20448
rect 30650 20408 30656 20420
rect 30708 20408 30714 20460
rect 22281 20383 22339 20389
rect 22281 20349 22293 20383
rect 22327 20349 22339 20383
rect 22281 20343 22339 20349
rect 23293 20383 23351 20389
rect 23293 20349 23305 20383
rect 23339 20349 23351 20383
rect 23293 20343 23351 20349
rect 23477 20383 23535 20389
rect 23477 20349 23489 20383
rect 23523 20349 23535 20383
rect 23477 20343 23535 20349
rect 21174 20312 21180 20324
rect 20824 20284 21180 20312
rect 21174 20272 21180 20284
rect 21232 20312 21238 20324
rect 22002 20312 22008 20324
rect 21232 20284 22008 20312
rect 21232 20272 21238 20284
rect 22002 20272 22008 20284
rect 22060 20312 22066 20324
rect 22296 20312 22324 20343
rect 22060 20284 22324 20312
rect 23492 20312 23520 20343
rect 23658 20340 23664 20392
rect 23716 20380 23722 20392
rect 23716 20352 23761 20380
rect 23716 20340 23722 20352
rect 23842 20340 23848 20392
rect 23900 20380 23906 20392
rect 24762 20380 24768 20392
rect 23900 20352 23945 20380
rect 24596 20352 24768 20380
rect 23900 20340 23906 20352
rect 24596 20312 24624 20352
rect 24762 20340 24768 20352
rect 24820 20340 24826 20392
rect 26234 20340 26240 20392
rect 26292 20380 26298 20392
rect 26881 20383 26939 20389
rect 26881 20380 26893 20383
rect 26292 20352 26893 20380
rect 26292 20340 26298 20352
rect 26881 20349 26893 20352
rect 26927 20380 26939 20383
rect 27341 20383 27399 20389
rect 27341 20380 27353 20383
rect 26927 20352 27353 20380
rect 26927 20349 26939 20352
rect 26881 20343 26939 20349
rect 27341 20349 27353 20352
rect 27387 20349 27399 20383
rect 27341 20343 27399 20349
rect 27608 20383 27666 20389
rect 27608 20349 27620 20383
rect 27654 20380 27666 20383
rect 27982 20380 27988 20392
rect 27654 20352 27988 20380
rect 27654 20349 27666 20352
rect 27608 20343 27666 20349
rect 27982 20340 27988 20352
rect 28040 20340 28046 20392
rect 28718 20340 28724 20392
rect 28776 20380 28782 20392
rect 29733 20383 29791 20389
rect 29733 20380 29745 20383
rect 28776 20352 29745 20380
rect 28776 20340 28782 20352
rect 29733 20349 29745 20352
rect 29779 20349 29791 20383
rect 29733 20343 29791 20349
rect 29825 20383 29883 20389
rect 29825 20349 29837 20383
rect 29871 20380 29883 20383
rect 30282 20380 30288 20392
rect 29871 20352 30288 20380
rect 29871 20349 29883 20352
rect 29825 20343 29883 20349
rect 30282 20340 30288 20352
rect 30340 20380 30346 20392
rect 30561 20383 30619 20389
rect 30561 20380 30573 20383
rect 30340 20352 30573 20380
rect 30340 20340 30346 20352
rect 30561 20349 30573 20352
rect 30607 20349 30619 20383
rect 30561 20343 30619 20349
rect 30745 20383 30803 20389
rect 30745 20349 30757 20383
rect 30791 20380 30803 20383
rect 30926 20380 30932 20392
rect 30791 20352 30932 20380
rect 30791 20349 30803 20352
rect 30745 20343 30803 20349
rect 23492 20284 24624 20312
rect 24673 20315 24731 20321
rect 22060 20272 22066 20284
rect 24673 20281 24685 20315
rect 24719 20312 24731 20315
rect 25130 20312 25136 20324
rect 24719 20284 25136 20312
rect 24719 20281 24731 20284
rect 24673 20275 24731 20281
rect 25130 20272 25136 20284
rect 25188 20272 25194 20324
rect 26602 20272 26608 20324
rect 26660 20321 26666 20324
rect 26660 20312 26672 20321
rect 26660 20284 26705 20312
rect 26660 20275 26672 20284
rect 26660 20272 26666 20275
rect 30466 20272 30472 20324
rect 30524 20312 30530 20324
rect 30760 20312 30788 20343
rect 30926 20340 30932 20352
rect 30984 20340 30990 20392
rect 30524 20284 30788 20312
rect 30524 20272 30530 20284
rect 20806 20244 20812 20256
rect 17175 20216 20812 20244
rect 17175 20213 17187 20216
rect 17129 20207 17187 20213
rect 20806 20204 20812 20216
rect 20864 20204 20870 20256
rect 21266 20244 21272 20256
rect 21227 20216 21272 20244
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 21358 20204 21364 20256
rect 21416 20244 21422 20256
rect 24946 20244 24952 20256
rect 21416 20216 24952 20244
rect 21416 20204 21422 20216
rect 24946 20204 24952 20216
rect 25004 20204 25010 20256
rect 1104 20154 32016 20176
rect 1104 20102 11253 20154
rect 11305 20102 11317 20154
rect 11369 20102 11381 20154
rect 11433 20102 11445 20154
rect 11497 20102 11509 20154
rect 11561 20102 21557 20154
rect 21609 20102 21621 20154
rect 21673 20102 21685 20154
rect 21737 20102 21749 20154
rect 21801 20102 21813 20154
rect 21865 20102 32016 20154
rect 1104 20080 32016 20102
rect 1302 20000 1308 20052
rect 1360 20040 1366 20052
rect 1486 20040 1492 20052
rect 1360 20012 1492 20040
rect 1360 20000 1366 20012
rect 1486 20000 1492 20012
rect 1544 20000 1550 20052
rect 2958 20040 2964 20052
rect 2919 20012 2964 20040
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 4246 20040 4252 20052
rect 4207 20012 4252 20040
rect 4246 20000 4252 20012
rect 4304 20000 4310 20052
rect 5350 20000 5356 20052
rect 5408 20040 5414 20052
rect 8202 20040 8208 20052
rect 5408 20012 5488 20040
rect 8163 20012 8208 20040
rect 5408 20000 5414 20012
rect 2406 19972 2412 19984
rect 2332 19944 2412 19972
rect 1486 19904 1492 19916
rect 1447 19876 1492 19904
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 1670 19864 1676 19916
rect 1728 19904 1734 19916
rect 2332 19913 2360 19944
rect 2406 19932 2412 19944
rect 2464 19932 2470 19984
rect 4614 19932 4620 19984
rect 4672 19972 4678 19984
rect 4890 19972 4896 19984
rect 4672 19944 4896 19972
rect 4672 19932 4678 19944
rect 4890 19932 4896 19944
rect 4948 19972 4954 19984
rect 5460 19972 5488 20012
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 10502 20000 10508 20052
rect 10560 20040 10566 20052
rect 10781 20043 10839 20049
rect 10781 20040 10793 20043
rect 10560 20012 10793 20040
rect 10560 20000 10566 20012
rect 10781 20009 10793 20012
rect 10827 20040 10839 20043
rect 10962 20040 10968 20052
rect 10827 20012 10968 20040
rect 10827 20009 10839 20012
rect 10781 20003 10839 20009
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 13446 20040 13452 20052
rect 12676 20012 13308 20040
rect 13407 20012 13452 20040
rect 12676 20000 12682 20012
rect 4948 19944 5396 19972
rect 4948 19932 4954 19944
rect 2317 19907 2375 19913
rect 2317 19904 2329 19907
rect 1728 19876 2329 19904
rect 1728 19864 1734 19876
rect 2317 19873 2329 19876
rect 2363 19873 2375 19907
rect 2498 19904 2504 19916
rect 2459 19876 2504 19904
rect 2317 19867 2375 19873
rect 2498 19864 2504 19876
rect 2556 19864 2562 19916
rect 2593 19907 2651 19913
rect 2593 19873 2605 19907
rect 2639 19873 2651 19907
rect 2593 19867 2651 19873
rect 2685 19907 2743 19913
rect 2685 19873 2697 19907
rect 2731 19904 2743 19907
rect 3418 19904 3424 19916
rect 2731 19876 2912 19904
rect 3379 19876 3424 19904
rect 2731 19873 2743 19876
rect 2685 19867 2743 19873
rect 2608 19768 2636 19867
rect 2884 19780 2912 19876
rect 3418 19864 3424 19876
rect 3476 19864 3482 19916
rect 3602 19904 3608 19916
rect 3563 19876 3608 19904
rect 3602 19864 3608 19876
rect 3660 19864 3666 19916
rect 4154 19904 4160 19916
rect 4115 19876 4160 19904
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 5368 19913 5396 19944
rect 5460 19944 6408 19972
rect 5460 19913 5488 19944
rect 6380 19913 6408 19944
rect 7650 19932 7656 19984
rect 7708 19972 7714 19984
rect 7708 19944 7880 19972
rect 7708 19932 7714 19944
rect 5261 19907 5319 19913
rect 5261 19904 5273 19907
rect 5092 19876 5273 19904
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 2608 19740 2774 19768
rect 1762 19700 1768 19712
rect 1723 19672 1768 19700
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 2746 19700 2774 19740
rect 2866 19728 2872 19780
rect 2924 19768 2930 19780
rect 3804 19768 3832 19799
rect 2924 19740 3832 19768
rect 5092 19768 5120 19876
rect 5261 19873 5273 19876
rect 5307 19873 5319 19907
rect 5261 19867 5319 19873
rect 5350 19907 5408 19913
rect 5350 19873 5362 19907
rect 5396 19873 5408 19907
rect 5350 19867 5408 19873
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19873 5687 19907
rect 5629 19867 5687 19873
rect 6365 19907 6423 19913
rect 6365 19873 6377 19907
rect 6411 19873 6423 19907
rect 6546 19904 6552 19916
rect 6507 19876 6552 19904
rect 6365 19867 6423 19873
rect 5166 19796 5172 19848
rect 5224 19836 5230 19848
rect 5644 19836 5672 19867
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 7561 19907 7619 19913
rect 7561 19873 7573 19907
rect 7607 19873 7619 19907
rect 7742 19904 7748 19916
rect 7703 19876 7748 19904
rect 7561 19867 7619 19873
rect 5224 19808 5672 19836
rect 5224 19796 5230 19808
rect 5258 19768 5264 19780
rect 5092 19740 5264 19768
rect 2924 19728 2930 19740
rect 5258 19728 5264 19740
rect 5316 19768 5322 19780
rect 5994 19768 6000 19780
rect 5316 19740 6000 19768
rect 5316 19728 5322 19740
rect 5994 19728 6000 19740
rect 6052 19728 6058 19780
rect 7576 19768 7604 19867
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 7852 19913 7880 19944
rect 8018 19932 8024 19984
rect 8076 19972 8082 19984
rect 12894 19972 12900 19984
rect 8076 19944 8708 19972
rect 8076 19932 8082 19944
rect 7837 19907 7895 19913
rect 7837 19873 7849 19907
rect 7883 19873 7895 19907
rect 7837 19867 7895 19873
rect 7926 19864 7932 19916
rect 7984 19904 7990 19916
rect 8680 19913 8708 19944
rect 12728 19944 12900 19972
rect 8665 19907 8723 19913
rect 7984 19876 8029 19904
rect 7984 19864 7990 19876
rect 8665 19873 8677 19907
rect 8711 19873 8723 19907
rect 8665 19867 8723 19873
rect 9122 19864 9128 19916
rect 9180 19904 9186 19916
rect 9401 19907 9459 19913
rect 9401 19904 9413 19907
rect 9180 19876 9413 19904
rect 9180 19864 9186 19876
rect 9401 19873 9413 19876
rect 9447 19873 9459 19907
rect 10410 19904 10416 19916
rect 10371 19876 10416 19904
rect 9401 19867 9459 19873
rect 10410 19864 10416 19876
rect 10468 19864 10474 19916
rect 11974 19904 11980 19916
rect 11935 19876 11980 19904
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12728 19913 12756 19944
rect 12894 19932 12900 19944
rect 12952 19932 12958 19984
rect 13280 19972 13308 20012
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 14093 20043 14151 20049
rect 14093 20009 14105 20043
rect 14139 20040 14151 20043
rect 14182 20040 14188 20052
rect 14139 20012 14188 20040
rect 14139 20009 14151 20012
rect 14093 20003 14151 20009
rect 14182 20000 14188 20012
rect 14240 20040 14246 20052
rect 14826 20040 14832 20052
rect 14240 20012 14832 20040
rect 14240 20000 14246 20012
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 18966 20000 18972 20052
rect 19024 20040 19030 20052
rect 19024 20012 19472 20040
rect 19024 20000 19030 20012
rect 13280 19944 15700 19972
rect 12161 19907 12219 19913
rect 12161 19873 12173 19907
rect 12207 19873 12219 19907
rect 12161 19867 12219 19873
rect 12713 19907 12771 19913
rect 12713 19873 12725 19907
rect 12759 19873 12771 19907
rect 13354 19904 13360 19916
rect 13315 19876 13360 19904
rect 12713 19867 12771 19873
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 8168 19808 8953 19836
rect 8168 19796 8174 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 8478 19768 8484 19780
rect 7576 19740 8484 19768
rect 8478 19728 8484 19740
rect 8536 19728 8542 19780
rect 10965 19771 11023 19777
rect 10965 19737 10977 19771
rect 11011 19768 11023 19771
rect 12176 19768 12204 19867
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 14274 19864 14280 19916
rect 14332 19904 14338 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14332 19876 14749 19904
rect 14332 19864 14338 19876
rect 14737 19873 14749 19876
rect 14783 19904 14795 19907
rect 15102 19904 15108 19916
rect 14783 19876 15108 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 15378 19904 15384 19916
rect 15339 19876 15384 19904
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 15672 19913 15700 19944
rect 16114 19932 16120 19984
rect 16172 19972 16178 19984
rect 17678 19972 17684 19984
rect 16172 19944 17684 19972
rect 16172 19932 16178 19944
rect 17678 19932 17684 19944
rect 17736 19932 17742 19984
rect 17896 19975 17954 19981
rect 17896 19941 17908 19975
rect 17942 19972 17954 19975
rect 19337 19975 19395 19981
rect 19337 19972 19349 19975
rect 17942 19944 19349 19972
rect 17942 19941 17954 19944
rect 17896 19935 17954 19941
rect 19337 19941 19349 19944
rect 19383 19941 19395 19975
rect 19444 19972 19472 20012
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 21269 20043 21327 20049
rect 21269 20040 21281 20043
rect 21232 20012 21281 20040
rect 21232 20000 21238 20012
rect 21269 20009 21281 20012
rect 21315 20009 21327 20043
rect 21269 20003 21327 20009
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 24581 20043 24639 20049
rect 24581 20040 24593 20043
rect 23716 20012 24593 20040
rect 23716 20000 23722 20012
rect 24581 20009 24593 20012
rect 24627 20040 24639 20043
rect 26142 20040 26148 20052
rect 24627 20012 26148 20040
rect 24627 20009 24639 20012
rect 24581 20003 24639 20009
rect 26142 20000 26148 20012
rect 26200 20000 26206 20052
rect 31110 20000 31116 20052
rect 31168 20040 31174 20052
rect 31205 20043 31263 20049
rect 31205 20040 31217 20043
rect 31168 20012 31217 20040
rect 31168 20000 31174 20012
rect 31205 20009 31217 20012
rect 31251 20009 31263 20043
rect 31205 20003 31263 20009
rect 22094 19972 22100 19984
rect 19444 19944 22100 19972
rect 19337 19935 19395 19941
rect 22094 19932 22100 19944
rect 22152 19932 22158 19984
rect 25716 19975 25774 19981
rect 25716 19941 25728 19975
rect 25762 19972 25774 19975
rect 26326 19972 26332 19984
rect 25762 19944 26332 19972
rect 25762 19941 25774 19944
rect 25716 19935 25774 19941
rect 26326 19932 26332 19944
rect 26384 19932 26390 19984
rect 31018 19972 31024 19984
rect 29012 19944 31024 19972
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19873 15623 19907
rect 15565 19867 15623 19873
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19904 15715 19907
rect 15838 19904 15844 19916
rect 15703 19876 15844 19904
rect 15703 19873 15715 19876
rect 15657 19867 15715 19873
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 13170 19836 13176 19848
rect 12943 19808 13176 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 15580 19836 15608 19867
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 15933 19907 15991 19913
rect 15933 19873 15945 19907
rect 15979 19904 15991 19907
rect 16206 19904 16212 19916
rect 15979 19876 16212 19904
rect 15979 19873 15991 19876
rect 15933 19867 15991 19873
rect 14875 19828 15148 19836
rect 15212 19828 15608 19836
rect 14875 19808 15608 19828
rect 15749 19839 15807 19845
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 15120 19800 15240 19808
rect 15749 19805 15761 19839
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 11011 19740 12204 19768
rect 11011 19737 11023 19740
rect 10965 19731 11023 19737
rect 15286 19728 15292 19780
rect 15344 19768 15350 19780
rect 15764 19768 15792 19799
rect 15344 19740 15792 19768
rect 15344 19728 15350 19740
rect 15838 19728 15844 19780
rect 15896 19768 15902 19780
rect 15948 19768 15976 19867
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 17126 19904 17132 19916
rect 16632 19876 17132 19904
rect 16632 19864 16638 19876
rect 17126 19864 17132 19876
rect 17184 19904 17190 19916
rect 18598 19904 18604 19916
rect 17184 19876 18276 19904
rect 18559 19876 18604 19904
rect 17184 19864 17190 19876
rect 16666 19836 16672 19848
rect 15896 19740 15976 19768
rect 16040 19808 16672 19836
rect 15896 19728 15902 19740
rect 3326 19700 3332 19712
rect 2746 19672 3332 19700
rect 3326 19660 3332 19672
rect 3384 19660 3390 19712
rect 4982 19700 4988 19712
rect 4943 19672 4988 19700
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 6549 19703 6607 19709
rect 6549 19669 6561 19703
rect 6595 19700 6607 19703
rect 6822 19700 6828 19712
rect 6595 19672 6828 19700
rect 6595 19669 6607 19672
rect 6549 19663 6607 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7006 19700 7012 19712
rect 6967 19672 7012 19700
rect 7006 19660 7012 19672
rect 7064 19660 7070 19712
rect 8570 19660 8576 19712
rect 8628 19700 8634 19712
rect 8754 19700 8760 19712
rect 8628 19672 8760 19700
rect 8628 19660 8634 19672
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 8849 19703 8907 19709
rect 8849 19669 8861 19703
rect 8895 19700 8907 19703
rect 9398 19700 9404 19712
rect 8895 19672 9404 19700
rect 8895 19669 8907 19672
rect 8849 19663 8907 19669
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 9493 19703 9551 19709
rect 9493 19669 9505 19703
rect 9539 19700 9551 19703
rect 9766 19700 9772 19712
rect 9539 19672 9772 19700
rect 9539 19669 9551 19672
rect 9493 19663 9551 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 10781 19703 10839 19709
rect 10781 19669 10793 19703
rect 10827 19700 10839 19703
rect 11146 19700 11152 19712
rect 10827 19672 11152 19700
rect 10827 19669 10839 19672
rect 10781 19663 10839 19669
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 16040 19700 16068 19808
rect 16666 19796 16672 19808
rect 16724 19796 16730 19848
rect 18138 19836 18144 19848
rect 18099 19808 18144 19836
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18248 19836 18276 19876
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19873 18843 19907
rect 18966 19904 18972 19916
rect 18927 19876 18972 19904
rect 18785 19867 18843 19873
rect 18800 19836 18828 19867
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 19153 19907 19211 19913
rect 19153 19904 19165 19907
rect 19076 19876 19165 19904
rect 18248 19808 18828 19836
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 16117 19771 16175 19777
rect 16117 19737 16129 19771
rect 16163 19768 16175 19771
rect 16850 19768 16856 19780
rect 16163 19740 16856 19768
rect 16163 19737 16175 19740
rect 16117 19731 16175 19737
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 18690 19728 18696 19780
rect 18748 19768 18754 19780
rect 18892 19768 18920 19799
rect 18748 19740 18920 19768
rect 18748 19728 18754 19740
rect 13872 19672 16068 19700
rect 16761 19703 16819 19709
rect 13872 19660 13878 19672
rect 16761 19669 16773 19703
rect 16807 19700 16819 19703
rect 17402 19700 17408 19712
rect 16807 19672 17408 19700
rect 16807 19669 16819 19672
rect 16761 19663 16819 19669
rect 17402 19660 17408 19672
rect 17460 19700 17466 19712
rect 19076 19700 19104 19876
rect 19153 19873 19165 19876
rect 19199 19873 19211 19907
rect 19153 19867 19211 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19889 19907 19947 19913
rect 19889 19904 19901 19907
rect 19668 19876 19901 19904
rect 19668 19864 19674 19876
rect 19889 19873 19901 19876
rect 19935 19873 19947 19907
rect 19889 19867 19947 19873
rect 20156 19907 20214 19913
rect 20156 19873 20168 19907
rect 20202 19904 20214 19907
rect 20898 19904 20904 19916
rect 20202 19876 20904 19904
rect 20202 19873 20214 19876
rect 20156 19867 20214 19873
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19904 22247 19907
rect 22278 19904 22284 19916
rect 22235 19876 22284 19904
rect 22235 19873 22247 19876
rect 22189 19867 22247 19873
rect 22278 19864 22284 19876
rect 22336 19864 22342 19916
rect 22462 19913 22468 19916
rect 22456 19867 22468 19913
rect 22520 19904 22526 19916
rect 27522 19904 27528 19916
rect 22520 19876 22556 19904
rect 27483 19876 27528 19904
rect 22462 19864 22468 19867
rect 22520 19864 22526 19876
rect 27522 19864 27528 19876
rect 27580 19864 27586 19916
rect 28074 19864 28080 19916
rect 28132 19904 28138 19916
rect 29012 19913 29040 19944
rect 31018 19932 31024 19944
rect 31076 19932 31082 19984
rect 31386 19972 31392 19984
rect 31128 19944 31392 19972
rect 28445 19907 28503 19913
rect 28445 19904 28457 19907
rect 28132 19876 28457 19904
rect 28132 19864 28138 19876
rect 28445 19873 28457 19876
rect 28491 19873 28503 19907
rect 28445 19867 28503 19873
rect 28997 19907 29055 19913
rect 28997 19873 29009 19907
rect 29043 19873 29055 19907
rect 28997 19867 29055 19873
rect 29825 19907 29883 19913
rect 29825 19873 29837 19907
rect 29871 19904 29883 19907
rect 30653 19907 30711 19913
rect 29871 19876 30512 19904
rect 29871 19873 29883 19876
rect 29825 19867 29883 19873
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19836 26019 19839
rect 26234 19836 26240 19848
rect 26007 19808 26240 19836
rect 26007 19805 26019 19808
rect 25961 19799 26019 19805
rect 26234 19796 26240 19808
rect 26292 19796 26298 19848
rect 27801 19839 27859 19845
rect 27801 19805 27813 19839
rect 27847 19836 27859 19839
rect 28902 19836 28908 19848
rect 27847 19808 28908 19836
rect 27847 19805 27859 19808
rect 27801 19799 27859 19805
rect 17460 19672 19104 19700
rect 17460 19660 17466 19672
rect 19150 19660 19156 19712
rect 19208 19700 19214 19712
rect 21358 19700 21364 19712
rect 19208 19672 21364 19700
rect 19208 19660 19214 19672
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 23290 19660 23296 19712
rect 23348 19700 23354 19712
rect 23569 19703 23627 19709
rect 23569 19700 23581 19703
rect 23348 19672 23581 19700
rect 23348 19660 23354 19672
rect 23569 19669 23581 19672
rect 23615 19669 23627 19703
rect 23569 19663 23627 19669
rect 24121 19703 24179 19709
rect 24121 19669 24133 19703
rect 24167 19700 24179 19703
rect 24394 19700 24400 19712
rect 24167 19672 24400 19700
rect 24167 19669 24179 19672
rect 24121 19663 24179 19669
rect 24394 19660 24400 19672
rect 24452 19700 24458 19712
rect 27816 19700 27844 19799
rect 28902 19796 28908 19808
rect 28960 19796 28966 19848
rect 30484 19777 30512 19876
rect 30653 19873 30665 19907
rect 30699 19904 30711 19907
rect 30742 19904 30748 19916
rect 30699 19876 30748 19904
rect 30699 19873 30711 19876
rect 30653 19867 30711 19873
rect 30742 19864 30748 19876
rect 30800 19904 30806 19916
rect 31128 19904 31156 19944
rect 31386 19932 31392 19944
rect 31444 19932 31450 19984
rect 31294 19904 31300 19916
rect 30800 19876 31156 19904
rect 31255 19876 31300 19904
rect 30800 19864 30806 19876
rect 31294 19864 31300 19876
rect 31352 19864 31358 19916
rect 30469 19771 30527 19777
rect 30469 19737 30481 19771
rect 30515 19737 30527 19771
rect 30469 19731 30527 19737
rect 31128 19740 31754 19768
rect 28350 19700 28356 19712
rect 24452 19672 27844 19700
rect 28311 19672 28356 19700
rect 24452 19660 24458 19672
rect 28350 19660 28356 19672
rect 28408 19660 28414 19712
rect 29181 19703 29239 19709
rect 29181 19669 29193 19703
rect 29227 19700 29239 19703
rect 29914 19700 29920 19712
rect 29227 19672 29920 19700
rect 29227 19669 29239 19672
rect 29181 19663 29239 19669
rect 29914 19660 29920 19672
rect 29972 19660 29978 19712
rect 30009 19703 30067 19709
rect 30009 19669 30021 19703
rect 30055 19700 30067 19703
rect 31128 19700 31156 19740
rect 30055 19672 31156 19700
rect 31726 19700 31754 19740
rect 31726 19672 32352 19700
rect 30055 19669 30067 19672
rect 30009 19663 30067 19669
rect 1104 19610 32016 19632
rect 1104 19558 6102 19610
rect 6154 19558 6166 19610
rect 6218 19558 6230 19610
rect 6282 19558 6294 19610
rect 6346 19558 6358 19610
rect 6410 19558 16405 19610
rect 16457 19558 16469 19610
rect 16521 19558 16533 19610
rect 16585 19558 16597 19610
rect 16649 19558 16661 19610
rect 16713 19558 26709 19610
rect 26761 19558 26773 19610
rect 26825 19558 26837 19610
rect 26889 19558 26901 19610
rect 26953 19558 26965 19610
rect 27017 19558 32016 19610
rect 32324 19564 32352 19672
rect 1104 19536 32016 19558
rect 32232 19536 32352 19564
rect 1762 19456 1768 19508
rect 1820 19496 1826 19508
rect 2682 19496 2688 19508
rect 1820 19468 2688 19496
rect 1820 19456 1826 19468
rect 2682 19456 2688 19468
rect 2740 19496 2746 19508
rect 2740 19456 2774 19496
rect 3602 19456 3608 19508
rect 3660 19496 3666 19508
rect 6917 19499 6975 19505
rect 6917 19496 6929 19499
rect 3660 19468 6929 19496
rect 3660 19456 3666 19468
rect 6917 19465 6929 19468
rect 6963 19496 6975 19499
rect 7006 19496 7012 19508
rect 6963 19468 7012 19496
rect 6963 19465 6975 19468
rect 6917 19459 6975 19465
rect 7006 19456 7012 19468
rect 7064 19496 7070 19508
rect 7282 19496 7288 19508
rect 7064 19468 7288 19496
rect 7064 19456 7070 19468
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 13354 19496 13360 19508
rect 12492 19468 13360 19496
rect 12492 19456 12498 19468
rect 0 19428 800 19442
rect 2746 19440 2774 19456
rect 1486 19428 1492 19440
rect 0 19400 1492 19428
rect 0 19386 800 19400
rect 1486 19388 1492 19400
rect 1544 19428 1550 19440
rect 2406 19428 2412 19440
rect 1544 19400 2412 19428
rect 1544 19388 1550 19400
rect 2406 19388 2412 19400
rect 2464 19388 2470 19440
rect 2746 19400 2780 19440
rect 2774 19388 2780 19400
rect 2832 19388 2838 19440
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 3476 19400 4108 19428
rect 3476 19388 3482 19400
rect 3878 19360 3884 19372
rect 2792 19332 3096 19360
rect 3839 19332 3884 19360
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 2038 19292 2044 19304
rect 1903 19264 2044 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2314 19252 2320 19304
rect 2372 19292 2378 19304
rect 2792 19301 2820 19332
rect 2489 19295 2547 19301
rect 2489 19294 2501 19295
rect 2424 19292 2501 19294
rect 2372 19266 2501 19292
rect 2372 19264 2452 19266
rect 2372 19252 2378 19264
rect 2489 19261 2501 19266
rect 2535 19261 2547 19295
rect 2489 19255 2547 19261
rect 2664 19292 2722 19298
rect 2664 19258 2676 19292
rect 2710 19258 2722 19292
rect 2664 19252 2722 19258
rect 2764 19295 2822 19301
rect 2764 19261 2776 19295
rect 2810 19261 2822 19295
rect 2764 19255 2822 19261
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 3068 19292 3096 19332
rect 3878 19320 3884 19332
rect 3936 19320 3942 19372
rect 4080 19369 4108 19400
rect 4614 19388 4620 19440
rect 4672 19428 4678 19440
rect 5166 19428 5172 19440
rect 4672 19400 5172 19428
rect 4672 19388 4678 19400
rect 5166 19388 5172 19400
rect 5224 19388 5230 19440
rect 5442 19388 5448 19440
rect 5500 19388 5506 19440
rect 6733 19431 6791 19437
rect 6733 19428 6745 19431
rect 6288 19400 6745 19428
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4246 19320 4252 19372
rect 4304 19360 4310 19372
rect 5460 19360 5488 19388
rect 6288 19369 6316 19400
rect 6733 19397 6745 19400
rect 6779 19397 6791 19431
rect 6733 19391 6791 19397
rect 9677 19431 9735 19437
rect 9677 19397 9689 19431
rect 9723 19428 9735 19431
rect 11698 19428 11704 19440
rect 9723 19400 9996 19428
rect 9723 19397 9735 19400
rect 9677 19391 9735 19397
rect 4304 19332 5488 19360
rect 6273 19363 6331 19369
rect 4304 19320 4310 19332
rect 6273 19329 6285 19363
rect 6319 19329 6331 19363
rect 8018 19360 8024 19372
rect 7979 19332 8024 19360
rect 6273 19323 6331 19329
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 8386 19360 8392 19372
rect 8347 19332 8392 19360
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 9456 19332 9505 19360
rect 9456 19320 9462 19332
rect 9493 19329 9505 19332
rect 9539 19329 9551 19363
rect 9766 19360 9772 19372
rect 9727 19332 9772 19360
rect 9493 19323 9551 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 3418 19292 3424 19304
rect 2924 19264 2969 19292
rect 3068 19264 3424 19292
rect 2924 19252 2930 19264
rect 3418 19252 3424 19264
rect 3476 19252 3482 19304
rect 4430 19252 4436 19304
rect 4488 19292 4494 19304
rect 5445 19295 5503 19301
rect 5445 19292 5457 19295
rect 4488 19264 5457 19292
rect 4488 19252 4494 19264
rect 5445 19261 5457 19264
rect 5491 19261 5503 19295
rect 5626 19292 5632 19304
rect 5587 19264 5632 19292
rect 5445 19255 5503 19261
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 5994 19292 6000 19304
rect 5955 19264 6000 19292
rect 5994 19252 6000 19264
rect 6052 19252 6058 19304
rect 6730 19252 6736 19304
rect 6788 19292 6794 19304
rect 7650 19292 7656 19304
rect 6788 19264 7144 19292
rect 7611 19264 7656 19292
rect 6788 19252 6794 19264
rect 2056 19224 2084 19252
rect 2679 19224 2707 19252
rect 3142 19224 3148 19236
rect 2056 19196 2707 19224
rect 3103 19196 3148 19224
rect 3142 19184 3148 19196
rect 3200 19184 3206 19236
rect 3436 19224 3464 19252
rect 3436 19196 6776 19224
rect 1949 19159 2007 19165
rect 1949 19125 1961 19159
rect 1995 19156 2007 19159
rect 2682 19156 2688 19168
rect 1995 19128 2688 19156
rect 1995 19125 2007 19128
rect 1949 19119 2007 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3050 19116 3056 19168
rect 3108 19156 3114 19168
rect 3786 19156 3792 19168
rect 3108 19128 3792 19156
rect 3108 19116 3114 19128
rect 3786 19116 3792 19128
rect 3844 19156 3850 19168
rect 4157 19159 4215 19165
rect 4157 19156 4169 19159
rect 3844 19128 4169 19156
rect 3844 19116 3850 19128
rect 4157 19125 4169 19128
rect 4203 19125 4215 19159
rect 4522 19156 4528 19168
rect 4483 19128 4528 19156
rect 4157 19119 4215 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 6546 19156 6552 19168
rect 6319 19128 6552 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 6748 19156 6776 19196
rect 6822 19184 6828 19236
rect 6880 19233 6886 19236
rect 7116 19233 7144 19264
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 7745 19295 7803 19301
rect 7745 19261 7757 19295
rect 7791 19261 7803 19295
rect 7745 19255 7803 19261
rect 6880 19227 6943 19233
rect 6880 19193 6897 19227
rect 6931 19193 6943 19227
rect 6880 19187 6943 19193
rect 7101 19227 7159 19233
rect 7101 19193 7113 19227
rect 7147 19193 7159 19227
rect 7101 19187 7159 19193
rect 6880 19184 6886 19187
rect 7760 19156 7788 19255
rect 8846 19252 8852 19304
rect 8904 19292 8910 19304
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 8904 19264 9229 19292
rect 8904 19252 8910 19264
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 8205 19227 8263 19233
rect 8205 19193 8217 19227
rect 8251 19224 8263 19227
rect 9876 19224 9904 19255
rect 8251 19196 9904 19224
rect 9968 19224 9996 19400
rect 11256 19400 11704 19428
rect 11256 19369 11284 19400
rect 11698 19388 11704 19400
rect 11756 19388 11762 19440
rect 12618 19428 12624 19440
rect 12452 19400 12624 19428
rect 12452 19369 12480 19400
rect 12618 19388 12624 19400
rect 12676 19388 12682 19440
rect 11241 19363 11299 19369
rect 11241 19329 11253 19363
rect 11287 19329 11299 19363
rect 11241 19323 11299 19329
rect 11333 19363 11391 19369
rect 11333 19329 11345 19363
rect 11379 19360 11391 19363
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 11379 19332 12449 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12584 19332 12629 19360
rect 12584 19320 12590 19332
rect 10502 19252 10508 19304
rect 10560 19292 10566 19304
rect 11057 19295 11115 19301
rect 11057 19292 11069 19295
rect 10560 19264 11069 19292
rect 10560 19252 10566 19264
rect 11057 19261 11069 19264
rect 11103 19261 11115 19295
rect 11057 19255 11115 19261
rect 11425 19295 11483 19301
rect 11425 19261 11437 19295
rect 11471 19292 11483 19295
rect 11514 19292 11520 19304
rect 11471 19264 11520 19292
rect 11471 19261 11483 19264
rect 11425 19255 11483 19261
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 11609 19295 11667 19301
rect 11609 19261 11621 19295
rect 11655 19292 11667 19295
rect 11655 19264 11928 19292
rect 11655 19261 11667 19264
rect 11609 19255 11667 19261
rect 11790 19224 11796 19236
rect 9968 19196 11796 19224
rect 8251 19193 8263 19196
rect 8205 19187 8263 19193
rect 11790 19184 11796 19196
rect 11848 19184 11854 19236
rect 11900 19224 11928 19264
rect 11974 19252 11980 19304
rect 12032 19292 12038 19304
rect 12728 19301 12756 19468
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 15378 19496 15384 19508
rect 15028 19468 15384 19496
rect 12894 19388 12900 19440
rect 12952 19428 12958 19440
rect 13449 19431 13507 19437
rect 13449 19428 13461 19431
rect 12952 19400 13461 19428
rect 12952 19388 12958 19400
rect 13449 19397 13461 19400
rect 13495 19428 13507 19431
rect 13538 19428 13544 19440
rect 13495 19400 13544 19428
rect 13495 19397 13507 19400
rect 13449 19391 13507 19397
rect 13538 19388 13544 19400
rect 13596 19388 13602 19440
rect 14734 19388 14740 19440
rect 14792 19388 14798 19440
rect 15028 19428 15056 19468
rect 15378 19456 15384 19468
rect 15436 19496 15442 19508
rect 15841 19499 15899 19505
rect 15841 19496 15853 19499
rect 15436 19468 15853 19496
rect 15436 19456 15442 19468
rect 15841 19465 15853 19468
rect 15887 19465 15899 19499
rect 17954 19496 17960 19508
rect 15841 19459 15899 19465
rect 16592 19468 17960 19496
rect 14936 19400 15056 19428
rect 14752 19301 14780 19388
rect 14936 19369 14964 19400
rect 15102 19388 15108 19440
rect 15160 19388 15166 19440
rect 15930 19388 15936 19440
rect 15988 19428 15994 19440
rect 15988 19400 16252 19428
rect 15988 19388 15994 19400
rect 14921 19363 14979 19369
rect 14921 19329 14933 19363
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15120 19360 15148 19388
rect 15838 19360 15844 19372
rect 15120 19332 15844 19360
rect 15120 19301 15148 19332
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 12032 19264 12173 19292
rect 12032 19252 12038 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 12345 19295 12403 19301
rect 12345 19261 12357 19295
rect 12391 19261 12403 19295
rect 12345 19255 12403 19261
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 14737 19295 14795 19301
rect 14737 19261 14749 19295
rect 14783 19261 14795 19295
rect 14737 19255 14795 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 15101 19295 15159 19301
rect 15101 19261 15113 19295
rect 15147 19261 15159 19295
rect 15101 19255 15159 19261
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19292 15347 19295
rect 15933 19295 15991 19301
rect 15335 19264 15893 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 12066 19224 12072 19236
rect 11900 19196 12072 19224
rect 6748 19128 7788 19156
rect 8110 19116 8116 19168
rect 8168 19156 8174 19168
rect 8754 19156 8760 19168
rect 8168 19128 8760 19156
rect 8168 19116 8174 19128
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 10870 19156 10876 19168
rect 10831 19128 10876 19156
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11900 19156 11928 19196
rect 12066 19184 12072 19196
rect 12124 19184 12130 19236
rect 11204 19128 11928 19156
rect 11204 19116 11210 19128
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 12360 19156 12388 19255
rect 13078 19184 13084 19236
rect 13136 19224 13142 19236
rect 14274 19224 14280 19236
rect 13136 19196 14280 19224
rect 13136 19184 13142 19196
rect 14274 19184 14280 19196
rect 14332 19184 14338 19236
rect 14918 19184 14924 19236
rect 14976 19224 14982 19236
rect 15028 19224 15056 19255
rect 14976 19196 15056 19224
rect 14976 19184 14982 19196
rect 12894 19156 12900 19168
rect 12216 19128 12388 19156
rect 12855 19128 12900 19156
rect 12216 19116 12222 19128
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 14550 19156 14556 19168
rect 14511 19128 14556 19156
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 15865 19156 15893 19264
rect 15933 19261 15945 19295
rect 15979 19292 15991 19295
rect 16114 19292 16120 19304
rect 15979 19264 16120 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16224 19224 16252 19400
rect 16592 19360 16620 19468
rect 17954 19456 17960 19468
rect 18012 19496 18018 19508
rect 18598 19496 18604 19508
rect 18012 19468 18604 19496
rect 18012 19456 18018 19468
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19496 20223 19499
rect 21174 19496 21180 19508
rect 20211 19468 21180 19496
rect 20211 19465 20223 19468
rect 20165 19459 20223 19465
rect 21174 19456 21180 19468
rect 21232 19496 21238 19508
rect 21232 19468 21588 19496
rect 21232 19456 21238 19468
rect 17126 19428 17132 19440
rect 16776 19400 17132 19428
rect 16776 19369 16804 19400
rect 17126 19388 17132 19400
rect 17184 19388 17190 19440
rect 17310 19388 17316 19440
rect 17368 19428 17374 19440
rect 19242 19428 19248 19440
rect 17368 19400 19248 19428
rect 17368 19388 17374 19400
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 19337 19431 19395 19437
rect 19337 19397 19349 19431
rect 19383 19428 19395 19431
rect 20346 19428 20352 19440
rect 19383 19400 20352 19428
rect 19383 19397 19395 19400
rect 19337 19391 19395 19397
rect 16500 19332 16620 19360
rect 16761 19363 16819 19369
rect 16500 19301 16528 19332
rect 16761 19329 16773 19363
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 17221 19363 17279 19369
rect 16899 19332 17172 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19261 16543 19295
rect 16666 19292 16672 19304
rect 16627 19264 16672 19292
rect 16485 19255 16543 19261
rect 16666 19252 16672 19264
rect 16724 19252 16730 19304
rect 17034 19292 17040 19304
rect 16995 19264 17040 19292
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 17144 19290 17172 19332
rect 17221 19329 17233 19363
rect 17267 19360 17279 19363
rect 17681 19363 17739 19369
rect 17267 19332 17632 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 17604 19292 17632 19332
rect 17681 19329 17693 19363
rect 17727 19360 17739 19363
rect 17862 19360 17868 19372
rect 17727 19332 17868 19360
rect 17727 19329 17739 19332
rect 17681 19323 17739 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 17957 19363 18015 19369
rect 17957 19329 17969 19363
rect 18003 19360 18015 19363
rect 18506 19360 18512 19372
rect 18003 19332 18512 19360
rect 18003 19329 18015 19332
rect 17957 19323 18015 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 17144 19262 17356 19290
rect 17604 19264 17724 19292
rect 16574 19224 16580 19236
rect 16224 19196 16580 19224
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 17328 19224 17356 19262
rect 17586 19224 17592 19236
rect 17328 19196 17592 19224
rect 17586 19184 17592 19196
rect 17644 19184 17650 19236
rect 17696 19224 17724 19264
rect 18598 19224 18604 19236
rect 17696 19196 18604 19224
rect 18598 19184 18604 19196
rect 18656 19184 18662 19236
rect 15930 19156 15936 19168
rect 15865 19128 15936 19156
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 17310 19156 17316 19168
rect 16448 19128 17316 19156
rect 16448 19116 16454 19128
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17494 19116 17500 19168
rect 17552 19156 17558 19168
rect 17770 19156 17776 19168
rect 17552 19128 17776 19156
rect 17552 19116 17558 19128
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 17862 19116 17868 19168
rect 17920 19156 17926 19168
rect 19352 19156 19380 19391
rect 20346 19388 20352 19400
rect 20404 19388 20410 19440
rect 21560 19360 21588 19468
rect 22002 19456 22008 19508
rect 22060 19496 22066 19508
rect 22373 19499 22431 19505
rect 22373 19496 22385 19499
rect 22060 19468 22385 19496
rect 22060 19456 22066 19468
rect 22373 19465 22385 19468
rect 22419 19465 22431 19499
rect 30742 19496 30748 19508
rect 22373 19459 22431 19465
rect 26344 19468 30748 19496
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21560 19332 22017 19360
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 23124 19332 23428 19360
rect 20254 19252 20260 19304
rect 20312 19292 20318 19304
rect 20312 19264 21128 19292
rect 20312 19252 20318 19264
rect 17920 19128 19380 19156
rect 21100 19156 21128 19264
rect 21266 19252 21272 19304
rect 21324 19301 21330 19304
rect 21324 19292 21336 19301
rect 21545 19295 21603 19301
rect 21324 19264 21369 19292
rect 21324 19255 21336 19264
rect 21545 19261 21557 19295
rect 21591 19292 21603 19295
rect 22278 19292 22284 19304
rect 21591 19264 22284 19292
rect 21591 19261 21603 19264
rect 21545 19255 21603 19261
rect 21324 19252 21330 19255
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 22370 19252 22376 19304
rect 22428 19252 22434 19304
rect 22738 19252 22744 19304
rect 22796 19292 22802 19304
rect 23124 19301 23152 19332
rect 23109 19295 23167 19301
rect 23109 19292 23121 19295
rect 22796 19264 23121 19292
rect 22796 19252 22802 19264
rect 23109 19261 23121 19264
rect 23155 19261 23167 19295
rect 23290 19292 23296 19304
rect 23251 19264 23296 19292
rect 23109 19255 23167 19261
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 23400 19292 23428 19332
rect 23474 19320 23480 19372
rect 23532 19360 23538 19372
rect 23842 19360 23848 19372
rect 23532 19332 23848 19360
rect 23532 19320 23538 19332
rect 23842 19320 23848 19332
rect 23900 19360 23906 19372
rect 24673 19363 24731 19369
rect 24673 19360 24685 19363
rect 23900 19332 24685 19360
rect 23900 19320 23906 19332
rect 24673 19329 24685 19332
rect 24719 19329 24731 19363
rect 24673 19323 24731 19329
rect 23750 19292 23756 19304
rect 23400 19264 23756 19292
rect 23750 19252 23756 19264
rect 23808 19252 23814 19304
rect 24394 19292 24400 19304
rect 24355 19264 24400 19292
rect 24394 19252 24400 19264
rect 24452 19252 24458 19304
rect 25590 19252 25596 19304
rect 25648 19292 25654 19304
rect 26237 19295 26295 19301
rect 26237 19292 26249 19295
rect 25648 19264 26249 19292
rect 25648 19252 25654 19264
rect 26237 19261 26249 19264
rect 26283 19261 26295 19295
rect 26237 19255 26295 19261
rect 22388 19224 22416 19252
rect 23201 19227 23259 19233
rect 23201 19224 23213 19227
rect 22388 19196 23213 19224
rect 23201 19193 23213 19196
rect 23247 19193 23259 19227
rect 26344 19224 26372 19468
rect 30742 19456 30748 19468
rect 30800 19456 30806 19508
rect 28166 19428 28172 19440
rect 27448 19400 28172 19428
rect 27338 19360 27344 19372
rect 27299 19332 27344 19360
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 27448 19369 27476 19400
rect 28166 19388 28172 19400
rect 28224 19428 28230 19440
rect 32232 19428 32260 19536
rect 32320 19428 33120 19442
rect 28224 19400 28672 19428
rect 32232 19400 33120 19428
rect 28224 19388 28230 19400
rect 28644 19369 28672 19400
rect 32320 19386 33120 19400
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19329 27491 19363
rect 28537 19363 28595 19369
rect 28537 19360 28549 19363
rect 27433 19323 27491 19329
rect 27540 19332 28549 19360
rect 27065 19295 27123 19301
rect 27065 19261 27077 19295
rect 27111 19261 27123 19295
rect 27246 19292 27252 19304
rect 27207 19264 27252 19292
rect 27065 19255 27123 19261
rect 23201 19187 23259 19193
rect 26068 19196 26372 19224
rect 27080 19224 27108 19255
rect 27246 19252 27252 19264
rect 27304 19252 27310 19304
rect 27356 19292 27384 19320
rect 27540 19292 27568 19332
rect 28537 19329 28549 19332
rect 28583 19329 28595 19363
rect 28537 19323 28595 19329
rect 28629 19363 28687 19369
rect 28629 19329 28641 19363
rect 28675 19329 28687 19363
rect 28629 19323 28687 19329
rect 28902 19320 28908 19372
rect 28960 19360 28966 19372
rect 30466 19360 30472 19372
rect 28960 19332 30472 19360
rect 28960 19320 28966 19332
rect 30466 19320 30472 19332
rect 30524 19320 30530 19372
rect 27356 19264 27568 19292
rect 27617 19295 27675 19301
rect 27617 19261 27629 19295
rect 27663 19261 27675 19295
rect 27617 19255 27675 19261
rect 27522 19224 27528 19236
rect 27080 19196 27528 19224
rect 22373 19159 22431 19165
rect 22373 19156 22385 19159
rect 21100 19128 22385 19156
rect 17920 19116 17926 19128
rect 22373 19125 22385 19128
rect 22419 19125 22431 19159
rect 22554 19156 22560 19168
rect 22515 19128 22560 19156
rect 22373 19119 22431 19125
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 22922 19116 22928 19168
rect 22980 19156 22986 19168
rect 25498 19156 25504 19168
rect 22980 19128 25504 19156
rect 22980 19116 22986 19128
rect 25498 19116 25504 19128
rect 25556 19156 25562 19168
rect 26068 19156 26096 19196
rect 27522 19184 27528 19196
rect 27580 19184 27586 19236
rect 27632 19224 27660 19255
rect 27706 19252 27712 19304
rect 27764 19292 27770 19304
rect 28261 19295 28319 19301
rect 28261 19292 28273 19295
rect 27764 19264 28273 19292
rect 27764 19252 27770 19264
rect 28261 19261 28273 19264
rect 28307 19292 28319 19295
rect 28350 19292 28356 19304
rect 28307 19264 28356 19292
rect 28307 19261 28319 19264
rect 28261 19255 28319 19261
rect 28350 19252 28356 19264
rect 28408 19252 28414 19304
rect 28445 19295 28503 19301
rect 28445 19261 28457 19295
rect 28491 19261 28503 19295
rect 28445 19255 28503 19261
rect 28460 19224 28488 19255
rect 28718 19252 28724 19304
rect 28776 19292 28782 19304
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28776 19264 28825 19292
rect 28776 19252 28782 19264
rect 28813 19261 28825 19264
rect 28859 19261 28871 19295
rect 28813 19255 28871 19261
rect 28994 19252 29000 19304
rect 29052 19292 29058 19304
rect 29549 19295 29607 19301
rect 29549 19292 29561 19295
rect 29052 19264 29561 19292
rect 29052 19252 29058 19264
rect 29549 19261 29561 19264
rect 29595 19261 29607 19295
rect 29549 19255 29607 19261
rect 30650 19224 30656 19236
rect 27632 19196 30656 19224
rect 30650 19184 30656 19196
rect 30708 19184 30714 19236
rect 25556 19128 26096 19156
rect 26145 19159 26203 19165
rect 25556 19116 25562 19128
rect 26145 19125 26157 19159
rect 26191 19156 26203 19159
rect 26326 19156 26332 19168
rect 26191 19128 26332 19156
rect 26191 19125 26203 19128
rect 26145 19119 26203 19125
rect 26326 19116 26332 19128
rect 26384 19116 26390 19168
rect 27798 19156 27804 19168
rect 27759 19128 27804 19156
rect 27798 19116 27804 19128
rect 27856 19116 27862 19168
rect 28810 19116 28816 19168
rect 28868 19156 28874 19168
rect 28997 19159 29055 19165
rect 28997 19156 29009 19159
rect 28868 19128 29009 19156
rect 28868 19116 28874 19128
rect 28997 19125 29009 19128
rect 29043 19125 29055 19159
rect 28997 19119 29055 19125
rect 29730 19116 29736 19168
rect 29788 19156 29794 19168
rect 30374 19156 30380 19168
rect 29788 19128 30380 19156
rect 29788 19116 29794 19128
rect 30374 19116 30380 19128
rect 30432 19156 30438 19168
rect 30837 19159 30895 19165
rect 30837 19156 30849 19159
rect 30432 19128 30849 19156
rect 30432 19116 30438 19128
rect 30837 19125 30849 19128
rect 30883 19125 30895 19159
rect 30837 19119 30895 19125
rect 1104 19066 32016 19088
rect 1104 19014 11253 19066
rect 11305 19014 11317 19066
rect 11369 19014 11381 19066
rect 11433 19014 11445 19066
rect 11497 19014 11509 19066
rect 11561 19014 21557 19066
rect 21609 19014 21621 19066
rect 21673 19014 21685 19066
rect 21737 19014 21749 19066
rect 21801 19014 21813 19066
rect 21865 19014 32016 19066
rect 1104 18992 32016 19014
rect 2222 18952 2228 18964
rect 1504 18924 2228 18952
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 1504 18825 1532 18924
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 2777 18955 2835 18961
rect 2777 18921 2789 18955
rect 2823 18952 2835 18955
rect 3050 18952 3056 18964
rect 2823 18924 3056 18952
rect 2823 18921 2835 18924
rect 2777 18915 2835 18921
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3292 18924 3801 18952
rect 3292 18912 3298 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 4430 18952 4436 18964
rect 4391 18924 4436 18952
rect 3789 18915 3847 18921
rect 4430 18912 4436 18924
rect 4488 18952 4494 18964
rect 6822 18952 6828 18964
rect 4488 18924 5580 18952
rect 6783 18924 6828 18952
rect 4488 18912 4494 18924
rect 2130 18884 2136 18896
rect 1780 18856 2136 18884
rect 1489 18819 1547 18825
rect 1489 18816 1501 18819
rect 1452 18788 1501 18816
rect 1452 18776 1458 18788
rect 1489 18785 1501 18788
rect 1535 18785 1547 18819
rect 1670 18816 1676 18828
rect 1631 18788 1676 18816
rect 1489 18779 1547 18785
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 1780 18760 1808 18856
rect 2130 18844 2136 18856
rect 2188 18844 2194 18896
rect 2314 18844 2320 18896
rect 2372 18884 2378 18896
rect 5552 18884 5580 18924
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 7650 18952 7656 18964
rect 7611 18924 7656 18952
rect 7650 18912 7656 18924
rect 7708 18952 7714 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 7708 18924 8493 18952
rect 7708 18912 7714 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 8481 18915 8539 18921
rect 8941 18955 8999 18961
rect 8941 18921 8953 18955
rect 8987 18952 8999 18955
rect 9122 18952 9128 18964
rect 8987 18924 9128 18952
rect 8987 18921 8999 18924
rect 8941 18915 8999 18921
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 13078 18952 13084 18964
rect 10652 18924 13084 18952
rect 10652 18912 10658 18924
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 13354 18912 13360 18964
rect 13412 18952 13418 18964
rect 13817 18955 13875 18961
rect 13817 18952 13829 18955
rect 13412 18924 13829 18952
rect 13412 18912 13418 18924
rect 13817 18921 13829 18924
rect 13863 18921 13875 18955
rect 13817 18915 13875 18921
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 15286 18952 15292 18964
rect 14148 18924 15292 18952
rect 14148 18912 14154 18924
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 15470 18912 15476 18964
rect 15528 18952 15534 18964
rect 15657 18955 15715 18961
rect 15657 18952 15669 18955
rect 15528 18924 15669 18952
rect 15528 18912 15534 18924
rect 15657 18921 15669 18924
rect 15703 18921 15715 18955
rect 15657 18915 15715 18921
rect 16666 18912 16672 18964
rect 16724 18912 16730 18964
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 18322 18952 18328 18964
rect 17736 18924 18328 18952
rect 17736 18912 17742 18924
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19300 18924 19717 18952
rect 19300 18912 19306 18924
rect 19705 18921 19717 18924
rect 19751 18921 19763 18955
rect 19705 18915 19763 18921
rect 6733 18887 6791 18893
rect 6733 18884 6745 18887
rect 2372 18856 2912 18884
rect 2372 18844 2378 18856
rect 2038 18816 2044 18828
rect 1999 18788 2044 18816
rect 2038 18776 2044 18788
rect 2096 18776 2102 18828
rect 2682 18816 2688 18828
rect 2643 18788 2688 18816
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 2884 18825 2912 18856
rect 4356 18856 5488 18884
rect 5552 18856 6745 18884
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18785 2927 18819
rect 2869 18779 2927 18785
rect 3234 18776 3240 18828
rect 3292 18816 3298 18828
rect 3602 18816 3608 18828
rect 3292 18788 3608 18816
rect 3292 18776 3298 18788
rect 3602 18776 3608 18788
rect 3660 18776 3666 18828
rect 3878 18816 3884 18828
rect 3839 18788 3884 18816
rect 3878 18776 3884 18788
rect 3936 18776 3942 18828
rect 4246 18776 4252 18828
rect 4304 18816 4310 18828
rect 4356 18825 4384 18856
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 4304 18788 4353 18816
rect 4304 18776 4310 18788
rect 4341 18785 4353 18788
rect 4387 18785 4399 18819
rect 4341 18779 4399 18785
rect 4525 18819 4583 18825
rect 4525 18785 4537 18819
rect 4571 18816 4583 18819
rect 4614 18816 4620 18828
rect 4571 18788 4620 18816
rect 4571 18785 4583 18788
rect 4525 18779 4583 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 5258 18816 5264 18828
rect 5219 18788 5264 18816
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5460 18825 5488 18856
rect 6733 18853 6745 18856
rect 6779 18853 6791 18887
rect 8110 18884 8116 18896
rect 6733 18847 6791 18853
rect 8036 18856 8116 18884
rect 8036 18828 8064 18856
rect 8110 18844 8116 18856
rect 8168 18844 8174 18896
rect 9668 18887 9726 18893
rect 9668 18853 9680 18887
rect 9714 18884 9726 18887
rect 10870 18884 10876 18896
rect 9714 18856 10876 18884
rect 9714 18853 9726 18856
rect 9668 18847 9726 18853
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11790 18844 11796 18896
rect 11848 18884 11854 18896
rect 12342 18884 12348 18896
rect 11848 18856 12348 18884
rect 11848 18844 11854 18856
rect 12342 18844 12348 18856
rect 12400 18844 12406 18896
rect 12704 18887 12762 18893
rect 12704 18853 12716 18887
rect 12750 18884 12762 18887
rect 12894 18884 12900 18896
rect 12750 18856 12900 18884
rect 12750 18853 12762 18856
rect 12704 18847 12762 18853
rect 12894 18844 12900 18856
rect 12952 18844 12958 18896
rect 16684 18884 16712 18912
rect 19334 18884 19340 18896
rect 16684 18856 19340 18884
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 19720 18884 19748 18915
rect 19794 18912 19800 18964
rect 19852 18952 19858 18964
rect 20898 18952 20904 18964
rect 19852 18924 20383 18952
rect 20859 18924 20904 18952
rect 19852 18912 19858 18924
rect 20355 18884 20383 18924
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 21910 18952 21916 18964
rect 21871 18924 21916 18952
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 22462 18912 22468 18964
rect 22520 18952 22526 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 22520 18924 22569 18952
rect 22520 18912 22526 18924
rect 22557 18921 22569 18924
rect 22603 18921 22615 18955
rect 22557 18915 22615 18921
rect 23566 18912 23572 18964
rect 23624 18952 23630 18964
rect 23624 18924 23704 18952
rect 23624 18912 23630 18924
rect 21450 18884 21456 18896
rect 19720 18856 20300 18884
rect 20355 18856 21456 18884
rect 5353 18819 5411 18825
rect 5353 18785 5365 18819
rect 5399 18785 5411 18819
rect 5460 18819 5524 18825
rect 5460 18788 5478 18819
rect 5353 18779 5411 18785
rect 5466 18785 5478 18788
rect 5512 18785 5524 18819
rect 5466 18779 5524 18785
rect 5629 18819 5687 18825
rect 5629 18785 5641 18819
rect 5675 18816 5687 18819
rect 5810 18816 5816 18828
rect 5675 18788 5816 18816
rect 5675 18785 5687 18788
rect 5629 18779 5687 18785
rect 1762 18748 1768 18760
rect 1723 18720 1768 18748
rect 1762 18708 1768 18720
rect 1820 18708 1826 18760
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18748 1915 18751
rect 1946 18748 1952 18760
rect 1903 18720 1952 18748
rect 1903 18717 1915 18720
rect 1857 18711 1915 18717
rect 1946 18708 1952 18720
rect 2004 18708 2010 18760
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 2774 18748 2780 18760
rect 2372 18720 2780 18748
rect 2372 18708 2378 18720
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 5381 18748 5409 18779
rect 5810 18776 5816 18788
rect 5868 18776 5874 18828
rect 7006 18776 7012 18828
rect 7064 18816 7070 18828
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 7064 18788 7573 18816
rect 7064 18776 7070 18788
rect 7561 18785 7573 18788
rect 7607 18816 7619 18819
rect 7650 18816 7656 18828
rect 7607 18788 7656 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 7745 18819 7803 18825
rect 7745 18785 7757 18819
rect 7791 18816 7803 18819
rect 7834 18816 7840 18828
rect 7791 18788 7840 18816
rect 7791 18785 7803 18788
rect 7745 18779 7803 18785
rect 6914 18748 6920 18760
rect 4856 18720 5409 18748
rect 6875 18720 6920 18748
rect 4856 18708 4862 18720
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 7760 18748 7788 18779
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 8018 18776 8024 18828
rect 8076 18776 8082 18828
rect 8202 18776 8208 18828
rect 8260 18816 8266 18828
rect 8573 18819 8631 18825
rect 8573 18816 8585 18819
rect 8260 18788 8585 18816
rect 8260 18776 8266 18788
rect 8573 18785 8585 18788
rect 8619 18785 8631 18819
rect 8573 18779 8631 18785
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 11238 18816 11244 18828
rect 11020 18788 11244 18816
rect 11020 18776 11026 18788
rect 11238 18776 11244 18788
rect 11296 18776 11302 18828
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 13446 18816 13452 18828
rect 11655 18788 13452 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 7524 18720 7788 18748
rect 8389 18751 8447 18757
rect 7524 18708 7530 18720
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 8938 18748 8944 18760
rect 8435 18720 8944 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 8938 18708 8944 18720
rect 8996 18708 9002 18760
rect 9398 18748 9404 18760
rect 9359 18720 9404 18748
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 11146 18748 11152 18760
rect 10928 18720 11152 18748
rect 10928 18708 10934 18720
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 3326 18640 3332 18692
rect 3384 18680 3390 18692
rect 7834 18680 7840 18692
rect 3384 18652 7840 18680
rect 3384 18640 3390 18652
rect 7834 18640 7840 18652
rect 7892 18640 7898 18692
rect 10962 18640 10968 18692
rect 11020 18680 11026 18692
rect 11624 18680 11652 18779
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 14366 18776 14372 18828
rect 14424 18776 14430 18828
rect 14550 18825 14556 18828
rect 14544 18816 14556 18825
rect 14511 18788 14556 18816
rect 14544 18779 14556 18788
rect 14550 18776 14556 18779
rect 14608 18776 14614 18828
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 15930 18816 15936 18828
rect 14976 18788 15936 18816
rect 14976 18776 14982 18788
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 16298 18776 16304 18828
rect 16356 18816 16362 18828
rect 16669 18819 16727 18825
rect 16669 18816 16681 18819
rect 16356 18788 16681 18816
rect 16356 18776 16362 18788
rect 16669 18785 16681 18788
rect 16715 18785 16727 18819
rect 16850 18816 16856 18828
rect 16811 18788 16856 18816
rect 16669 18779 16727 18785
rect 12342 18708 12348 18760
rect 12400 18748 12406 18760
rect 12437 18751 12495 18757
rect 12437 18748 12449 18751
rect 12400 18720 12449 18748
rect 12400 18708 12406 18720
rect 12437 18717 12449 18720
rect 12483 18717 12495 18751
rect 12437 18711 12495 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14384 18748 14412 18776
rect 14323 18720 14412 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 11020 18652 11652 18680
rect 11020 18640 11026 18652
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 1670 18612 1676 18624
rect 1544 18584 1676 18612
rect 1544 18572 1550 18584
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 2222 18612 2228 18624
rect 2183 18584 2228 18612
rect 2222 18572 2228 18584
rect 2280 18572 2286 18624
rect 4985 18615 5043 18621
rect 4985 18581 4997 18615
rect 5031 18612 5043 18615
rect 5166 18612 5172 18624
rect 5031 18584 5172 18612
rect 5031 18581 5043 18584
rect 4985 18575 5043 18581
rect 5166 18572 5172 18584
rect 5224 18572 5230 18624
rect 6365 18615 6423 18621
rect 6365 18581 6377 18615
rect 6411 18612 6423 18615
rect 6454 18612 6460 18624
rect 6411 18584 6460 18612
rect 6411 18581 6423 18584
rect 6365 18575 6423 18581
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 8110 18572 8116 18624
rect 8168 18612 8174 18624
rect 8754 18612 8760 18624
rect 8168 18584 8760 18612
rect 8168 18572 8174 18584
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 10502 18572 10508 18624
rect 10560 18612 10566 18624
rect 10781 18615 10839 18621
rect 10781 18612 10793 18615
rect 10560 18584 10793 18612
rect 10560 18572 10566 18584
rect 10781 18581 10793 18584
rect 10827 18581 10839 18615
rect 14292 18612 14320 18711
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15838 18748 15844 18760
rect 15344 18720 15844 18748
rect 15344 18708 15350 18720
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 16684 18748 16712 18779
rect 16850 18776 16856 18788
rect 16908 18776 16914 18828
rect 17037 18819 17095 18825
rect 17037 18785 17049 18819
rect 17083 18816 17095 18819
rect 17218 18816 17224 18828
rect 17083 18788 17224 18816
rect 17083 18785 17095 18788
rect 17037 18779 17095 18785
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 17310 18776 17316 18828
rect 17368 18816 17374 18828
rect 17773 18819 17831 18825
rect 17512 18816 17724 18818
rect 17773 18816 17785 18819
rect 17368 18790 17785 18816
rect 17368 18788 17540 18790
rect 17696 18788 17785 18790
rect 17368 18776 17374 18788
rect 17773 18785 17785 18788
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 17873 18809 17931 18815
rect 17873 18775 17885 18809
rect 17919 18806 17931 18809
rect 17919 18775 17939 18806
rect 18138 18776 18144 18828
rect 18196 18816 18202 18828
rect 18598 18825 18604 18828
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 18196 18788 18337 18816
rect 18196 18776 18202 18788
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 18592 18816 18604 18825
rect 18559 18788 18604 18816
rect 18325 18779 18383 18785
rect 18592 18779 18604 18788
rect 18598 18776 18604 18779
rect 18656 18776 18662 18828
rect 18874 18776 18880 18828
rect 18932 18816 18938 18828
rect 18932 18788 19380 18816
rect 18932 18776 18938 18788
rect 17873 18769 17939 18775
rect 17126 18748 17132 18760
rect 16684 18720 17132 18748
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17911 18748 17939 18769
rect 17911 18720 18368 18748
rect 18340 18692 18368 18720
rect 16574 18640 16580 18692
rect 16632 18680 16638 18692
rect 16942 18680 16948 18692
rect 16632 18652 16948 18680
rect 16632 18640 16638 18652
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 17218 18640 17224 18692
rect 17276 18640 17282 18692
rect 18322 18640 18328 18692
rect 18380 18640 18386 18692
rect 19352 18680 19380 18788
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 20162 18816 20168 18828
rect 19484 18788 20168 18816
rect 19484 18776 19490 18788
rect 20162 18776 20168 18788
rect 20220 18776 20226 18828
rect 20272 18816 20300 18856
rect 21450 18844 21456 18856
rect 21508 18844 21514 18896
rect 23676 18884 23704 18924
rect 24578 18912 24584 18964
rect 24636 18952 24642 18964
rect 24636 18924 26004 18952
rect 24636 18912 24642 18924
rect 23676 18856 24900 18884
rect 20346 18816 20352 18828
rect 20272 18788 20352 18816
rect 20346 18776 20352 18788
rect 20404 18816 20410 18828
rect 20717 18819 20775 18825
rect 20404 18788 20497 18816
rect 20404 18776 20410 18788
rect 20717 18785 20729 18819
rect 20763 18816 20775 18819
rect 22002 18816 22008 18828
rect 20763 18788 22008 18816
rect 20763 18785 20775 18788
rect 20717 18779 20775 18785
rect 22002 18776 22008 18788
rect 22060 18776 22066 18828
rect 22738 18816 22744 18828
rect 22699 18788 22744 18816
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 23385 18819 23443 18825
rect 23385 18785 23397 18819
rect 23431 18816 23443 18819
rect 23474 18816 23480 18828
rect 23431 18788 23480 18816
rect 23431 18785 23443 18788
rect 23385 18779 23443 18785
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 23676 18825 23704 18856
rect 24872 18825 24900 18856
rect 25976 18825 26004 18924
rect 27798 18912 27804 18964
rect 27856 18952 27862 18964
rect 27856 18924 29040 18952
rect 27856 18912 27862 18924
rect 27154 18844 27160 18896
rect 27212 18884 27218 18896
rect 28074 18884 28080 18896
rect 27212 18856 28080 18884
rect 27212 18844 27218 18856
rect 28074 18844 28080 18856
rect 28132 18844 28138 18896
rect 28810 18844 28816 18896
rect 28868 18893 28874 18896
rect 28868 18884 28880 18893
rect 29012 18884 29040 18924
rect 30650 18912 30656 18964
rect 30708 18952 30714 18964
rect 30929 18955 30987 18961
rect 30929 18952 30941 18955
rect 30708 18924 30941 18952
rect 30708 18912 30714 18924
rect 30929 18921 30941 18924
rect 30975 18921 30987 18955
rect 30929 18915 30987 18921
rect 29794 18887 29852 18893
rect 29794 18884 29806 18887
rect 28868 18856 28913 18884
rect 29012 18856 29806 18884
rect 28868 18847 28880 18856
rect 29794 18853 29806 18856
rect 29840 18853 29852 18887
rect 29794 18847 29852 18853
rect 28868 18844 28874 18847
rect 23569 18819 23627 18825
rect 23569 18785 23581 18819
rect 23615 18785 23627 18819
rect 23569 18779 23627 18785
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18785 23719 18819
rect 23661 18779 23719 18785
rect 23937 18819 23995 18825
rect 23937 18785 23949 18819
rect 23983 18816 23995 18819
rect 24857 18819 24915 18825
rect 23983 18788 24808 18816
rect 23983 18785 23995 18788
rect 23937 18779 23995 18785
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 20441 18751 20499 18757
rect 20441 18748 20453 18751
rect 19668 18720 20453 18748
rect 19668 18708 19674 18720
rect 20441 18717 20453 18720
rect 20487 18717 20499 18751
rect 20441 18711 20499 18717
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18748 20591 18751
rect 20806 18748 20812 18760
rect 20579 18720 20812 18748
rect 20579 18717 20591 18720
rect 20533 18711 20591 18717
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 23584 18748 23612 18779
rect 20956 18720 23612 18748
rect 23753 18751 23811 18757
rect 20956 18708 20962 18720
rect 23753 18717 23765 18751
rect 23799 18717 23811 18751
rect 24578 18748 24584 18760
rect 24539 18720 24584 18748
rect 23753 18711 23811 18717
rect 23658 18680 23664 18692
rect 19352 18652 23664 18680
rect 23658 18640 23664 18652
rect 23716 18640 23722 18692
rect 23768 18680 23796 18711
rect 24578 18708 24584 18720
rect 24636 18708 24642 18760
rect 24780 18748 24808 18788
rect 24857 18785 24869 18819
rect 24903 18785 24915 18819
rect 24857 18779 24915 18785
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18816 26019 18819
rect 27982 18816 27988 18828
rect 26007 18788 27988 18816
rect 26007 18785 26019 18788
rect 25961 18779 26019 18785
rect 27982 18776 27988 18788
rect 28040 18776 28046 18828
rect 29089 18819 29147 18825
rect 29089 18785 29101 18819
rect 29135 18816 29147 18819
rect 29549 18819 29607 18825
rect 29549 18816 29561 18819
rect 29135 18788 29561 18816
rect 29135 18785 29147 18788
rect 29089 18779 29147 18785
rect 29549 18785 29561 18788
rect 29595 18816 29607 18819
rect 29638 18816 29644 18828
rect 29595 18788 29644 18816
rect 29595 18785 29607 18788
rect 29549 18779 29607 18785
rect 29638 18776 29644 18788
rect 29696 18776 29702 18828
rect 26418 18748 26424 18760
rect 24780 18720 26424 18748
rect 26418 18708 26424 18720
rect 26476 18708 26482 18760
rect 26326 18680 26332 18692
rect 23768 18652 26332 18680
rect 26326 18640 26332 18652
rect 26384 18640 26390 18692
rect 16114 18612 16120 18624
rect 14292 18584 16120 18612
rect 10781 18575 10839 18581
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16758 18612 16764 18624
rect 16719 18584 16764 18612
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 17236 18612 17264 18640
rect 17310 18612 17316 18624
rect 17236 18584 17316 18612
rect 17310 18572 17316 18584
rect 17368 18572 17374 18624
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 17586 18612 17592 18624
rect 17460 18584 17592 18612
rect 17460 18572 17466 18584
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 19794 18612 19800 18624
rect 19392 18584 19800 18612
rect 19392 18572 19398 18584
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 19886 18572 19892 18624
rect 19944 18612 19950 18624
rect 23106 18612 23112 18624
rect 19944 18584 23112 18612
rect 19944 18572 19950 18584
rect 23106 18572 23112 18584
rect 23164 18572 23170 18624
rect 24121 18615 24179 18621
rect 24121 18581 24133 18615
rect 24167 18612 24179 18615
rect 25314 18612 25320 18624
rect 24167 18584 25320 18612
rect 24167 18581 24179 18584
rect 24121 18575 24179 18581
rect 25314 18572 25320 18584
rect 25372 18572 25378 18624
rect 27154 18612 27160 18624
rect 27115 18584 27160 18612
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 27709 18615 27767 18621
rect 27709 18581 27721 18615
rect 27755 18612 27767 18615
rect 28718 18612 28724 18624
rect 27755 18584 28724 18612
rect 27755 18581 27767 18584
rect 27709 18575 27767 18581
rect 28718 18572 28724 18584
rect 28776 18572 28782 18624
rect 1104 18522 32016 18544
rect 1104 18470 6102 18522
rect 6154 18470 6166 18522
rect 6218 18470 6230 18522
rect 6282 18470 6294 18522
rect 6346 18470 6358 18522
rect 6410 18470 16405 18522
rect 16457 18470 16469 18522
rect 16521 18470 16533 18522
rect 16585 18470 16597 18522
rect 16649 18470 16661 18522
rect 16713 18470 26709 18522
rect 26761 18470 26773 18522
rect 26825 18470 26837 18522
rect 26889 18470 26901 18522
rect 26953 18470 26965 18522
rect 27017 18470 32016 18522
rect 1104 18448 32016 18470
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 5626 18408 5632 18420
rect 4120 18380 5632 18408
rect 4120 18368 4126 18380
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 8110 18408 8116 18420
rect 7576 18380 7972 18408
rect 8071 18380 8116 18408
rect 5534 18300 5540 18352
rect 5592 18340 5598 18352
rect 7576 18340 7604 18380
rect 7944 18340 7972 18380
rect 8110 18368 8116 18380
rect 8168 18368 8174 18420
rect 8846 18368 8852 18420
rect 8904 18408 8910 18420
rect 9398 18408 9404 18420
rect 8904 18380 9404 18408
rect 8904 18368 8910 18380
rect 9398 18368 9404 18380
rect 9456 18408 9462 18420
rect 11054 18408 11060 18420
rect 9456 18380 11060 18408
rect 9456 18368 9462 18380
rect 11054 18368 11060 18380
rect 11112 18408 11118 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 11112 18380 11805 18408
rect 11112 18368 11118 18380
rect 11793 18377 11805 18380
rect 11839 18408 11851 18411
rect 12342 18408 12348 18420
rect 11839 18380 12348 18408
rect 11839 18377 11851 18380
rect 11793 18371 11851 18377
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 13998 18368 14004 18420
rect 14056 18408 14062 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 14056 18380 14105 18408
rect 14056 18368 14062 18380
rect 14093 18377 14105 18380
rect 14139 18408 14151 18411
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 14139 18380 14841 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 14829 18377 14841 18380
rect 14875 18377 14887 18411
rect 15930 18408 15936 18420
rect 14829 18371 14887 18377
rect 14933 18380 15700 18408
rect 15891 18380 15936 18408
rect 8757 18343 8815 18349
rect 8757 18340 8769 18343
rect 5592 18312 7604 18340
rect 7668 18312 7880 18340
rect 7944 18312 8769 18340
rect 5592 18300 5598 18312
rect 4982 18272 4988 18284
rect 4943 18244 4988 18272
rect 4982 18232 4988 18244
rect 5040 18232 5046 18284
rect 5626 18272 5632 18284
rect 5276 18244 5632 18272
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2510 18207 2568 18213
rect 2510 18204 2522 18207
rect 2280 18176 2522 18204
rect 2280 18164 2286 18176
rect 2510 18173 2522 18176
rect 2556 18173 2568 18207
rect 2510 18167 2568 18173
rect 2682 18164 2688 18216
rect 2740 18204 2746 18216
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2740 18176 2789 18204
rect 2740 18164 2746 18176
rect 2777 18173 2789 18176
rect 2823 18173 2835 18207
rect 2777 18167 2835 18173
rect 4522 18164 4528 18216
rect 4580 18204 4586 18216
rect 5276 18213 5304 18244
rect 5626 18232 5632 18244
rect 5684 18272 5690 18284
rect 6730 18272 6736 18284
rect 5684 18244 6736 18272
rect 5684 18232 5690 18244
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 7668 18272 7696 18312
rect 6963 18244 7696 18272
rect 7852 18272 7880 18312
rect 8757 18309 8769 18312
rect 8803 18309 8815 18343
rect 8757 18303 8815 18309
rect 9122 18300 9128 18352
rect 9180 18340 9186 18352
rect 9490 18340 9496 18352
rect 9180 18312 9496 18340
rect 9180 18300 9186 18312
rect 9490 18300 9496 18312
rect 9548 18300 9554 18352
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 12802 18340 12808 18352
rect 10284 18312 12808 18340
rect 10284 18300 10290 18312
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 13357 18343 13415 18349
rect 13357 18340 13369 18343
rect 13320 18312 13369 18340
rect 13320 18300 13326 18312
rect 13357 18309 13369 18312
rect 13403 18340 13415 18343
rect 14933 18340 14961 18380
rect 15562 18340 15568 18352
rect 13403 18312 14961 18340
rect 15523 18312 15568 18340
rect 13403 18309 13415 18312
rect 13357 18303 13415 18309
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 15672 18340 15700 18380
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16206 18368 16212 18420
rect 16264 18408 16270 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 16264 18380 16957 18408
rect 16264 18368 16270 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 16945 18371 17003 18377
rect 17129 18411 17187 18417
rect 17129 18377 17141 18411
rect 17175 18408 17187 18411
rect 17310 18408 17316 18420
rect 17175 18380 17316 18408
rect 17175 18377 17187 18380
rect 17129 18371 17187 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 17681 18411 17739 18417
rect 17681 18377 17693 18411
rect 17727 18408 17739 18411
rect 18322 18408 18328 18420
rect 17727 18380 18328 18408
rect 17727 18377 17739 18380
rect 17681 18371 17739 18377
rect 18322 18368 18328 18380
rect 18380 18408 18386 18420
rect 19242 18408 19248 18420
rect 18380 18380 19248 18408
rect 18380 18368 18386 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 20438 18408 20444 18420
rect 19352 18380 20444 18408
rect 15672 18312 16712 18340
rect 9858 18272 9864 18284
rect 7852 18244 9168 18272
rect 9771 18244 9864 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 5169 18207 5227 18213
rect 5169 18204 5181 18207
rect 4580 18176 5181 18204
rect 4580 18164 4586 18176
rect 5169 18173 5181 18176
rect 5215 18173 5227 18207
rect 5169 18167 5227 18173
rect 5261 18207 5319 18213
rect 5261 18173 5273 18207
rect 5307 18173 5319 18207
rect 5261 18167 5319 18173
rect 6089 18207 6147 18213
rect 6089 18173 6101 18207
rect 6135 18204 6147 18207
rect 6454 18204 6460 18216
rect 6135 18176 6460 18204
rect 6135 18173 6147 18176
rect 6089 18167 6147 18173
rect 6454 18164 6460 18176
rect 6512 18164 6518 18216
rect 7006 18204 7012 18216
rect 6967 18176 7012 18204
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 7466 18204 7472 18216
rect 7427 18176 7472 18204
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 7668 18213 7696 18244
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 7926 18204 7932 18216
rect 7883 18176 7932 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 7760 18136 7788 18167
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 8478 18164 8484 18216
rect 8536 18204 8542 18216
rect 9140 18213 9168 18244
rect 9858 18232 9864 18244
rect 9916 18272 9922 18284
rect 9916 18244 13584 18272
rect 9916 18232 9922 18244
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 8536 18176 8953 18204
rect 8536 18164 8542 18176
rect 8941 18173 8953 18176
rect 8987 18173 8999 18207
rect 8941 18167 8999 18173
rect 9125 18207 9183 18213
rect 9125 18173 9137 18207
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 10410 18164 10416 18216
rect 10468 18204 10474 18216
rect 11698 18204 11704 18216
rect 10468 18176 11704 18204
rect 10468 18164 10474 18176
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 13556 18213 13584 18244
rect 14642 18232 14648 18284
rect 14700 18272 14706 18284
rect 14918 18272 14924 18284
rect 14700 18244 14924 18272
rect 14700 18232 14706 18244
rect 14918 18232 14924 18244
rect 14976 18232 14982 18284
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 16577 18275 16635 18281
rect 16577 18272 16589 18275
rect 15528 18244 16589 18272
rect 15528 18232 15534 18244
rect 16577 18241 16589 18244
rect 16623 18241 16635 18275
rect 16684 18272 16712 18312
rect 17218 18300 17224 18352
rect 17276 18340 17282 18352
rect 19352 18340 19380 18380
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 27062 18408 27068 18420
rect 23716 18380 27068 18408
rect 23716 18368 23722 18380
rect 27062 18368 27068 18380
rect 27120 18368 27126 18420
rect 28902 18408 28908 18420
rect 27172 18380 28908 18408
rect 19886 18340 19892 18352
rect 17276 18312 19380 18340
rect 19444 18312 19892 18340
rect 17276 18300 17282 18312
rect 18601 18275 18659 18281
rect 16684 18244 18460 18272
rect 16577 18235 16635 18241
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 13998 18204 14004 18216
rect 13587 18176 14004 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 13998 18164 14004 18176
rect 14056 18164 14062 18216
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14148 18176 16436 18204
rect 14148 18164 14154 18176
rect 8294 18136 8300 18148
rect 2792 18108 8300 18136
rect 2792 18080 2820 18108
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 8757 18139 8815 18145
rect 8757 18105 8769 18139
rect 8803 18136 8815 18139
rect 9490 18136 9496 18148
rect 8803 18108 9496 18136
rect 8803 18105 8815 18108
rect 8757 18099 8815 18105
rect 9490 18096 9496 18108
rect 9548 18136 9554 18148
rect 10505 18139 10563 18145
rect 10505 18136 10517 18139
rect 9548 18108 10517 18136
rect 9548 18096 9554 18108
rect 10505 18105 10517 18108
rect 10551 18136 10563 18139
rect 14182 18136 14188 18148
rect 10551 18108 14188 18136
rect 10551 18105 10563 18108
rect 10505 18099 10563 18105
rect 14182 18096 14188 18108
rect 14240 18096 14246 18148
rect 14737 18139 14795 18145
rect 14737 18105 14749 18139
rect 14783 18136 14795 18139
rect 14918 18136 14924 18148
rect 14783 18108 14924 18136
rect 14783 18105 14795 18108
rect 14737 18099 14795 18105
rect 14918 18096 14924 18108
rect 14976 18136 14982 18148
rect 16298 18136 16304 18148
rect 14976 18108 16304 18136
rect 14976 18096 14982 18108
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 1397 18071 1455 18077
rect 1397 18037 1409 18071
rect 1443 18068 1455 18071
rect 1486 18068 1492 18080
rect 1443 18040 1492 18068
rect 1443 18037 1455 18040
rect 1397 18031 1455 18037
rect 1486 18028 1492 18040
rect 1544 18068 1550 18080
rect 2038 18068 2044 18080
rect 1544 18040 2044 18068
rect 1544 18028 1550 18040
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 2774 18028 2780 18080
rect 2832 18028 2838 18080
rect 3973 18071 4031 18077
rect 3973 18037 3985 18071
rect 4019 18068 4031 18071
rect 4062 18068 4068 18080
rect 4019 18040 4068 18068
rect 4019 18037 4031 18040
rect 3973 18031 4031 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4433 18071 4491 18077
rect 4433 18068 4445 18071
rect 4304 18040 4445 18068
rect 4304 18028 4310 18040
rect 4433 18037 4445 18040
rect 4479 18068 4491 18071
rect 4706 18068 4712 18080
rect 4479 18040 4712 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 4985 18071 5043 18077
rect 4985 18037 4997 18071
rect 5031 18068 5043 18071
rect 5718 18068 5724 18080
rect 5031 18040 5724 18068
rect 5031 18037 5043 18040
rect 4985 18031 5043 18037
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 5994 18068 6000 18080
rect 5955 18040 6000 18068
rect 5994 18028 6000 18040
rect 6052 18028 6058 18080
rect 8202 18028 8208 18080
rect 8260 18068 8266 18080
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 8260 18040 9045 18068
rect 8260 18028 8266 18040
rect 9033 18037 9045 18040
rect 9079 18037 9091 18071
rect 9033 18031 9091 18037
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 11606 18068 11612 18080
rect 10100 18040 11612 18068
rect 10100 18028 10106 18040
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 11790 18028 11796 18080
rect 11848 18068 11854 18080
rect 12713 18071 12771 18077
rect 12713 18068 12725 18071
rect 11848 18040 12725 18068
rect 11848 18028 11854 18040
rect 12713 18037 12725 18040
rect 12759 18037 12771 18071
rect 12713 18031 12771 18037
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 14550 18068 14556 18080
rect 12860 18040 14556 18068
rect 12860 18028 12866 18040
rect 14550 18028 14556 18040
rect 14608 18068 14614 18080
rect 15746 18068 15752 18080
rect 14608 18040 15752 18068
rect 14608 18028 14614 18040
rect 15746 18028 15752 18040
rect 15804 18068 15810 18080
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 15804 18040 15945 18068
rect 15804 18028 15810 18040
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 16117 18071 16175 18077
rect 16117 18037 16129 18071
rect 16163 18068 16175 18071
rect 16206 18068 16212 18080
rect 16163 18040 16212 18068
rect 16163 18037 16175 18040
rect 16117 18031 16175 18037
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16408 18068 16436 18176
rect 16666 18164 16672 18216
rect 16724 18164 16730 18216
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17218 18204 17224 18216
rect 16816 18176 17224 18204
rect 16816 18164 16822 18176
rect 17218 18164 17224 18176
rect 17276 18164 17282 18216
rect 17678 18204 17684 18216
rect 17420 18176 17684 18204
rect 16684 18136 16712 18164
rect 17420 18136 17448 18176
rect 17678 18164 17684 18176
rect 17736 18164 17742 18216
rect 17770 18164 17776 18216
rect 17828 18204 17834 18216
rect 18141 18207 18199 18213
rect 18141 18204 18153 18207
rect 17828 18176 18153 18204
rect 17828 18164 17834 18176
rect 18141 18173 18153 18176
rect 18187 18173 18199 18207
rect 18322 18204 18328 18216
rect 18283 18176 18328 18204
rect 18141 18167 18199 18173
rect 18322 18164 18328 18176
rect 18380 18164 18386 18216
rect 18432 18204 18460 18244
rect 18601 18241 18613 18275
rect 18647 18272 18659 18275
rect 18690 18272 18696 18284
rect 18647 18244 18696 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 19444 18272 19472 18312
rect 19886 18300 19892 18312
rect 19944 18300 19950 18352
rect 20530 18300 20536 18352
rect 20588 18340 20594 18352
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 20588 18312 22017 18340
rect 20588 18300 20594 18312
rect 22005 18309 22017 18312
rect 22051 18340 22063 18343
rect 27172 18340 27200 18380
rect 28902 18368 28908 18380
rect 28960 18368 28966 18420
rect 22051 18312 27200 18340
rect 22051 18309 22063 18312
rect 22005 18303 22063 18309
rect 18800 18244 19472 18272
rect 19613 18275 19671 18281
rect 18800 18204 18828 18244
rect 19613 18241 19625 18275
rect 19659 18272 19671 18275
rect 20806 18272 20812 18284
rect 19659 18244 20812 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 24397 18275 24455 18281
rect 24397 18272 24409 18275
rect 23124 18244 24409 18272
rect 18432 18176 18828 18204
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19334 18204 19340 18216
rect 19291 18176 19340 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 19429 18207 19487 18213
rect 19429 18173 19441 18207
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18204 19579 18207
rect 19794 18204 19800 18216
rect 19567 18176 19656 18204
rect 19755 18176 19800 18204
rect 19567 18173 19579 18176
rect 19521 18167 19579 18173
rect 18046 18136 18052 18148
rect 16684 18108 17448 18136
rect 17512 18108 18052 18136
rect 16945 18071 17003 18077
rect 16945 18068 16957 18071
rect 16408 18040 16957 18068
rect 16945 18037 16957 18040
rect 16991 18068 17003 18071
rect 17512 18068 17540 18108
rect 18046 18096 18052 18108
rect 18104 18096 18110 18148
rect 18506 18096 18512 18148
rect 18564 18136 18570 18148
rect 18693 18139 18751 18145
rect 18693 18136 18705 18139
rect 18564 18108 18705 18136
rect 18564 18096 18570 18108
rect 18693 18105 18705 18108
rect 18739 18136 18751 18139
rect 18874 18136 18880 18148
rect 18739 18108 18880 18136
rect 18739 18105 18751 18108
rect 18693 18099 18751 18105
rect 18874 18096 18880 18108
rect 18932 18096 18938 18148
rect 19150 18096 19156 18148
rect 19208 18136 19214 18148
rect 19444 18136 19472 18167
rect 19628 18148 19656 18176
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 20441 18207 20499 18213
rect 20441 18173 20453 18207
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 21177 18207 21235 18213
rect 21177 18173 21189 18207
rect 21223 18204 21235 18207
rect 21223 18176 22094 18204
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 19208 18108 19472 18136
rect 19208 18096 19214 18108
rect 19610 18096 19616 18148
rect 19668 18096 19674 18148
rect 20456 18136 20484 18167
rect 22066 18148 22094 18176
rect 22646 18164 22652 18216
rect 22704 18204 22710 18216
rect 23124 18213 23152 18244
rect 24397 18241 24409 18244
rect 24443 18241 24455 18275
rect 24397 18235 24455 18241
rect 25332 18244 27660 18272
rect 23109 18207 23167 18213
rect 23109 18204 23121 18207
rect 22704 18176 23121 18204
rect 22704 18164 22710 18176
rect 23109 18173 23121 18176
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23382 18164 23388 18216
rect 23440 18204 23446 18216
rect 25332 18213 25360 18244
rect 25317 18207 25375 18213
rect 25317 18204 25329 18207
rect 23440 18176 25329 18204
rect 23440 18164 23446 18176
rect 25317 18173 25329 18176
rect 25363 18173 25375 18207
rect 27525 18207 27583 18213
rect 27525 18204 27537 18207
rect 25317 18167 25375 18173
rect 26620 18176 27537 18204
rect 19812 18108 20484 18136
rect 21729 18139 21787 18145
rect 16991 18040 17540 18068
rect 16991 18037 17003 18040
rect 16945 18031 17003 18037
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 19812 18068 19840 18108
rect 21729 18105 21741 18139
rect 21775 18105 21787 18139
rect 21729 18099 21787 18105
rect 17644 18040 19840 18068
rect 17644 18028 17650 18040
rect 19886 18028 19892 18080
rect 19944 18068 19950 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19944 18040 19993 18068
rect 19944 18028 19950 18040
rect 19981 18037 19993 18040
rect 20027 18037 20039 18071
rect 20530 18068 20536 18080
rect 20491 18040 20536 18068
rect 19981 18031 20039 18037
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 21082 18028 21088 18080
rect 21140 18068 21146 18080
rect 21744 18068 21772 18099
rect 22002 18096 22008 18148
rect 22060 18136 22094 18148
rect 23750 18136 23756 18148
rect 22060 18108 23756 18136
rect 22060 18096 22066 18108
rect 23750 18096 23756 18108
rect 23808 18096 23814 18148
rect 22186 18068 22192 18080
rect 21140 18040 22192 18068
rect 21140 18028 21146 18040
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 22830 18028 22836 18080
rect 22888 18068 22894 18080
rect 22925 18071 22983 18077
rect 22925 18068 22937 18071
rect 22888 18040 22937 18068
rect 22888 18028 22894 18040
rect 22925 18037 22937 18040
rect 22971 18037 22983 18071
rect 23658 18068 23664 18080
rect 23619 18040 23664 18068
rect 22925 18031 22983 18037
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 26234 18068 26240 18080
rect 25280 18040 26240 18068
rect 25280 18028 25286 18040
rect 26234 18028 26240 18040
rect 26292 18068 26298 18080
rect 26620 18077 26648 18176
rect 27525 18173 27537 18176
rect 27571 18173 27583 18207
rect 27632 18204 27660 18244
rect 28994 18204 29000 18216
rect 27632 18176 29000 18204
rect 27525 18167 27583 18173
rect 28994 18164 29000 18176
rect 29052 18164 29058 18216
rect 29730 18164 29736 18216
rect 29788 18204 29794 18216
rect 29917 18207 29975 18213
rect 29917 18204 29929 18207
rect 29788 18176 29929 18204
rect 29788 18164 29794 18176
rect 29917 18173 29929 18176
rect 29963 18173 29975 18207
rect 29917 18167 29975 18173
rect 27798 18145 27804 18148
rect 27792 18099 27804 18145
rect 27856 18136 27862 18148
rect 30184 18139 30242 18145
rect 27856 18108 27892 18136
rect 27798 18096 27804 18099
rect 27856 18096 27862 18108
rect 30184 18105 30196 18139
rect 30230 18136 30242 18139
rect 30282 18136 30288 18148
rect 30230 18108 30288 18136
rect 30230 18105 30242 18108
rect 30184 18099 30242 18105
rect 30282 18096 30288 18108
rect 30340 18096 30346 18148
rect 26605 18071 26663 18077
rect 26605 18068 26617 18071
rect 26292 18040 26617 18068
rect 26292 18028 26298 18040
rect 26605 18037 26617 18040
rect 26651 18037 26663 18071
rect 26605 18031 26663 18037
rect 27246 18028 27252 18080
rect 27304 18068 27310 18080
rect 28905 18071 28963 18077
rect 28905 18068 28917 18071
rect 27304 18040 28917 18068
rect 27304 18028 27310 18040
rect 28905 18037 28917 18040
rect 28951 18037 28963 18071
rect 28905 18031 28963 18037
rect 30466 18028 30472 18080
rect 30524 18068 30530 18080
rect 31294 18068 31300 18080
rect 30524 18040 31300 18068
rect 30524 18028 30530 18040
rect 31294 18028 31300 18040
rect 31352 18028 31358 18080
rect 1104 17978 32016 18000
rect 1104 17926 11253 17978
rect 11305 17926 11317 17978
rect 11369 17926 11381 17978
rect 11433 17926 11445 17978
rect 11497 17926 11509 17978
rect 11561 17926 21557 17978
rect 21609 17926 21621 17978
rect 21673 17926 21685 17978
rect 21737 17926 21749 17978
rect 21801 17926 21813 17978
rect 21865 17926 32016 17978
rect 1104 17904 32016 17926
rect 1946 17824 1952 17876
rect 2004 17824 2010 17876
rect 3878 17824 3884 17876
rect 3936 17864 3942 17876
rect 3973 17867 4031 17873
rect 3973 17864 3985 17867
rect 3936 17836 3985 17864
rect 3936 17824 3942 17836
rect 3973 17833 3985 17836
rect 4019 17833 4031 17867
rect 3973 17827 4031 17833
rect 1762 17796 1768 17808
rect 1688 17768 1768 17796
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 1486 17688 1492 17740
rect 1544 17728 1550 17740
rect 1688 17737 1716 17768
rect 1762 17756 1768 17768
rect 1820 17756 1826 17808
rect 1964 17796 1992 17824
rect 1872 17768 1992 17796
rect 2133 17799 2191 17805
rect 1581 17731 1639 17737
rect 1581 17728 1593 17731
rect 1544 17700 1593 17728
rect 1544 17688 1550 17700
rect 1581 17697 1593 17700
rect 1627 17697 1639 17731
rect 1581 17691 1639 17697
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17697 1731 17731
rect 1673 17691 1731 17697
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 1872 17660 1900 17768
rect 2133 17765 2145 17799
rect 2179 17796 2191 17799
rect 2838 17799 2896 17805
rect 2838 17796 2850 17799
rect 2179 17768 2850 17796
rect 2179 17765 2191 17768
rect 2133 17759 2191 17765
rect 2838 17765 2850 17768
rect 2884 17765 2896 17799
rect 3988 17796 4016 17827
rect 8202 17824 8208 17876
rect 8260 17873 8266 17876
rect 8260 17867 8279 17873
rect 8267 17833 8279 17867
rect 8386 17864 8392 17876
rect 8347 17836 8392 17864
rect 8260 17827 8279 17833
rect 8260 17824 8266 17827
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 10594 17864 10600 17876
rect 8496 17836 10600 17864
rect 4617 17799 4675 17805
rect 4617 17796 4629 17799
rect 3988 17768 4629 17796
rect 2838 17759 2896 17765
rect 4617 17765 4629 17768
rect 4663 17765 4675 17799
rect 4617 17759 4675 17765
rect 7926 17756 7932 17808
rect 7984 17796 7990 17808
rect 8021 17799 8079 17805
rect 8021 17796 8033 17799
rect 7984 17768 8033 17796
rect 7984 17756 7990 17768
rect 8021 17765 8033 17768
rect 8067 17765 8079 17799
rect 8021 17759 8079 17765
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2593 17731 2651 17737
rect 1995 17700 2553 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 1811 17632 1900 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 2525 17524 2553 17700
rect 2593 17697 2605 17731
rect 2639 17728 2651 17731
rect 2682 17728 2688 17740
rect 2639 17700 2688 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17728 5503 17731
rect 5626 17728 5632 17740
rect 5491 17700 5632 17728
rect 5491 17697 5503 17700
rect 5445 17691 5503 17697
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 6914 17728 6920 17740
rect 6875 17700 6920 17728
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5534 17620 5540 17672
rect 5592 17660 5598 17672
rect 8496 17660 8524 17836
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 11606 17824 11612 17876
rect 11664 17824 11670 17876
rect 12986 17824 12992 17876
rect 13044 17864 13050 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 13044 17836 13737 17864
rect 13044 17824 13050 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 18598 17864 18604 17876
rect 17000 17836 18604 17864
rect 17000 17824 17006 17836
rect 8662 17756 8668 17808
rect 8720 17796 8726 17808
rect 9217 17799 9275 17805
rect 9217 17796 9229 17799
rect 8720 17768 9229 17796
rect 8720 17756 8726 17768
rect 9217 17765 9229 17768
rect 9263 17765 9275 17799
rect 9217 17759 9275 17765
rect 9585 17799 9643 17805
rect 9585 17765 9597 17799
rect 9631 17796 9643 17799
rect 9858 17796 9864 17808
rect 9631 17768 9864 17796
rect 9631 17765 9643 17768
rect 9585 17759 9643 17765
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 10502 17756 10508 17808
rect 10560 17796 10566 17808
rect 11624 17796 11652 17824
rect 15746 17796 15752 17808
rect 10560 17768 11560 17796
rect 11624 17768 15752 17796
rect 10560 17756 10566 17768
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 10321 17731 10379 17737
rect 10321 17728 10333 17731
rect 10008 17700 10333 17728
rect 10008 17688 10014 17700
rect 10321 17697 10333 17700
rect 10367 17697 10379 17731
rect 10321 17691 10379 17697
rect 10410 17688 10416 17740
rect 10468 17688 10474 17740
rect 10704 17737 10732 17768
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17697 10747 17731
rect 10689 17691 10747 17697
rect 10870 17688 10876 17740
rect 10928 17728 10934 17740
rect 11532 17737 11560 17768
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 15933 17799 15991 17805
rect 15933 17765 15945 17799
rect 15979 17796 15991 17799
rect 16114 17796 16120 17808
rect 15979 17768 16120 17796
rect 15979 17765 15991 17768
rect 15933 17759 15991 17765
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 17126 17796 17132 17808
rect 17052 17768 17132 17796
rect 11517 17731 11575 17737
rect 10928 17700 10973 17728
rect 10928 17688 10934 17700
rect 11517 17697 11529 17731
rect 11563 17697 11575 17731
rect 12342 17728 12348 17740
rect 12303 17700 12348 17728
rect 11517 17691 11575 17697
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 12612 17731 12670 17737
rect 12612 17697 12624 17731
rect 12658 17728 12670 17731
rect 13078 17728 13084 17740
rect 12658 17700 13084 17728
rect 12658 17697 12670 17700
rect 12612 17691 12670 17697
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 14182 17728 14188 17740
rect 14095 17700 14188 17728
rect 14182 17688 14188 17700
rect 14240 17728 14246 17740
rect 15102 17728 15108 17740
rect 14240 17700 15108 17728
rect 14240 17688 14246 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 17052 17737 17080 17768
rect 17126 17756 17132 17768
rect 17184 17756 17190 17808
rect 17328 17737 17356 17836
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 18966 17824 18972 17876
rect 19024 17864 19030 17876
rect 19518 17864 19524 17876
rect 19024 17836 19524 17864
rect 19024 17824 19030 17836
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 20070 17864 20076 17876
rect 19983 17836 20076 17864
rect 17770 17796 17776 17808
rect 17731 17768 17776 17796
rect 17770 17756 17776 17768
rect 17828 17756 17834 17808
rect 18230 17796 18236 17808
rect 18191 17768 18236 17796
rect 18230 17756 18236 17768
rect 18288 17756 18294 17808
rect 19996 17805 20024 17836
rect 20070 17824 20076 17836
rect 20128 17864 20134 17876
rect 20622 17864 20628 17876
rect 20128 17836 20628 17864
rect 20128 17824 20134 17836
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 23014 17864 23020 17876
rect 20732 17836 23020 17864
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17765 20039 17799
rect 19981 17759 20039 17765
rect 20162 17756 20168 17808
rect 20220 17796 20226 17808
rect 20732 17796 20760 17836
rect 23014 17824 23020 17836
rect 23072 17864 23078 17876
rect 23382 17864 23388 17876
rect 23072 17836 23388 17864
rect 23072 17824 23078 17836
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 24210 17824 24216 17876
rect 24268 17864 24274 17876
rect 27709 17867 27767 17873
rect 24268 17836 27660 17864
rect 24268 17824 24274 17836
rect 27632 17808 27660 17836
rect 27709 17833 27721 17867
rect 27755 17864 27767 17867
rect 27798 17864 27804 17876
rect 27755 17836 27804 17864
rect 27755 17833 27767 17836
rect 27709 17827 27767 17833
rect 27798 17824 27804 17836
rect 27856 17824 27862 17876
rect 30834 17864 30840 17876
rect 28612 17836 30840 17864
rect 25314 17805 25320 17808
rect 24305 17799 24363 17805
rect 24305 17796 24317 17799
rect 20220 17768 20760 17796
rect 21008 17768 24317 17796
rect 20220 17756 20226 17768
rect 17037 17731 17095 17737
rect 17037 17697 17049 17731
rect 17083 17697 17095 17731
rect 17037 17691 17095 17697
rect 17221 17731 17279 17737
rect 17221 17697 17233 17731
rect 17267 17697 17279 17731
rect 17221 17691 17279 17697
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17697 17371 17731
rect 17586 17728 17592 17740
rect 17547 17700 17592 17728
rect 17313 17691 17371 17697
rect 5592 17632 8524 17660
rect 5592 17620 5598 17632
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 10042 17660 10048 17672
rect 9456 17632 10048 17660
rect 9456 17620 9462 17632
rect 10042 17620 10048 17632
rect 10100 17620 10106 17672
rect 10428 17660 10456 17688
rect 10505 17663 10563 17669
rect 10505 17660 10517 17663
rect 10428 17632 10517 17660
rect 10505 17629 10517 17632
rect 10551 17629 10563 17663
rect 10505 17623 10563 17629
rect 10597 17663 10655 17669
rect 10597 17629 10609 17663
rect 10643 17660 10655 17663
rect 11882 17660 11888 17672
rect 10643 17632 11888 17660
rect 10643 17629 10655 17632
rect 10597 17623 10655 17629
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 15470 17660 15476 17672
rect 13596 17632 15476 17660
rect 13596 17620 13602 17632
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 3878 17552 3884 17604
rect 3936 17592 3942 17604
rect 4433 17595 4491 17601
rect 4433 17592 4445 17595
rect 3936 17564 4445 17592
rect 3936 17552 3942 17564
rect 4433 17561 4445 17564
rect 4479 17561 4491 17595
rect 4433 17555 4491 17561
rect 6454 17552 6460 17604
rect 6512 17592 6518 17604
rect 6733 17595 6791 17601
rect 6733 17592 6745 17595
rect 6512 17564 6745 17592
rect 6512 17552 6518 17564
rect 6733 17561 6745 17564
rect 6779 17561 6791 17595
rect 6733 17555 6791 17561
rect 6914 17552 6920 17604
rect 6972 17592 6978 17604
rect 7190 17592 7196 17604
rect 6972 17564 7196 17592
rect 6972 17552 6978 17564
rect 7190 17552 7196 17564
rect 7248 17592 7254 17604
rect 7561 17595 7619 17601
rect 7561 17592 7573 17595
rect 7248 17564 7573 17592
rect 7248 17552 7254 17564
rect 7561 17561 7573 17564
rect 7607 17592 7619 17595
rect 10410 17592 10416 17604
rect 7607 17564 10416 17592
rect 7607 17561 7619 17564
rect 7561 17555 7619 17561
rect 10410 17552 10416 17564
rect 10468 17552 10474 17604
rect 10870 17552 10876 17604
rect 10928 17592 10934 17604
rect 16850 17592 16856 17604
rect 10928 17564 11744 17592
rect 10928 17552 10934 17564
rect 2866 17524 2872 17536
rect 2525 17496 2872 17524
rect 2866 17484 2872 17496
rect 2924 17524 2930 17536
rect 3896 17524 3924 17552
rect 5258 17524 5264 17536
rect 2924 17496 3924 17524
rect 5219 17496 5264 17524
rect 2924 17484 2930 17496
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 5353 17527 5411 17533
rect 5353 17493 5365 17527
rect 5399 17524 5411 17527
rect 5902 17524 5908 17536
rect 5399 17496 5908 17524
rect 5399 17493 5411 17496
rect 5353 17487 5411 17493
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 8205 17527 8263 17533
rect 8205 17524 8217 17527
rect 7892 17496 8217 17524
rect 7892 17484 7898 17496
rect 8205 17493 8217 17496
rect 8251 17493 8263 17527
rect 8205 17487 8263 17493
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 10137 17527 10195 17533
rect 10137 17524 10149 17527
rect 9640 17496 10149 17524
rect 9640 17484 9646 17496
rect 10137 17493 10149 17496
rect 10183 17493 10195 17527
rect 10137 17487 10195 17493
rect 10594 17484 10600 17536
rect 10652 17524 10658 17536
rect 11609 17527 11667 17533
rect 11609 17524 11621 17527
rect 10652 17496 11621 17524
rect 10652 17484 10658 17496
rect 11609 17493 11621 17496
rect 11655 17493 11667 17527
rect 11716 17524 11744 17564
rect 13280 17564 16856 17592
rect 13280 17524 13308 17564
rect 16850 17552 16856 17564
rect 16908 17552 16914 17604
rect 17236 17592 17264 17691
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 20346 17688 20352 17740
rect 20404 17728 20410 17740
rect 21008 17737 21036 17768
rect 24305 17765 24317 17768
rect 24351 17765 24363 17799
rect 24305 17759 24363 17765
rect 25308 17759 25320 17805
rect 25372 17796 25378 17808
rect 25372 17768 25408 17796
rect 25314 17756 25320 17759
rect 25372 17756 25378 17768
rect 25866 17756 25872 17808
rect 25924 17796 25930 17808
rect 25924 17768 27108 17796
rect 25924 17756 25930 17768
rect 20441 17731 20499 17737
rect 20441 17728 20453 17731
rect 20404 17700 20453 17728
rect 20404 17688 20410 17700
rect 20441 17697 20453 17700
rect 20487 17697 20499 17731
rect 20441 17691 20499 17697
rect 20625 17731 20683 17737
rect 20625 17697 20637 17731
rect 20671 17697 20683 17731
rect 20625 17691 20683 17697
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 20993 17731 21051 17737
rect 20763 17700 20944 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17660 17463 17663
rect 18046 17660 18052 17672
rect 17451 17632 18052 17660
rect 17451 17629 17463 17632
rect 17405 17623 17463 17629
rect 18046 17620 18052 17632
rect 18104 17620 18110 17672
rect 20530 17660 20536 17672
rect 19306 17632 20536 17660
rect 19306 17592 19334 17632
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 17236 17564 19334 17592
rect 19794 17552 19800 17604
rect 19852 17592 19858 17604
rect 20254 17592 20260 17604
rect 19852 17564 20260 17592
rect 19852 17552 19858 17564
rect 20254 17552 20260 17564
rect 20312 17592 20318 17604
rect 20640 17592 20668 17691
rect 20806 17660 20812 17672
rect 20767 17632 20812 17660
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 20916 17660 20944 17700
rect 20993 17697 21005 17731
rect 21039 17697 21051 17731
rect 22278 17728 22284 17740
rect 22239 17700 22284 17728
rect 20993 17691 21051 17697
rect 22278 17688 22284 17700
rect 22336 17688 22342 17740
rect 22554 17737 22560 17740
rect 22548 17691 22560 17737
rect 22612 17728 22618 17740
rect 24210 17728 24216 17740
rect 22612 17700 22648 17728
rect 24171 17700 24216 17728
rect 22554 17688 22560 17691
rect 22612 17688 22618 17700
rect 24210 17688 24216 17700
rect 24268 17688 24274 17740
rect 26510 17688 26516 17740
rect 26568 17728 26574 17740
rect 26973 17731 27031 17737
rect 26973 17728 26985 17731
rect 26568 17700 26985 17728
rect 26568 17688 26574 17700
rect 26973 17697 26985 17700
rect 27019 17697 27031 17731
rect 26973 17691 27031 17697
rect 21358 17660 21364 17672
rect 20916 17632 21364 17660
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 25041 17663 25099 17669
rect 25041 17629 25053 17663
rect 25087 17629 25099 17663
rect 25041 17623 25099 17629
rect 20312 17564 20668 17592
rect 20312 17552 20318 17564
rect 11716 17496 13308 17524
rect 11609 17487 11667 17493
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 18230 17524 18236 17536
rect 14516 17496 18236 17524
rect 14516 17484 14522 17496
rect 18230 17484 18236 17496
rect 18288 17524 18294 17536
rect 18506 17524 18512 17536
rect 18288 17496 18512 17524
rect 18288 17484 18294 17496
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 20990 17524 20996 17536
rect 18656 17496 20996 17524
rect 18656 17484 18662 17496
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 21174 17524 21180 17536
rect 21135 17496 21180 17524
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 23661 17527 23719 17533
rect 23661 17524 23673 17527
rect 22152 17496 23673 17524
rect 22152 17484 22158 17496
rect 23661 17493 23673 17496
rect 23707 17524 23719 17527
rect 23934 17524 23940 17536
rect 23707 17496 23940 17524
rect 23707 17493 23719 17496
rect 23661 17487 23719 17493
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 25056 17524 25084 17623
rect 27080 17592 27108 17768
rect 27246 17756 27252 17808
rect 27304 17796 27310 17808
rect 27304 17768 27568 17796
rect 27304 17756 27310 17768
rect 27540 17737 27568 17768
rect 27614 17756 27620 17808
rect 27672 17796 27678 17808
rect 28612 17805 28640 17836
rect 30834 17824 30840 17836
rect 30892 17824 30898 17876
rect 30926 17824 30932 17876
rect 30984 17864 30990 17876
rect 31297 17867 31355 17873
rect 31297 17864 31309 17867
rect 30984 17836 31309 17864
rect 30984 17824 30990 17836
rect 31297 17833 31309 17836
rect 31343 17833 31355 17867
rect 31297 17827 31355 17833
rect 28597 17799 28655 17805
rect 28597 17796 28609 17799
rect 27672 17768 28609 17796
rect 27672 17756 27678 17768
rect 28597 17765 28609 17768
rect 28643 17765 28655 17799
rect 28597 17759 28655 17765
rect 28813 17799 28871 17805
rect 28813 17765 28825 17799
rect 28859 17796 28871 17799
rect 28859 17768 29408 17796
rect 28859 17765 28871 17768
rect 28813 17759 28871 17765
rect 27157 17731 27215 17737
rect 27157 17697 27169 17731
rect 27203 17728 27215 17731
rect 27525 17731 27583 17737
rect 27203 17700 27476 17728
rect 27203 17697 27215 17700
rect 27157 17691 27215 17697
rect 27246 17660 27252 17672
rect 27207 17632 27252 17660
rect 27246 17620 27252 17632
rect 27304 17620 27310 17672
rect 27341 17663 27399 17669
rect 27341 17629 27353 17663
rect 27387 17629 27399 17663
rect 27448 17660 27476 17700
rect 27525 17697 27537 17731
rect 27571 17728 27583 17731
rect 29273 17731 29331 17737
rect 29273 17728 29285 17731
rect 27571 17700 29285 17728
rect 27571 17697 27583 17700
rect 27525 17691 27583 17697
rect 29273 17697 29285 17700
rect 29319 17697 29331 17731
rect 29273 17691 29331 17697
rect 27448 17632 28672 17660
rect 27341 17623 27399 17629
rect 27356 17592 27384 17623
rect 27080 17564 27384 17592
rect 28644 17536 28672 17632
rect 25222 17524 25228 17536
rect 25056 17496 25228 17524
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 26418 17524 26424 17536
rect 26379 17496 26424 17524
rect 26418 17484 26424 17496
rect 26476 17484 26482 17536
rect 28442 17524 28448 17536
rect 28403 17496 28448 17524
rect 28442 17484 28448 17496
rect 28500 17484 28506 17536
rect 28626 17524 28632 17536
rect 28587 17496 28632 17524
rect 28626 17484 28632 17496
rect 28684 17484 28690 17536
rect 29380 17533 29408 17768
rect 29914 17756 29920 17808
rect 29972 17796 29978 17808
rect 29972 17768 32352 17796
rect 29972 17756 29978 17768
rect 30190 17737 30196 17740
rect 30184 17691 30196 17737
rect 30248 17728 30254 17740
rect 30248 17700 30284 17728
rect 30190 17688 30196 17691
rect 30248 17688 30254 17700
rect 29730 17620 29736 17672
rect 29788 17660 29794 17672
rect 29917 17663 29975 17669
rect 29917 17660 29929 17663
rect 29788 17632 29929 17660
rect 29788 17620 29794 17632
rect 29917 17629 29929 17632
rect 29963 17629 29975 17663
rect 29917 17623 29975 17629
rect 29365 17527 29423 17533
rect 29365 17493 29377 17527
rect 29411 17524 29423 17527
rect 30650 17524 30656 17536
rect 29411 17496 30656 17524
rect 29411 17493 29423 17496
rect 29365 17487 29423 17493
rect 30650 17484 30656 17496
rect 30708 17484 30714 17536
rect 32324 17524 32352 17768
rect 32232 17496 32352 17524
rect 1104 17434 32016 17456
rect 0 17388 800 17402
rect 0 17360 888 17388
rect 1104 17382 6102 17434
rect 6154 17382 6166 17434
rect 6218 17382 6230 17434
rect 6282 17382 6294 17434
rect 6346 17382 6358 17434
rect 6410 17382 16405 17434
rect 16457 17382 16469 17434
rect 16521 17382 16533 17434
rect 16585 17382 16597 17434
rect 16649 17382 16661 17434
rect 16713 17382 26709 17434
rect 26761 17382 26773 17434
rect 26825 17382 26837 17434
rect 26889 17382 26901 17434
rect 26953 17382 26965 17434
rect 27017 17382 32016 17434
rect 1104 17360 32016 17382
rect 32232 17388 32260 17496
rect 32320 17388 33120 17402
rect 32232 17360 33120 17388
rect 0 17346 800 17360
rect 860 17116 888 17360
rect 32320 17346 33120 17360
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 2133 17323 2191 17329
rect 2133 17320 2145 17323
rect 1820 17292 2145 17320
rect 1820 17280 1826 17292
rect 2133 17289 2145 17292
rect 2179 17289 2191 17323
rect 2133 17283 2191 17289
rect 7469 17323 7527 17329
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 8478 17320 8484 17332
rect 7515 17292 8484 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 9398 17320 9404 17332
rect 9359 17292 9404 17320
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 10008 17292 11376 17320
rect 10008 17280 10014 17292
rect 1581 17255 1639 17261
rect 1581 17221 1593 17255
rect 1627 17252 1639 17255
rect 4062 17252 4068 17264
rect 1627 17224 4068 17252
rect 1627 17221 1639 17224
rect 1581 17215 1639 17221
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 5258 17212 5264 17264
rect 5316 17252 5322 17264
rect 5316 17224 5672 17252
rect 5316 17212 5322 17224
rect 3602 17144 3608 17196
rect 3660 17184 3666 17196
rect 3970 17184 3976 17196
rect 3660 17156 3976 17184
rect 3660 17144 3666 17156
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 5534 17184 5540 17196
rect 5491 17156 5540 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 5644 17184 5672 17224
rect 5994 17212 6000 17264
rect 6052 17252 6058 17264
rect 10962 17252 10968 17264
rect 6052 17224 6316 17252
rect 6052 17212 6058 17224
rect 6288 17193 6316 17224
rect 10244 17224 10968 17252
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 5644 17156 6101 17184
rect 6089 17153 6101 17156
rect 6135 17153 6147 17187
rect 6089 17147 6147 17153
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17153 6331 17187
rect 6273 17147 6331 17153
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 10244 17193 10272 17224
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 10229 17187 10287 17193
rect 9916 17156 10088 17184
rect 9916 17144 9922 17156
rect 2777 17119 2835 17125
rect 2777 17116 2789 17119
rect 860 17088 2789 17116
rect 2777 17085 2789 17088
rect 2823 17116 2835 17119
rect 3050 17116 3056 17128
rect 2823 17088 3056 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 4614 17116 4620 17128
rect 4575 17088 4620 17116
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 4798 17076 4804 17128
rect 4856 17116 4862 17128
rect 5350 17116 5356 17128
rect 4856 17088 5356 17116
rect 4856 17076 4862 17088
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 5718 17116 5724 17128
rect 5679 17088 5724 17116
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 6546 17116 6552 17128
rect 6507 17088 6552 17116
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 7377 17119 7435 17125
rect 7377 17085 7389 17119
rect 7423 17116 7435 17119
rect 7466 17116 7472 17128
rect 7423 17088 7472 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 9950 17116 9956 17128
rect 9911 17088 9956 17116
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 10060 17116 10088 17156
rect 10229 17153 10241 17187
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10870 17184 10876 17196
rect 10367 17156 10876 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 10060 17088 10149 17116
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 10505 17119 10563 17125
rect 10505 17106 10517 17119
rect 10551 17106 10563 17119
rect 10137 17079 10195 17085
rect 2225 17051 2283 17057
rect 2225 17017 2237 17051
rect 2271 17048 2283 17051
rect 3142 17048 3148 17060
rect 2271 17020 3148 17048
rect 2271 17017 2283 17020
rect 2225 17011 2283 17017
rect 3142 17008 3148 17020
rect 3200 17048 3206 17060
rect 5994 17048 6000 17060
rect 3200 17020 6000 17048
rect 3200 17008 3206 17020
rect 5994 17008 6000 17020
rect 6052 17048 6058 17060
rect 6454 17048 6460 17060
rect 6052 17020 6460 17048
rect 6052 17008 6058 17020
rect 6454 17008 6460 17020
rect 6512 17008 6518 17060
rect 8389 17051 8447 17057
rect 10502 17054 10508 17106
rect 10560 17054 10566 17106
rect 8389 17017 8401 17051
rect 8435 17048 8447 17051
rect 8435 17020 9674 17048
rect 8435 17017 8447 17020
rect 8389 17011 8447 17017
rect 2774 16940 2780 16992
rect 2832 16980 2838 16992
rect 2961 16983 3019 16989
rect 2961 16980 2973 16983
rect 2832 16952 2973 16980
rect 2832 16940 2838 16952
rect 2961 16949 2973 16952
rect 3007 16949 3019 16983
rect 2961 16943 3019 16949
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 3878 16980 3884 16992
rect 3476 16952 3884 16980
rect 3476 16940 3482 16952
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 4154 16980 4160 16992
rect 4115 16952 4160 16980
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 4709 16983 4767 16989
rect 4709 16949 4721 16983
rect 4755 16980 4767 16983
rect 5258 16980 5264 16992
rect 4755 16952 5264 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 9646 16980 9674 17020
rect 10612 16980 10640 17156
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11348 17125 11376 17292
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 12526 17320 12532 17332
rect 11664 17292 12532 17320
rect 11664 17280 11670 17292
rect 12526 17280 12532 17292
rect 12584 17320 12590 17332
rect 13078 17320 13084 17332
rect 12584 17292 12747 17320
rect 13039 17292 13084 17320
rect 12584 17280 12590 17292
rect 11882 17252 11888 17264
rect 11440 17224 11888 17252
rect 11440 17193 11468 17224
rect 11882 17212 11888 17224
rect 11940 17252 11946 17264
rect 11940 17224 12664 17252
rect 11940 17212 11946 17224
rect 12636 17196 12664 17224
rect 11425 17187 11483 17193
rect 11425 17153 11437 17187
rect 11471 17153 11483 17187
rect 11425 17147 11483 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 11606 17184 11612 17196
rect 11563 17156 11612 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 12618 17184 12624 17196
rect 12032 17156 12388 17184
rect 12579 17156 12624 17184
rect 12032 17144 12038 17156
rect 12360 17128 12388 17156
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 11112 17088 11161 17116
rect 11112 17076 11118 17088
rect 11149 17085 11161 17088
rect 11195 17085 11207 17119
rect 11149 17079 11207 17085
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17085 11391 17119
rect 11333 17079 11391 17085
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17116 11759 17119
rect 12066 17116 12072 17128
rect 11747 17088 12072 17116
rect 11747 17085 11759 17088
rect 11701 17079 11759 17085
rect 12066 17076 12072 17088
rect 12124 17076 12130 17128
rect 12342 17116 12348 17128
rect 12303 17088 12348 17116
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12719 17125 12747 17292
rect 13078 17280 13084 17292
rect 13136 17280 13142 17332
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 16758 17320 16764 17332
rect 15344 17292 16764 17320
rect 15344 17280 15350 17292
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 17218 17280 17224 17332
rect 17276 17320 17282 17332
rect 17494 17320 17500 17332
rect 17276 17292 17500 17320
rect 17276 17280 17282 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 18509 17323 18567 17329
rect 18509 17320 18521 17323
rect 17644 17292 18521 17320
rect 17644 17280 17650 17292
rect 18509 17289 18521 17292
rect 18555 17289 18567 17323
rect 18509 17283 18567 17289
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19300 17292 21772 17320
rect 19300 17280 19306 17292
rect 14274 17252 14280 17264
rect 14235 17224 14280 17252
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 14375 17224 18276 17252
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 14375 17184 14403 17224
rect 12860 17156 14403 17184
rect 12860 17144 12866 17156
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 16390 17184 16396 17196
rect 15528 17156 16396 17184
rect 15528 17144 15534 17156
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 17862 17184 17868 17196
rect 17144 17156 17868 17184
rect 17144 17128 17172 17156
rect 17862 17144 17868 17156
rect 17920 17184 17926 17196
rect 18141 17187 18199 17193
rect 18141 17184 18153 17187
rect 17920 17156 18153 17184
rect 17920 17144 17926 17156
rect 18141 17153 18153 17156
rect 18187 17153 18199 17187
rect 18248 17184 18276 17224
rect 18322 17212 18328 17264
rect 18380 17252 18386 17264
rect 18693 17255 18751 17261
rect 18693 17252 18705 17255
rect 18380 17224 18705 17252
rect 18380 17212 18386 17224
rect 18693 17221 18705 17224
rect 18739 17221 18751 17255
rect 21744 17252 21772 17292
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 24210 17320 24216 17332
rect 22520 17292 24216 17320
rect 22520 17280 22526 17292
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 30098 17320 30104 17332
rect 24320 17292 30104 17320
rect 24320 17252 24348 17292
rect 30098 17280 30104 17292
rect 30156 17280 30162 17332
rect 30282 17320 30288 17332
rect 30243 17292 30288 17320
rect 30282 17280 30288 17292
rect 30340 17280 30346 17332
rect 30650 17280 30656 17332
rect 30708 17320 30714 17332
rect 30708 17292 31064 17320
rect 30708 17280 30714 17292
rect 21744 17224 23152 17252
rect 18693 17215 18751 17221
rect 20530 17184 20536 17196
rect 18248 17156 20536 17184
rect 18141 17147 18199 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 12492 17088 12541 17116
rect 12492 17076 12498 17088
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 12713 17119 12771 17125
rect 12713 17085 12725 17119
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 12986 17116 12992 17128
rect 12943 17088 12992 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 14093 17119 14151 17125
rect 14093 17085 14105 17119
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 10689 17051 10747 17057
rect 10689 17017 10701 17051
rect 10735 17048 10747 17051
rect 14108 17048 14136 17079
rect 10735 17020 14136 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 11882 16980 11888 16992
rect 9646 16952 10640 16980
rect 11843 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 14292 16980 14320 17079
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 15105 17119 15163 17125
rect 15105 17116 15117 17119
rect 14424 17088 15117 17116
rect 14424 17076 14430 17088
rect 15105 17085 15117 17088
rect 15151 17085 15163 17119
rect 15105 17079 15163 17085
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17085 15347 17119
rect 15289 17079 15347 17085
rect 15565 17119 15623 17125
rect 15565 17085 15577 17119
rect 15611 17116 15623 17119
rect 16209 17119 16267 17125
rect 15611 17088 16160 17116
rect 15611 17085 15623 17088
rect 15565 17079 15623 17085
rect 14458 17008 14464 17060
rect 14516 17048 14522 17060
rect 14645 17051 14703 17057
rect 14645 17048 14657 17051
rect 14516 17020 14657 17048
rect 14516 17008 14522 17020
rect 14645 17017 14657 17020
rect 14691 17017 14703 17051
rect 14645 17011 14703 17017
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 15304 17048 15332 17079
rect 14792 17020 15332 17048
rect 14792 17008 14798 17020
rect 15470 17008 15476 17060
rect 15528 17048 15534 17060
rect 15657 17051 15715 17057
rect 15657 17048 15669 17051
rect 15528 17020 15669 17048
rect 15528 17008 15534 17020
rect 15657 17017 15669 17020
rect 15703 17048 15715 17051
rect 15838 17048 15844 17060
rect 15703 17020 15844 17048
rect 15703 17017 15715 17020
rect 15657 17011 15715 17017
rect 15838 17008 15844 17020
rect 15896 17008 15902 17060
rect 16132 17048 16160 17088
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 16298 17116 16304 17128
rect 16255 17088 16304 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 17126 17116 17132 17128
rect 16500 17088 16988 17116
rect 17087 17088 17132 17116
rect 16500 17048 16528 17088
rect 16132 17020 16528 17048
rect 16960 17048 16988 17088
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 17497 17119 17555 17125
rect 17497 17085 17509 17119
rect 17543 17116 17555 17119
rect 17586 17116 17592 17128
rect 17543 17088 17592 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 16960 17020 17172 17048
rect 17144 16992 17172 17020
rect 12032 16952 14320 16980
rect 12032 16940 12038 16952
rect 15746 16940 15752 16992
rect 15804 16980 15810 16992
rect 16393 16983 16451 16989
rect 16393 16980 16405 16983
rect 15804 16952 16405 16980
rect 15804 16940 15810 16952
rect 16393 16949 16405 16952
rect 16439 16949 16451 16983
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 16393 16943 16451 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17126 16940 17132 16992
rect 17184 16940 17190 16992
rect 17328 16980 17356 17079
rect 17420 17048 17448 17079
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17681 17119 17739 17125
rect 17681 17085 17693 17119
rect 17727 17116 17739 17119
rect 17954 17116 17960 17128
rect 17727 17088 17960 17116
rect 17727 17085 17739 17088
rect 17681 17079 17739 17085
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18782 17116 18788 17128
rect 18064 17088 18788 17116
rect 18064 17048 18092 17088
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 19429 17119 19487 17125
rect 19429 17085 19441 17119
rect 19475 17085 19487 17119
rect 19610 17116 19616 17128
rect 19571 17088 19616 17116
rect 19429 17079 19487 17085
rect 18506 17048 18512 17060
rect 17420 17020 18092 17048
rect 18419 17020 18512 17048
rect 18506 17008 18512 17020
rect 18564 17048 18570 17060
rect 19058 17048 19064 17060
rect 18564 17020 19064 17048
rect 18564 17008 18570 17020
rect 19058 17008 19064 17020
rect 19116 17008 19122 17060
rect 19444 17048 19472 17079
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 20165 17119 20223 17125
rect 20165 17085 20177 17119
rect 20211 17116 20223 17119
rect 20438 17116 20444 17128
rect 20211 17088 20444 17116
rect 20211 17085 20223 17088
rect 20165 17079 20223 17085
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 20806 17116 20812 17128
rect 20767 17088 20812 17116
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 23124 17125 23152 17224
rect 23308 17224 24348 17252
rect 24397 17255 24455 17261
rect 23308 17125 23336 17224
rect 24397 17221 24409 17255
rect 24443 17221 24455 17255
rect 24397 17215 24455 17221
rect 23385 17187 23443 17193
rect 23385 17153 23397 17187
rect 23431 17184 23443 17187
rect 23842 17184 23848 17196
rect 23431 17156 23848 17184
rect 23431 17153 23443 17156
rect 23385 17147 23443 17153
rect 23842 17144 23848 17156
rect 23900 17144 23906 17196
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17085 23167 17119
rect 23109 17079 23167 17085
rect 23293 17119 23351 17125
rect 23293 17085 23305 17119
rect 23339 17085 23351 17119
rect 23293 17079 23351 17085
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 23661 17119 23719 17125
rect 23532 17088 23577 17116
rect 23532 17076 23538 17088
rect 23661 17085 23673 17119
rect 23707 17116 23719 17119
rect 24412 17116 24440 17215
rect 28626 17212 28632 17264
rect 28684 17252 28690 17264
rect 30837 17255 30895 17261
rect 30837 17252 30849 17255
rect 28684 17224 30849 17252
rect 28684 17212 28690 17224
rect 30837 17221 30849 17224
rect 30883 17221 30895 17255
rect 30837 17215 30895 17221
rect 27154 17184 27160 17196
rect 26252 17156 27160 17184
rect 23707 17088 24440 17116
rect 23707 17085 23719 17088
rect 23661 17079 23719 17085
rect 19518 17048 19524 17060
rect 19444 17020 19524 17048
rect 19518 17008 19524 17020
rect 19576 17008 19582 17060
rect 20349 17051 20407 17057
rect 20349 17017 20361 17051
rect 20395 17017 20407 17051
rect 20349 17011 20407 17017
rect 21076 17051 21134 17057
rect 21076 17017 21088 17051
rect 21122 17048 21134 17051
rect 21450 17048 21456 17060
rect 21122 17020 21456 17048
rect 21122 17017 21134 17020
rect 21076 17011 21134 17017
rect 17770 16980 17776 16992
rect 17328 16952 17776 16980
rect 17770 16940 17776 16952
rect 17828 16980 17834 16992
rect 18874 16980 18880 16992
rect 17828 16952 18880 16980
rect 17828 16940 17834 16952
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 20364 16980 20392 17011
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 23198 17008 23204 17060
rect 23256 17048 23262 17060
rect 23676 17048 23704 17079
rect 25222 17076 25228 17128
rect 25280 17116 25286 17128
rect 25777 17119 25835 17125
rect 25777 17116 25789 17119
rect 25280 17088 25789 17116
rect 25280 17076 25286 17088
rect 25777 17085 25789 17088
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 26142 17076 26148 17128
rect 26200 17116 26206 17128
rect 26252 17125 26280 17156
rect 27154 17144 27160 17156
rect 27212 17184 27218 17196
rect 27525 17187 27583 17193
rect 27525 17184 27537 17187
rect 27212 17156 27537 17184
rect 27212 17144 27218 17156
rect 27525 17153 27537 17156
rect 27571 17184 27583 17187
rect 28169 17187 28227 17193
rect 28169 17184 28181 17187
rect 27571 17156 28181 17184
rect 27571 17153 27583 17156
rect 27525 17147 27583 17153
rect 28169 17153 28181 17156
rect 28215 17184 28227 17187
rect 29270 17184 29276 17196
rect 28215 17156 29276 17184
rect 28215 17153 28227 17156
rect 28169 17147 28227 17153
rect 29270 17144 29276 17156
rect 29328 17144 29334 17196
rect 29638 17184 29644 17196
rect 29564 17156 29644 17184
rect 26237 17119 26295 17125
rect 26237 17116 26249 17119
rect 26200 17088 26249 17116
rect 26200 17076 26206 17088
rect 26237 17085 26249 17088
rect 26283 17085 26295 17119
rect 26510 17116 26516 17128
rect 26471 17088 26516 17116
rect 26237 17079 26295 17085
rect 26510 17076 26516 17088
rect 26568 17076 26574 17128
rect 29564 17125 29592 17156
rect 29638 17144 29644 17156
rect 29696 17144 29702 17196
rect 30282 17184 30288 17196
rect 29748 17156 30288 17184
rect 29748 17127 29776 17156
rect 30282 17144 30288 17156
rect 30340 17184 30346 17196
rect 30926 17184 30932 17196
rect 30340 17156 30932 17184
rect 30340 17144 30346 17156
rect 30926 17144 30932 17156
rect 30984 17144 30990 17196
rect 31036 17193 31064 17292
rect 31021 17187 31079 17193
rect 31021 17153 31033 17187
rect 31067 17153 31079 17187
rect 31021 17147 31079 17153
rect 28445 17119 28503 17125
rect 28445 17085 28457 17119
rect 28491 17116 28503 17119
rect 29549 17119 29607 17125
rect 29549 17116 29561 17119
rect 28491 17088 29561 17116
rect 28491 17085 28503 17088
rect 28445 17079 28503 17085
rect 29549 17085 29561 17088
rect 29595 17085 29607 17119
rect 29549 17079 29607 17085
rect 29733 17121 29791 17127
rect 29733 17087 29745 17121
rect 29779 17087 29791 17121
rect 29733 17081 29791 17087
rect 29822 17076 29828 17128
rect 29880 17116 29886 17128
rect 30006 17125 30012 17128
rect 29963 17119 30012 17125
rect 29880 17088 29925 17116
rect 29880 17076 29886 17088
rect 29963 17085 29975 17119
rect 30009 17085 30012 17119
rect 29963 17079 30012 17085
rect 30006 17076 30012 17079
rect 30064 17076 30070 17128
rect 30098 17076 30104 17128
rect 30156 17116 30162 17128
rect 30466 17116 30472 17128
rect 30156 17088 30472 17116
rect 30156 17076 30162 17088
rect 30466 17076 30472 17088
rect 30524 17076 30530 17128
rect 30650 17076 30656 17128
rect 30708 17116 30714 17128
rect 30745 17119 30803 17125
rect 30745 17116 30757 17119
rect 30708 17088 30757 17116
rect 30708 17076 30714 17088
rect 30745 17085 30757 17088
rect 30791 17085 30803 17119
rect 30745 17079 30803 17085
rect 23256 17020 23704 17048
rect 23845 17051 23903 17057
rect 23256 17008 23262 17020
rect 23845 17017 23857 17051
rect 23891 17048 23903 17051
rect 25510 17051 25568 17057
rect 25510 17048 25522 17051
rect 23891 17020 25522 17048
rect 23891 17017 23903 17020
rect 23845 17011 23903 17017
rect 25510 17017 25522 17020
rect 25556 17017 25568 17051
rect 25510 17011 25568 17017
rect 21910 16980 21916 16992
rect 20364 16952 21916 16980
rect 21910 16940 21916 16952
rect 21968 16940 21974 16992
rect 22186 16980 22192 16992
rect 22147 16952 22192 16980
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 23106 16940 23112 16992
rect 23164 16980 23170 16992
rect 26970 16980 26976 16992
rect 23164 16952 26976 16980
rect 23164 16940 23170 16952
rect 26970 16940 26976 16952
rect 27028 16940 27034 16992
rect 28810 16940 28816 16992
rect 28868 16980 28874 16992
rect 30745 16983 30803 16989
rect 30745 16980 30757 16983
rect 28868 16952 30757 16980
rect 28868 16940 28874 16952
rect 30745 16949 30757 16952
rect 30791 16949 30803 16983
rect 30745 16943 30803 16949
rect 1104 16890 32016 16912
rect 1104 16838 11253 16890
rect 11305 16838 11317 16890
rect 11369 16838 11381 16890
rect 11433 16838 11445 16890
rect 11497 16838 11509 16890
rect 11561 16838 21557 16890
rect 21609 16838 21621 16890
rect 21673 16838 21685 16890
rect 21737 16838 21749 16890
rect 21801 16838 21813 16890
rect 21865 16838 32016 16890
rect 1104 16816 32016 16838
rect 1210 16736 1216 16788
rect 1268 16776 1274 16788
rect 1397 16779 1455 16785
rect 1397 16776 1409 16779
rect 1268 16748 1409 16776
rect 1268 16736 1274 16748
rect 1397 16745 1409 16748
rect 1443 16776 1455 16779
rect 2590 16776 2596 16788
rect 1443 16748 2596 16776
rect 1443 16745 1455 16748
rect 1397 16739 1455 16745
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 3329 16779 3387 16785
rect 3329 16745 3341 16779
rect 3375 16776 3387 16779
rect 3418 16776 3424 16788
rect 3375 16748 3424 16776
rect 3375 16745 3387 16748
rect 3329 16739 3387 16745
rect 3418 16736 3424 16748
rect 3476 16776 3482 16788
rect 3694 16776 3700 16788
rect 3476 16748 3700 16776
rect 3476 16736 3482 16748
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 4154 16776 4160 16788
rect 4067 16748 4160 16776
rect 4154 16736 4160 16748
rect 4212 16776 4218 16788
rect 6457 16779 6515 16785
rect 4212 16748 5580 16776
rect 4212 16736 4218 16748
rect 1394 16600 1400 16652
rect 1452 16640 1458 16652
rect 1946 16640 1952 16652
rect 1452 16612 1952 16640
rect 1452 16600 1458 16612
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2130 16640 2136 16652
rect 2091 16612 2136 16640
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 2222 16600 2228 16652
rect 2280 16640 2286 16652
rect 2501 16643 2559 16649
rect 2280 16612 2325 16640
rect 2280 16600 2286 16612
rect 2501 16609 2513 16643
rect 2547 16609 2559 16643
rect 2501 16603 2559 16609
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2317 16575 2375 16581
rect 2317 16572 2329 16575
rect 2096 16544 2329 16572
rect 2096 16532 2102 16544
rect 2317 16541 2329 16544
rect 2363 16541 2375 16575
rect 2516 16572 2544 16603
rect 3142 16600 3148 16652
rect 3200 16640 3206 16652
rect 4172 16649 4200 16736
rect 5074 16668 5080 16720
rect 5132 16708 5138 16720
rect 5445 16711 5503 16717
rect 5445 16708 5457 16711
rect 5132 16680 5457 16708
rect 5132 16668 5138 16680
rect 5445 16677 5457 16680
rect 5491 16677 5503 16711
rect 5552 16708 5580 16748
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 6730 16776 6736 16788
rect 6503 16748 6736 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 6730 16736 6736 16748
rect 6788 16776 6794 16788
rect 7374 16776 7380 16788
rect 6788 16748 7380 16776
rect 6788 16736 6794 16748
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 9214 16736 9220 16788
rect 9272 16776 9278 16788
rect 9272 16748 9628 16776
rect 9272 16736 9278 16748
rect 5552 16680 9444 16708
rect 5445 16671 5503 16677
rect 9416 16652 9444 16680
rect 4157 16643 4215 16649
rect 3200 16612 3245 16640
rect 3200 16600 3206 16612
rect 4157 16609 4169 16643
rect 4203 16609 4215 16643
rect 4706 16640 4712 16652
rect 4667 16612 4712 16640
rect 4157 16603 4215 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 4798 16600 4804 16652
rect 4856 16640 4862 16652
rect 4856 16612 4901 16640
rect 4856 16600 4862 16612
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 7570 16643 7628 16649
rect 7570 16640 7582 16643
rect 7064 16612 7582 16640
rect 7064 16600 7070 16612
rect 7570 16609 7582 16612
rect 7616 16609 7628 16643
rect 8938 16640 8944 16652
rect 8899 16612 8944 16640
rect 7570 16603 7628 16609
rect 8938 16600 8944 16612
rect 8996 16600 9002 16652
rect 9398 16640 9404 16652
rect 9359 16612 9404 16640
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 4246 16572 4252 16584
rect 2516 16544 4252 16572
rect 2317 16535 2375 16541
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16572 7895 16575
rect 8846 16572 8852 16584
rect 7883 16544 8852 16572
rect 7883 16541 7895 16544
rect 7837 16535 7895 16541
rect 8846 16532 8852 16544
rect 8904 16572 8910 16584
rect 9214 16572 9220 16584
rect 8904 16544 9220 16572
rect 8904 16532 8910 16544
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 9600 16572 9628 16748
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10594 16776 10600 16788
rect 9916 16748 10600 16776
rect 9916 16736 9922 16748
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 10689 16779 10747 16785
rect 10689 16745 10701 16779
rect 10735 16776 10747 16779
rect 11974 16776 11980 16788
rect 10735 16748 11980 16776
rect 10735 16745 10747 16748
rect 10689 16739 10747 16745
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 12342 16776 12348 16788
rect 12176 16748 12348 16776
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 10505 16711 10563 16717
rect 10505 16708 10517 16711
rect 10284 16680 10517 16708
rect 10284 16668 10290 16680
rect 10505 16677 10517 16680
rect 10551 16677 10563 16711
rect 10505 16671 10563 16677
rect 11054 16668 11060 16720
rect 11112 16708 11118 16720
rect 12176 16708 12204 16748
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 13538 16776 13544 16788
rect 12492 16748 13544 16776
rect 12492 16736 12498 16748
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 14001 16779 14059 16785
rect 14001 16745 14013 16779
rect 14047 16776 14059 16779
rect 14366 16776 14372 16788
rect 14047 16748 14372 16776
rect 14047 16745 14059 16748
rect 14001 16739 14059 16745
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 14645 16779 14703 16785
rect 14645 16745 14657 16779
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 11112 16680 12204 16708
rect 11112 16668 11118 16680
rect 13906 16668 13912 16720
rect 13964 16708 13970 16720
rect 14550 16708 14556 16720
rect 13964 16680 14556 16708
rect 13964 16668 13970 16680
rect 14550 16668 14556 16680
rect 14608 16708 14614 16720
rect 14660 16708 14688 16739
rect 15562 16736 15568 16788
rect 15620 16736 15626 16788
rect 15838 16736 15844 16788
rect 15896 16776 15902 16788
rect 17402 16776 17408 16788
rect 15896 16748 17408 16776
rect 15896 16736 15902 16748
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 17586 16736 17592 16788
rect 17644 16776 17650 16788
rect 17862 16776 17868 16788
rect 17644 16748 17868 16776
rect 17644 16736 17650 16748
rect 17862 16736 17868 16748
rect 17920 16776 17926 16788
rect 18049 16779 18107 16785
rect 18049 16776 18061 16779
rect 17920 16748 18061 16776
rect 17920 16736 17926 16748
rect 18049 16745 18061 16748
rect 18095 16745 18107 16779
rect 18049 16739 18107 16745
rect 20254 16736 20260 16788
rect 20312 16776 20318 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 20312 16748 21189 16776
rect 20312 16736 20318 16748
rect 21177 16745 21189 16748
rect 21223 16776 21235 16779
rect 22462 16776 22468 16788
rect 21223 16748 22468 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 22554 16736 22560 16788
rect 22612 16776 22618 16788
rect 22649 16779 22707 16785
rect 22649 16776 22661 16779
rect 22612 16748 22661 16776
rect 22612 16736 22618 16748
rect 22649 16745 22661 16748
rect 22695 16745 22707 16779
rect 23750 16776 23756 16788
rect 23711 16748 23756 16776
rect 22649 16739 22707 16745
rect 23750 16736 23756 16748
rect 23808 16736 23814 16788
rect 26142 16776 26148 16788
rect 24504 16748 26148 16776
rect 15580 16708 15608 16736
rect 18138 16708 18144 16720
rect 14608 16680 14688 16708
rect 15396 16680 15608 16708
rect 16684 16680 18144 16708
rect 14608 16668 14614 16680
rect 11517 16643 11575 16649
rect 10336 16612 11468 16640
rect 10336 16572 10364 16612
rect 9600 16544 10364 16572
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 3973 16507 4031 16513
rect 3973 16504 3985 16507
rect 2648 16476 3985 16504
rect 2648 16464 2654 16476
rect 3973 16473 3985 16476
rect 4019 16473 4031 16507
rect 3973 16467 4031 16473
rect 5629 16507 5687 16513
rect 5629 16473 5641 16507
rect 5675 16504 5687 16507
rect 6546 16504 6552 16516
rect 5675 16476 6552 16504
rect 5675 16473 5687 16476
rect 5629 16467 5687 16473
rect 6546 16464 6552 16476
rect 6604 16464 6610 16516
rect 9600 16513 9628 16544
rect 10410 16532 10416 16584
rect 10468 16572 10474 16584
rect 11440 16572 11468 16612
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 11698 16640 11704 16652
rect 11563 16612 11704 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 11698 16600 11704 16612
rect 11756 16640 11762 16652
rect 11974 16640 11980 16652
rect 11756 16612 11980 16640
rect 11756 16600 11762 16612
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12158 16600 12164 16652
rect 12216 16640 12222 16652
rect 12894 16640 12900 16652
rect 12216 16612 12900 16640
rect 12216 16600 12222 16612
rect 12894 16600 12900 16612
rect 12952 16640 12958 16652
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 12952 16612 13277 16640
rect 12952 16600 12958 16612
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 13446 16640 13452 16652
rect 13407 16612 13452 16640
rect 13265 16603 13323 16609
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16640 13875 16643
rect 13998 16640 14004 16652
rect 13863 16612 14004 16640
rect 13863 16609 13875 16612
rect 13817 16603 13875 16609
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14829 16643 14887 16649
rect 14829 16609 14841 16643
rect 14875 16640 14887 16643
rect 14918 16640 14924 16652
rect 14875 16612 14924 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15396 16649 15424 16680
rect 15381 16643 15439 16649
rect 15381 16640 15393 16643
rect 15252 16612 15393 16640
rect 15252 16600 15258 16612
rect 15381 16609 15393 16612
rect 15427 16609 15439 16643
rect 15562 16640 15568 16652
rect 15523 16612 15568 16640
rect 15381 16603 15439 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 15930 16640 15936 16652
rect 15891 16612 15936 16640
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 16684 16649 16712 16680
rect 18138 16668 18144 16680
rect 18196 16708 18202 16720
rect 20806 16708 20812 16720
rect 18196 16680 20812 16708
rect 18196 16668 18202 16680
rect 16942 16649 16948 16652
rect 16669 16643 16727 16649
rect 16669 16609 16681 16643
rect 16715 16609 16727 16643
rect 16936 16640 16948 16649
rect 16903 16612 16948 16640
rect 16669 16603 16727 16609
rect 16936 16603 16948 16612
rect 16942 16600 16948 16603
rect 17000 16600 17006 16652
rect 17402 16600 17408 16652
rect 17460 16640 17466 16652
rect 17954 16640 17960 16652
rect 17460 16612 17960 16640
rect 17460 16600 17466 16612
rect 17954 16600 17960 16612
rect 18012 16640 18018 16652
rect 18509 16643 18567 16649
rect 18509 16640 18521 16643
rect 18012 16612 18521 16640
rect 18012 16600 18018 16612
rect 18509 16609 18521 16612
rect 18555 16609 18567 16643
rect 18509 16603 18567 16609
rect 18598 16600 18604 16652
rect 18656 16640 18662 16652
rect 18693 16643 18751 16649
rect 18693 16640 18705 16643
rect 18656 16612 18705 16640
rect 18656 16600 18662 16612
rect 18693 16609 18705 16612
rect 18739 16609 18751 16643
rect 18874 16640 18880 16652
rect 18835 16612 18880 16640
rect 18693 16603 18751 16609
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 19058 16640 19064 16652
rect 18971 16612 19064 16640
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 19812 16649 19840 16680
rect 20806 16668 20812 16680
rect 20864 16668 20870 16720
rect 24504 16708 24532 16748
rect 26142 16736 26148 16748
rect 26200 16736 26206 16788
rect 26970 16776 26976 16788
rect 26931 16748 26976 16776
rect 26970 16736 26976 16748
rect 27028 16736 27034 16788
rect 28902 16736 28908 16788
rect 28960 16776 28966 16788
rect 28960 16748 30144 16776
rect 28960 16736 28966 16748
rect 27709 16711 27767 16717
rect 27709 16708 27721 16711
rect 21836 16680 24532 16708
rect 24596 16680 27721 16708
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 19886 16600 19892 16652
rect 19944 16640 19950 16652
rect 20053 16643 20111 16649
rect 20053 16640 20065 16643
rect 19944 16612 20065 16640
rect 19944 16600 19950 16612
rect 20053 16609 20065 16612
rect 20099 16609 20111 16643
rect 20053 16603 20111 16609
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 21836 16640 21864 16680
rect 22002 16640 22008 16652
rect 20588 16612 21864 16640
rect 21963 16612 22008 16640
rect 20588 16600 20594 16612
rect 22002 16600 22008 16612
rect 22060 16600 22066 16652
rect 22186 16640 22192 16652
rect 22147 16612 22192 16640
rect 22186 16600 22192 16612
rect 22244 16600 22250 16652
rect 22830 16640 22836 16652
rect 22791 16612 22836 16640
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 23106 16640 23112 16652
rect 23067 16612 23112 16640
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 23293 16643 23351 16649
rect 23293 16609 23305 16643
rect 23339 16640 23351 16643
rect 23566 16640 23572 16652
rect 23339 16612 23572 16640
rect 23339 16609 23351 16612
rect 23293 16603 23351 16609
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 23842 16600 23848 16652
rect 23900 16640 23906 16652
rect 24596 16649 24624 16680
rect 27709 16677 27721 16680
rect 27755 16708 27767 16711
rect 27755 16680 29224 16708
rect 27755 16677 27767 16680
rect 27709 16671 27767 16677
rect 24581 16643 24639 16649
rect 24581 16640 24593 16643
rect 23900 16612 24593 16640
rect 23900 16600 23906 16612
rect 24581 16609 24593 16612
rect 24627 16609 24639 16643
rect 24581 16603 24639 16609
rect 24670 16600 24676 16652
rect 24728 16640 24734 16652
rect 25593 16643 25651 16649
rect 25593 16640 25605 16643
rect 24728 16612 25605 16640
rect 24728 16600 24734 16612
rect 25593 16609 25605 16612
rect 25639 16609 25651 16643
rect 25866 16640 25872 16652
rect 25827 16612 25872 16640
rect 25593 16603 25651 16609
rect 25866 16600 25872 16612
rect 25924 16640 25930 16652
rect 26142 16640 26148 16652
rect 25924 16612 26148 16640
rect 25924 16600 25930 16612
rect 26142 16600 26148 16612
rect 26200 16600 26206 16652
rect 28442 16600 28448 16652
rect 28500 16640 28506 16652
rect 28721 16643 28779 16649
rect 28721 16640 28733 16643
rect 28500 16612 28733 16640
rect 28500 16600 28506 16612
rect 28721 16609 28733 16612
rect 28767 16609 28779 16643
rect 28902 16640 28908 16652
rect 28815 16612 28908 16640
rect 28721 16603 28779 16609
rect 28902 16600 28908 16612
rect 28960 16600 28966 16652
rect 29196 16640 29224 16680
rect 29270 16668 29276 16720
rect 29328 16708 29334 16720
rect 29454 16708 29460 16720
rect 29328 16680 29460 16708
rect 29328 16668 29334 16680
rect 29454 16668 29460 16680
rect 29512 16668 29518 16720
rect 30116 16708 30144 16748
rect 30190 16736 30196 16788
rect 30248 16776 30254 16788
rect 30285 16779 30343 16785
rect 30285 16776 30297 16779
rect 30248 16748 30297 16776
rect 30248 16736 30254 16748
rect 30285 16745 30297 16748
rect 30331 16745 30343 16779
rect 30285 16739 30343 16745
rect 30558 16736 30564 16788
rect 30616 16776 30622 16788
rect 30834 16776 30840 16788
rect 30616 16748 30840 16776
rect 30616 16736 30622 16748
rect 30834 16736 30840 16748
rect 30892 16736 30898 16788
rect 31018 16736 31024 16788
rect 31076 16776 31082 16788
rect 31113 16779 31171 16785
rect 31113 16776 31125 16779
rect 31076 16748 31125 16776
rect 31076 16736 31082 16748
rect 31113 16745 31125 16748
rect 31159 16745 31171 16779
rect 31113 16739 31171 16745
rect 30466 16708 30472 16720
rect 30116 16680 30472 16708
rect 30466 16668 30472 16680
rect 30524 16668 30530 16720
rect 29549 16643 29607 16649
rect 29196 16612 29316 16640
rect 11790 16572 11796 16584
rect 10468 16544 10824 16572
rect 11440 16544 11652 16572
rect 11751 16544 11796 16572
rect 10468 16532 10474 16544
rect 9585 16507 9643 16513
rect 9585 16473 9597 16507
rect 9631 16473 9643 16507
rect 9585 16467 9643 16473
rect 9950 16464 9956 16516
rect 10008 16504 10014 16516
rect 10137 16507 10195 16513
rect 10137 16504 10149 16507
rect 10008 16476 10149 16504
rect 10008 16464 10014 16476
rect 10137 16473 10149 16476
rect 10183 16504 10195 16507
rect 10686 16504 10692 16516
rect 10183 16476 10692 16504
rect 10183 16473 10195 16476
rect 10137 16467 10195 16473
rect 10686 16464 10692 16476
rect 10744 16464 10750 16516
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 2685 16439 2743 16445
rect 2685 16436 2697 16439
rect 2556 16408 2697 16436
rect 2556 16396 2562 16408
rect 2685 16405 2697 16408
rect 2731 16405 2743 16439
rect 2685 16399 2743 16405
rect 3694 16396 3700 16448
rect 3752 16436 3758 16448
rect 4062 16436 4068 16448
rect 3752 16408 4068 16436
rect 3752 16396 3758 16408
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 8846 16436 8852 16448
rect 8807 16408 8852 16436
rect 8846 16396 8852 16408
rect 8904 16396 8910 16448
rect 10502 16436 10508 16448
rect 10463 16408 10508 16436
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 10796 16436 10824 16544
rect 11624 16504 11652 16544
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 12802 16572 12808 16584
rect 12176 16544 12808 16572
rect 12176 16504 12204 16544
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 13136 16544 13553 16572
rect 13136 16532 13142 16544
rect 13541 16541 13553 16544
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16572 13691 16575
rect 14182 16572 14188 16584
rect 13679 16544 14188 16572
rect 13679 16541 13691 16544
rect 13633 16535 13691 16541
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 15286 16572 15292 16584
rect 14424 16544 15292 16572
rect 14424 16532 14430 16544
rect 15286 16532 15292 16544
rect 15344 16572 15350 16584
rect 15657 16575 15715 16581
rect 15657 16572 15669 16575
rect 15344 16544 15669 16572
rect 15344 16532 15350 16544
rect 15657 16541 15669 16544
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16572 15807 16575
rect 15838 16572 15844 16584
rect 15795 16544 15844 16572
rect 15795 16541 15807 16544
rect 15749 16535 15807 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 18782 16572 18788 16584
rect 18196 16544 18788 16572
rect 18196 16532 18202 16544
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 11624 16476 12204 16504
rect 12259 16476 16427 16504
rect 12259 16436 12287 16476
rect 10796 16408 12287 16436
rect 12802 16396 12808 16448
rect 12860 16436 12866 16448
rect 13262 16436 13268 16448
rect 12860 16408 13268 16436
rect 12860 16396 12866 16408
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 16117 16439 16175 16445
rect 16117 16405 16129 16439
rect 16163 16436 16175 16439
rect 16298 16436 16304 16448
rect 16163 16408 16304 16436
rect 16163 16405 16175 16408
rect 16117 16399 16175 16405
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16399 16436 16427 16476
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 19076 16504 19104 16600
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16572 23075 16575
rect 23198 16572 23204 16584
rect 23063 16544 23204 16572
rect 23063 16541 23075 16544
rect 23017 16535 23075 16541
rect 18288 16476 19104 16504
rect 18288 16464 18294 16476
rect 19150 16464 19156 16516
rect 19208 16504 19214 16516
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 19208 16476 19257 16504
rect 19208 16464 19214 16476
rect 19245 16473 19257 16476
rect 19291 16473 19303 16507
rect 19245 16467 19303 16473
rect 21836 16436 21864 16535
rect 23198 16532 23204 16544
rect 23256 16532 23262 16584
rect 24302 16572 24308 16584
rect 24263 16544 24308 16572
rect 24302 16532 24308 16544
rect 24360 16532 24366 16584
rect 27246 16532 27252 16584
rect 27304 16572 27310 16584
rect 27893 16575 27951 16581
rect 27893 16572 27905 16575
rect 27304 16544 27905 16572
rect 27304 16532 27310 16544
rect 27893 16541 27905 16544
rect 27939 16541 27951 16575
rect 27893 16535 27951 16541
rect 28629 16575 28687 16581
rect 28629 16541 28641 16575
rect 28675 16572 28687 16575
rect 28810 16572 28816 16584
rect 28675 16544 28816 16572
rect 28675 16541 28687 16544
rect 28629 16535 28687 16541
rect 28810 16532 28816 16544
rect 28868 16532 28874 16584
rect 22922 16504 22928 16516
rect 22883 16476 22928 16504
rect 22922 16464 22928 16476
rect 22980 16464 22986 16516
rect 24486 16464 24492 16516
rect 24544 16504 24550 16516
rect 28074 16504 28080 16516
rect 24544 16476 28080 16504
rect 24544 16464 24550 16476
rect 28074 16464 28080 16476
rect 28132 16464 28138 16516
rect 16399 16408 21864 16436
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 27338 16436 27344 16448
rect 22888 16408 27344 16436
rect 22888 16396 22894 16408
rect 27338 16396 27344 16408
rect 27396 16436 27402 16448
rect 28920 16436 28948 16600
rect 29288 16584 29316 16612
rect 29549 16609 29561 16643
rect 29595 16640 29607 16643
rect 29638 16640 29644 16652
rect 29595 16612 29644 16640
rect 29595 16609 29607 16612
rect 29549 16603 29607 16609
rect 29638 16600 29644 16612
rect 29696 16600 29702 16652
rect 29733 16643 29791 16649
rect 29733 16609 29745 16643
rect 29779 16640 29791 16643
rect 30006 16640 30012 16652
rect 29779 16612 30012 16640
rect 29779 16609 29791 16612
rect 29733 16603 29791 16609
rect 30006 16600 30012 16612
rect 30064 16600 30070 16652
rect 30101 16643 30159 16649
rect 30101 16609 30113 16643
rect 30147 16640 30159 16643
rect 30282 16640 30288 16652
rect 30147 16612 30288 16640
rect 30147 16609 30159 16612
rect 30101 16603 30159 16609
rect 30282 16600 30288 16612
rect 30340 16600 30346 16652
rect 31297 16643 31355 16649
rect 31297 16609 31309 16643
rect 31343 16640 31355 16643
rect 31386 16640 31392 16652
rect 31343 16612 31392 16640
rect 31343 16609 31355 16612
rect 31297 16603 31355 16609
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 29086 16572 29092 16584
rect 29047 16544 29092 16572
rect 29086 16532 29092 16544
rect 29144 16532 29150 16584
rect 29270 16532 29276 16584
rect 29328 16572 29334 16584
rect 29822 16572 29828 16584
rect 29328 16544 29828 16572
rect 29328 16532 29334 16544
rect 29822 16532 29828 16544
rect 29880 16532 29886 16584
rect 29917 16575 29975 16581
rect 29917 16541 29929 16575
rect 29963 16541 29975 16575
rect 29917 16535 29975 16541
rect 29178 16464 29184 16516
rect 29236 16504 29242 16516
rect 29932 16504 29960 16535
rect 29236 16476 29960 16504
rect 29236 16464 29242 16476
rect 27396 16408 28948 16436
rect 27396 16396 27402 16408
rect 1104 16346 32016 16368
rect 1104 16294 6102 16346
rect 6154 16294 6166 16346
rect 6218 16294 6230 16346
rect 6282 16294 6294 16346
rect 6346 16294 6358 16346
rect 6410 16294 16405 16346
rect 16457 16294 16469 16346
rect 16521 16294 16533 16346
rect 16585 16294 16597 16346
rect 16649 16294 16661 16346
rect 16713 16294 26709 16346
rect 26761 16294 26773 16346
rect 26825 16294 26837 16346
rect 26889 16294 26901 16346
rect 26953 16294 26965 16346
rect 27017 16294 32016 16346
rect 1104 16272 32016 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 3053 16235 3111 16241
rect 3053 16232 3065 16235
rect 2096 16204 3065 16232
rect 2096 16192 2102 16204
rect 3053 16201 3065 16204
rect 3099 16201 3111 16235
rect 3053 16195 3111 16201
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4341 16235 4399 16241
rect 4341 16232 4353 16235
rect 4304 16204 4353 16232
rect 4304 16192 4310 16204
rect 4341 16201 4353 16204
rect 4387 16201 4399 16235
rect 4341 16195 4399 16201
rect 4890 16192 4896 16244
rect 4948 16232 4954 16244
rect 5166 16232 5172 16244
rect 4948 16204 5172 16232
rect 4948 16192 4954 16204
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 6917 16235 6975 16241
rect 6917 16201 6929 16235
rect 6963 16232 6975 16235
rect 7006 16232 7012 16244
rect 6963 16204 7012 16232
rect 6963 16201 6975 16204
rect 6917 16195 6975 16201
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8754 16232 8760 16244
rect 8352 16204 8760 16232
rect 8352 16192 8358 16204
rect 8754 16192 8760 16204
rect 8812 16192 8818 16244
rect 12066 16232 12072 16244
rect 11164 16204 12072 16232
rect 9306 16164 9312 16176
rect 6380 16136 9312 16164
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2225 16099 2283 16105
rect 2225 16096 2237 16099
rect 2004 16068 2237 16096
rect 2004 16056 2010 16068
rect 2225 16065 2237 16068
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 2590 16096 2596 16108
rect 2547 16068 2596 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 4890 16096 4896 16108
rect 4851 16068 4896 16096
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5442 16096 5448 16108
rect 5123 16068 5448 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 5442 16056 5448 16068
rect 5500 16096 5506 16108
rect 5629 16099 5687 16105
rect 5629 16096 5641 16099
rect 5500 16068 5641 16096
rect 5500 16056 5506 16068
rect 5629 16065 5641 16068
rect 5675 16065 5687 16099
rect 5629 16059 5687 16065
rect 4246 16028 4252 16040
rect 4159 16000 4252 16028
rect 4246 15988 4252 16000
rect 4304 16028 4310 16040
rect 4614 16028 4620 16040
rect 4304 16000 4620 16028
rect 4304 15988 4310 16000
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5258 16028 5264 16040
rect 5215 16000 5264 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 3142 15960 3148 15972
rect 3055 15932 3148 15960
rect 3142 15920 3148 15932
rect 3200 15960 3206 15972
rect 4982 15960 4988 15972
rect 3200 15932 4988 15960
rect 3200 15920 3206 15932
rect 4982 15920 4988 15932
rect 5040 15920 5046 15972
rect 1302 15852 1308 15904
rect 1360 15892 1366 15904
rect 4062 15892 4068 15904
rect 1360 15864 4068 15892
rect 1360 15852 1366 15864
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4893 15895 4951 15901
rect 4893 15861 4905 15895
rect 4939 15892 4951 15895
rect 5534 15892 5540 15904
rect 4939 15864 5540 15892
rect 4939 15861 4951 15864
rect 4893 15855 4951 15861
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 5644 15892 5672 16059
rect 6380 16037 6408 16136
rect 9306 16124 9312 16136
rect 9364 16124 9370 16176
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7248 16068 7941 16096
rect 7248 16056 7254 16068
rect 7929 16065 7941 16068
rect 7975 16096 7987 16099
rect 8202 16096 8208 16108
rect 7975 16068 8208 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 8343 16068 9352 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 15997 6239 16031
rect 6181 15991 6239 15997
rect 6365 16031 6423 16037
rect 6365 15997 6377 16031
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 6196 15960 6224 15991
rect 6454 15988 6460 16040
rect 6512 16028 6518 16040
rect 6730 16028 6736 16040
rect 6512 16000 6557 16028
rect 6691 16000 6736 16028
rect 6512 15988 6518 16000
rect 6730 15988 6736 16000
rect 6788 15988 6794 16040
rect 7650 16028 7656 16040
rect 7611 16000 7656 16028
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 15997 7803 16031
rect 8386 16028 8392 16040
rect 8347 16000 8392 16028
rect 7745 15991 7803 15997
rect 6822 15960 6828 15972
rect 6196 15932 6828 15960
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 7282 15920 7288 15972
rect 7340 15960 7346 15972
rect 7760 15960 7788 15991
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 8846 15988 8852 16040
rect 8904 16028 8910 16040
rect 9324 16037 9352 16068
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 10284 16068 10425 16096
rect 10284 16056 10290 16068
rect 10413 16065 10425 16068
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 9033 16031 9091 16037
rect 9033 16028 9045 16031
rect 8904 16000 9045 16028
rect 8904 15988 8910 16000
rect 9033 15997 9045 16000
rect 9079 15997 9091 16031
rect 9033 15991 9091 15997
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 15997 9367 16031
rect 9674 16028 9680 16040
rect 9635 16000 9680 16028
rect 9309 15991 9367 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10042 16028 10048 16040
rect 10003 16000 10048 16028
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11054 16028 11060 16040
rect 11011 16000 11060 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11164 16037 11192 16204
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 14366 16232 14372 16244
rect 13136 16204 14372 16232
rect 13136 16192 13142 16204
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 15194 16232 15200 16244
rect 14507 16204 15200 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 15528 16204 16436 16232
rect 15528 16192 15534 16204
rect 16408 16176 16436 16204
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 18046 16232 18052 16244
rect 17368 16204 18052 16232
rect 17368 16192 17374 16204
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 19150 16232 19156 16244
rect 18840 16204 19156 16232
rect 18840 16192 18846 16204
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 20806 16192 20812 16244
rect 20864 16232 20870 16244
rect 20901 16235 20959 16241
rect 20901 16232 20913 16235
rect 20864 16204 20913 16232
rect 20864 16192 20870 16204
rect 20901 16201 20913 16204
rect 20947 16201 20959 16235
rect 20901 16195 20959 16201
rect 21450 16192 21456 16244
rect 21508 16232 21514 16244
rect 21821 16235 21879 16241
rect 21821 16232 21833 16235
rect 21508 16204 21833 16232
rect 21508 16192 21514 16204
rect 21821 16201 21833 16204
rect 21867 16201 21879 16235
rect 21821 16195 21879 16201
rect 23474 16192 23480 16244
rect 23532 16232 23538 16244
rect 24670 16232 24676 16244
rect 23532 16204 24676 16232
rect 23532 16192 23538 16204
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 27430 16192 27436 16244
rect 27488 16232 27494 16244
rect 28445 16235 28503 16241
rect 28445 16232 28457 16235
rect 27488 16204 28457 16232
rect 27488 16192 27494 16204
rect 28445 16201 28457 16204
rect 28491 16232 28503 16235
rect 28626 16232 28632 16244
rect 28491 16204 28632 16232
rect 28491 16201 28503 16204
rect 28445 16195 28503 16201
rect 28626 16192 28632 16204
rect 28684 16192 28690 16244
rect 28997 16235 29055 16241
rect 28997 16201 29009 16235
rect 29043 16232 29055 16235
rect 29454 16232 29460 16244
rect 29043 16204 29460 16232
rect 29043 16201 29055 16204
rect 28997 16195 29055 16201
rect 29454 16192 29460 16204
rect 29512 16192 29518 16244
rect 30098 16232 30104 16244
rect 30059 16204 30104 16232
rect 30098 16192 30104 16204
rect 30156 16192 30162 16244
rect 11330 16124 11336 16176
rect 11388 16164 11394 16176
rect 11388 16136 12204 16164
rect 11388 16124 11394 16136
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16096 11299 16099
rect 11790 16096 11796 16108
rect 11287 16068 11796 16096
rect 11287 16065 11299 16068
rect 11241 16059 11299 16065
rect 11790 16056 11796 16068
rect 11848 16056 11854 16108
rect 12176 16096 12204 16136
rect 16390 16124 16396 16176
rect 16448 16124 16454 16176
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 16816 16136 22876 16164
rect 16816 16124 16822 16136
rect 15841 16099 15899 16105
rect 12176 16068 12296 16096
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11333 16031 11391 16037
rect 11333 15997 11345 16031
rect 11379 16028 11391 16031
rect 11422 16028 11428 16040
rect 11379 16000 11428 16028
rect 11379 15997 11391 16000
rect 11333 15991 11391 15997
rect 11422 15988 11428 16000
rect 11480 15988 11486 16040
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 7340 15932 7788 15960
rect 7340 15920 7346 15932
rect 7558 15892 7564 15904
rect 5644 15864 7564 15892
rect 7558 15852 7564 15864
rect 7616 15852 7622 15904
rect 11532 15892 11560 15991
rect 12066 15988 12072 16040
rect 12124 16028 12130 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 12124 16000 12173 16028
rect 12124 15988 12130 16000
rect 12161 15997 12173 16000
rect 12207 15997 12219 16031
rect 12268 16028 12296 16068
rect 15841 16065 15853 16099
rect 15887 16096 15899 16099
rect 16114 16096 16120 16108
rect 15887 16068 16120 16096
rect 15887 16065 15899 16068
rect 15841 16059 15899 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16298 16096 16304 16108
rect 16259 16068 16304 16096
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 17310 16096 17316 16108
rect 16908 16068 17316 16096
rect 16908 16056 16914 16068
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16096 17831 16099
rect 18138 16096 18144 16108
rect 17819 16068 18144 16096
rect 17819 16065 17831 16068
rect 17773 16059 17831 16065
rect 18138 16056 18144 16068
rect 18196 16056 18202 16108
rect 18322 16056 18328 16108
rect 18380 16096 18386 16108
rect 18874 16096 18880 16108
rect 18380 16068 18880 16096
rect 18380 16056 18386 16068
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19886 16096 19892 16108
rect 19392 16068 19892 16096
rect 19392 16056 19398 16068
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 12268 16000 13860 16028
rect 12161 15991 12219 15997
rect 11701 15963 11759 15969
rect 11701 15929 11713 15963
rect 11747 15960 11759 15963
rect 12406 15963 12464 15969
rect 12406 15960 12418 15963
rect 11747 15932 12418 15960
rect 11747 15929 11759 15932
rect 11701 15923 11759 15929
rect 12406 15929 12418 15932
rect 12452 15929 12464 15963
rect 12406 15923 12464 15929
rect 12618 15920 12624 15972
rect 12676 15960 12682 15972
rect 13262 15960 13268 15972
rect 12676 15932 13268 15960
rect 12676 15920 12682 15932
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 13832 15960 13860 16000
rect 13906 15988 13912 16040
rect 13964 16028 13970 16040
rect 14826 16028 14832 16040
rect 13964 16000 14832 16028
rect 13964 15988 13970 16000
rect 14826 15988 14832 16000
rect 14884 16028 14890 16040
rect 14884 16000 15792 16028
rect 14884 15988 14890 16000
rect 14918 15960 14924 15972
rect 13832 15932 14924 15960
rect 14918 15920 14924 15932
rect 14976 15920 14982 15972
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 15574 15963 15632 15969
rect 15574 15960 15586 15963
rect 15436 15932 15586 15960
rect 15436 15920 15442 15932
rect 15574 15929 15586 15932
rect 15620 15929 15632 15963
rect 15764 15960 15792 16000
rect 16206 15988 16212 16040
rect 16264 16028 16270 16040
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 16264 16000 16497 16028
rect 16264 15988 16270 16000
rect 16485 15997 16497 16000
rect 16531 15997 16543 16031
rect 16485 15991 16543 15997
rect 16761 16031 16819 16037
rect 16761 15997 16773 16031
rect 16807 16028 16819 16031
rect 16942 16028 16948 16040
rect 16807 16000 16948 16028
rect 16807 15997 16819 16000
rect 16761 15991 16819 15997
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 17402 15988 17408 16040
rect 17460 16028 17466 16040
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17460 16000 17509 16028
rect 17460 15988 17466 16000
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 17681 16031 17739 16037
rect 17681 16028 17693 16031
rect 17644 16000 17693 16028
rect 17644 15988 17650 16000
rect 17681 15997 17693 16000
rect 17727 15997 17739 16031
rect 17681 15991 17739 15997
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 17920 16000 17965 16028
rect 17920 15988 17926 16000
rect 18046 15988 18052 16040
rect 18104 16028 18110 16040
rect 18598 16028 18604 16040
rect 18104 16000 18604 16028
rect 18104 15988 18110 16000
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 19613 16031 19671 16037
rect 19613 15997 19625 16031
rect 19659 16028 19671 16031
rect 20162 16028 20168 16040
rect 19659 16000 20168 16028
rect 19659 15997 19671 16000
rect 19613 15991 19671 15997
rect 16666 15960 16672 15972
rect 15764 15932 16672 15960
rect 15574 15923 15632 15929
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 16850 15960 16856 15972
rect 16811 15932 16856 15960
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 19628 15960 19656 15991
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 22005 16031 22063 16037
rect 22005 15997 22017 16031
rect 22051 16028 22063 16031
rect 22094 16028 22100 16040
rect 22051 16000 22100 16028
rect 22051 15997 22063 16000
rect 22005 15991 22063 15997
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 16951 15932 19656 15960
rect 12894 15892 12900 15904
rect 11532 15864 12900 15892
rect 12894 15852 12900 15864
rect 12952 15892 12958 15904
rect 13354 15892 13360 15904
rect 12952 15864 13360 15892
rect 12952 15852 12958 15864
rect 13354 15852 13360 15864
rect 13412 15892 13418 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 13412 15864 13553 15892
rect 13412 15852 13418 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 16206 15892 16212 15904
rect 15160 15864 16212 15892
rect 15160 15852 15166 15864
rect 16206 15852 16212 15864
rect 16264 15892 16270 15904
rect 16951 15892 16979 15932
rect 16264 15864 16979 15892
rect 16264 15852 16270 15864
rect 18046 15852 18052 15904
rect 18104 15892 18110 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 18104 15864 18245 15892
rect 18104 15852 18110 15864
rect 18233 15861 18245 15864
rect 18279 15861 18291 15895
rect 22462 15892 22468 15904
rect 22423 15864 22468 15892
rect 18233 15855 18291 15861
rect 22462 15852 22468 15864
rect 22520 15852 22526 15904
rect 22848 15892 22876 16136
rect 25222 16096 25228 16108
rect 23860 16068 25228 16096
rect 23860 16037 23888 16068
rect 25222 16056 25228 16068
rect 25280 16056 25286 16108
rect 30006 16056 30012 16108
rect 30064 16096 30070 16108
rect 30064 16068 30696 16096
rect 30064 16056 30070 16068
rect 23845 16031 23903 16037
rect 23845 16028 23857 16031
rect 23492 16000 23857 16028
rect 23492 15972 23520 16000
rect 23845 15997 23857 16000
rect 23891 15997 23903 16031
rect 23845 15991 23903 15997
rect 24302 15988 24308 16040
rect 24360 16028 24366 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24360 16000 24593 16028
rect 24360 15988 24366 16000
rect 24581 15997 24593 16000
rect 24627 15997 24639 16031
rect 24581 15991 24639 15997
rect 26050 15988 26056 16040
rect 26108 16028 26114 16040
rect 30668 16037 30696 16068
rect 27065 16031 27123 16037
rect 27065 16028 27077 16031
rect 26108 16000 27077 16028
rect 26108 15988 26114 16000
rect 27065 15997 27077 16000
rect 27111 15997 27123 16031
rect 27065 15991 27123 15997
rect 30653 16031 30711 16037
rect 30653 15997 30665 16031
rect 30699 15997 30711 16031
rect 30653 15991 30711 15997
rect 23474 15920 23480 15972
rect 23532 15920 23538 15972
rect 23600 15963 23658 15969
rect 23600 15929 23612 15963
rect 23646 15960 23658 15963
rect 23750 15960 23756 15972
rect 23646 15932 23756 15960
rect 23646 15929 23658 15932
rect 23600 15923 23658 15929
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 25492 15963 25550 15969
rect 25492 15929 25504 15963
rect 25538 15960 25550 15963
rect 25774 15960 25780 15972
rect 25538 15932 25780 15960
rect 25538 15929 25550 15932
rect 25492 15923 25550 15929
rect 25774 15920 25780 15932
rect 25832 15920 25838 15972
rect 27332 15963 27390 15969
rect 25884 15932 26740 15960
rect 25884 15892 25912 15932
rect 26602 15892 26608 15904
rect 22848 15864 25912 15892
rect 26563 15864 26608 15892
rect 26602 15852 26608 15864
rect 26660 15852 26666 15904
rect 26712 15892 26740 15932
rect 27332 15929 27344 15963
rect 27378 15960 27390 15963
rect 27706 15960 27712 15972
rect 27378 15932 27712 15960
rect 27378 15929 27390 15932
rect 27332 15923 27390 15929
rect 27706 15920 27712 15932
rect 27764 15920 27770 15972
rect 29178 15920 29184 15972
rect 29236 15960 29242 15972
rect 30009 15963 30067 15969
rect 30009 15960 30021 15963
rect 29236 15932 30021 15960
rect 29236 15920 29242 15932
rect 30009 15929 30021 15932
rect 30055 15929 30067 15963
rect 30009 15923 30067 15929
rect 27522 15892 27528 15904
rect 26712 15864 27528 15892
rect 27522 15852 27528 15864
rect 27580 15852 27586 15904
rect 30745 15895 30803 15901
rect 30745 15861 30757 15895
rect 30791 15892 30803 15895
rect 30926 15892 30932 15904
rect 30791 15864 30932 15892
rect 30791 15861 30803 15864
rect 30745 15855 30803 15861
rect 30926 15852 30932 15864
rect 30984 15852 30990 15904
rect 1104 15802 32016 15824
rect 1104 15750 11253 15802
rect 11305 15750 11317 15802
rect 11369 15750 11381 15802
rect 11433 15750 11445 15802
rect 11497 15750 11509 15802
rect 11561 15750 21557 15802
rect 21609 15750 21621 15802
rect 21673 15750 21685 15802
rect 21737 15750 21749 15802
rect 21801 15750 21813 15802
rect 21865 15750 32016 15802
rect 1104 15728 32016 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 2958 15688 2964 15700
rect 1627 15660 2964 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 4801 15691 4859 15697
rect 4801 15688 4813 15691
rect 4764 15660 4813 15688
rect 4764 15648 4770 15660
rect 4801 15657 4813 15660
rect 4847 15657 4859 15691
rect 4801 15651 4859 15657
rect 7009 15691 7067 15697
rect 7009 15657 7021 15691
rect 7055 15688 7067 15691
rect 8386 15688 8392 15700
rect 7055 15660 8392 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 8849 15691 8907 15697
rect 8849 15657 8861 15691
rect 8895 15688 8907 15691
rect 9674 15688 9680 15700
rect 8895 15660 9680 15688
rect 8895 15657 8907 15660
rect 8849 15651 8907 15657
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10686 15688 10692 15700
rect 10647 15660 10692 15688
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 15378 15688 15384 15700
rect 10796 15660 15240 15688
rect 15339 15660 15384 15688
rect 2682 15620 2688 15632
rect 2240 15592 2688 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1486 15552 1492 15564
rect 1443 15524 1492 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1486 15512 1492 15524
rect 1544 15512 1550 15564
rect 2240 15561 2268 15592
rect 2682 15580 2688 15592
rect 2740 15580 2746 15632
rect 3694 15580 3700 15632
rect 3752 15620 3758 15632
rect 6181 15623 6239 15629
rect 6181 15620 6193 15623
rect 3752 15592 6193 15620
rect 3752 15580 3758 15592
rect 6181 15589 6193 15592
rect 6227 15589 6239 15623
rect 6181 15583 6239 15589
rect 6641 15623 6699 15629
rect 6641 15589 6653 15623
rect 6687 15589 6699 15623
rect 6641 15583 6699 15589
rect 6857 15623 6915 15629
rect 6857 15589 6869 15623
rect 6903 15620 6915 15623
rect 8478 15620 8484 15632
rect 6903 15592 8484 15620
rect 6903 15589 6915 15592
rect 6857 15583 6915 15589
rect 2498 15561 2504 15564
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15521 2283 15555
rect 2492 15552 2504 15561
rect 2459 15524 2504 15552
rect 2225 15515 2283 15521
rect 2492 15515 2504 15524
rect 2498 15512 2504 15515
rect 2556 15512 2562 15564
rect 3786 15512 3792 15564
rect 3844 15552 3850 15564
rect 4433 15555 4491 15561
rect 4433 15552 4445 15555
rect 3844 15524 4445 15552
rect 3844 15512 3850 15524
rect 4433 15521 4445 15524
rect 4479 15521 4491 15555
rect 5258 15552 5264 15564
rect 5219 15524 5264 15552
rect 4433 15515 4491 15521
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 6656 15552 6684 15583
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 9582 15629 9588 15632
rect 9576 15620 9588 15629
rect 9543 15592 9588 15620
rect 9576 15583 9588 15592
rect 9582 15580 9588 15583
rect 9640 15580 9646 15632
rect 7374 15552 7380 15564
rect 6656 15524 7380 15552
rect 7374 15512 7380 15524
rect 7432 15552 7438 15564
rect 7745 15555 7803 15561
rect 7745 15552 7757 15555
rect 7432 15524 7757 15552
rect 7432 15512 7438 15524
rect 7745 15521 7757 15524
rect 7791 15521 7803 15555
rect 7745 15515 7803 15521
rect 7837 15555 7895 15561
rect 7837 15521 7849 15555
rect 7883 15521 7895 15555
rect 7837 15515 7895 15521
rect 4246 15484 4252 15496
rect 3620 15456 4252 15484
rect 3620 15425 3648 15456
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15484 4399 15487
rect 4982 15484 4988 15496
rect 4387 15456 4988 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15484 5595 15487
rect 5626 15484 5632 15496
rect 5583 15456 5632 15484
rect 5583 15453 5595 15456
rect 5537 15447 5595 15453
rect 5626 15444 5632 15456
rect 5684 15444 5690 15496
rect 7558 15444 7564 15496
rect 7616 15484 7622 15496
rect 7852 15484 7880 15515
rect 7926 15512 7932 15564
rect 7984 15552 7990 15564
rect 7984 15524 8029 15552
rect 7984 15512 7990 15524
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 8573 15555 8631 15561
rect 8168 15524 8213 15552
rect 8168 15512 8174 15524
rect 8573 15521 8585 15555
rect 8619 15552 8631 15555
rect 10796 15552 10824 15660
rect 11784 15623 11842 15629
rect 11784 15589 11796 15623
rect 11830 15620 11842 15623
rect 11882 15620 11888 15632
rect 11830 15592 11888 15620
rect 11830 15589 11842 15592
rect 11784 15583 11842 15589
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 13262 15580 13268 15632
rect 13320 15620 13326 15632
rect 13725 15623 13783 15629
rect 13725 15620 13737 15623
rect 13320 15592 13737 15620
rect 13320 15580 13326 15592
rect 13725 15589 13737 15592
rect 13771 15620 13783 15623
rect 14090 15620 14096 15632
rect 13771 15592 14096 15620
rect 13771 15589 13783 15592
rect 13725 15583 13783 15589
rect 14090 15580 14096 15592
rect 14148 15580 14154 15632
rect 15102 15620 15108 15632
rect 14936 15592 15108 15620
rect 8619 15524 8708 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 7616 15456 7880 15484
rect 7616 15444 7622 15456
rect 3605 15419 3663 15425
rect 3605 15385 3617 15419
rect 3651 15385 3663 15419
rect 3605 15379 3663 15385
rect 3878 15376 3884 15428
rect 3936 15416 3942 15428
rect 7852 15416 7880 15456
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8680 15484 8708 15524
rect 8956 15524 10824 15552
rect 11517 15555 11575 15561
rect 8846 15484 8852 15496
rect 8352 15456 8708 15484
rect 8807 15456 8852 15484
rect 8352 15444 8358 15456
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 8956 15416 8984 15524
rect 11517 15521 11529 15555
rect 11563 15552 11575 15555
rect 12066 15552 12072 15564
rect 11563 15524 12072 15552
rect 11563 15521 11575 15524
rect 11517 15515 11575 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 13354 15552 13360 15564
rect 13315 15524 13360 15552
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 14642 15552 14648 15564
rect 14603 15524 14648 15552
rect 14642 15512 14648 15524
rect 14700 15512 14706 15564
rect 14936 15561 14964 15592
rect 15102 15580 15108 15592
rect 15160 15580 15166 15632
rect 15212 15620 15240 15660
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 15562 15648 15568 15700
rect 15620 15688 15626 15700
rect 15933 15691 15991 15697
rect 15933 15688 15945 15691
rect 15620 15660 15945 15688
rect 15620 15648 15626 15660
rect 15933 15657 15945 15660
rect 15979 15657 15991 15691
rect 15933 15651 15991 15657
rect 16390 15648 16396 15700
rect 16448 15688 16454 15700
rect 16448 15660 20300 15688
rect 16448 15648 16454 15660
rect 15212 15592 20208 15620
rect 14829 15555 14887 15561
rect 14829 15521 14841 15555
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 14921 15555 14979 15561
rect 14921 15521 14933 15555
rect 14967 15521 14979 15555
rect 15194 15552 15200 15564
rect 15155 15524 15200 15552
rect 14921 15515 14979 15521
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 9272 15456 9321 15484
rect 9272 15444 9278 15456
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 3936 15388 7788 15416
rect 7852 15388 8984 15416
rect 3936 15376 3942 15388
rect 0 15348 800 15362
rect 1486 15348 1492 15360
rect 0 15320 1492 15348
rect 0 15306 800 15320
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 4706 15348 4712 15360
rect 4396 15320 4712 15348
rect 4396 15308 4402 15320
rect 4706 15308 4712 15320
rect 4764 15348 4770 15360
rect 5353 15351 5411 15357
rect 5353 15348 5365 15351
rect 4764 15320 5365 15348
rect 4764 15308 4770 15320
rect 5353 15317 5365 15320
rect 5399 15317 5411 15351
rect 5353 15311 5411 15317
rect 5445 15351 5503 15357
rect 5445 15317 5457 15351
rect 5491 15348 5503 15351
rect 5810 15348 5816 15360
rect 5491 15320 5816 15348
rect 5491 15317 5503 15320
rect 5445 15311 5503 15317
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 6181 15351 6239 15357
rect 6181 15317 6193 15351
rect 6227 15348 6239 15351
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6227 15320 6837 15348
rect 6227 15317 6239 15320
rect 6181 15311 6239 15317
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 7282 15308 7288 15360
rect 7340 15348 7346 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 7340 15320 7481 15348
rect 7340 15308 7346 15320
rect 7469 15317 7481 15320
rect 7515 15317 7527 15351
rect 7760 15348 7788 15388
rect 8665 15351 8723 15357
rect 8665 15348 8677 15351
rect 7760 15320 8677 15348
rect 7469 15311 7527 15317
rect 8665 15317 8677 15320
rect 8711 15317 8723 15351
rect 9324 15348 9352 15447
rect 13909 15419 13967 15425
rect 13909 15385 13921 15419
rect 13955 15416 13967 15419
rect 14734 15416 14740 15428
rect 13955 15388 14740 15416
rect 13955 15385 13967 15388
rect 13909 15379 13967 15385
rect 14734 15376 14740 15388
rect 14792 15376 14798 15428
rect 14844 15416 14872 15515
rect 15194 15512 15200 15524
rect 15252 15512 15258 15564
rect 15841 15555 15899 15561
rect 15841 15521 15853 15555
rect 15887 15552 15899 15555
rect 15930 15552 15936 15564
rect 15887 15524 15936 15552
rect 15887 15521 15899 15524
rect 15841 15515 15899 15521
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15484 15071 15487
rect 15286 15484 15292 15496
rect 15059 15456 15292 15484
rect 15059 15453 15071 15456
rect 15013 15447 15071 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 15470 15416 15476 15428
rect 14844 15388 15476 15416
rect 15470 15376 15476 15388
rect 15528 15416 15534 15428
rect 15856 15416 15884 15515
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 16761 15555 16819 15561
rect 16761 15552 16773 15555
rect 16724 15524 16773 15552
rect 16724 15512 16730 15524
rect 16761 15521 16773 15524
rect 16807 15521 16819 15555
rect 16761 15515 16819 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15552 17555 15555
rect 17954 15552 17960 15564
rect 17543 15524 17960 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 18138 15552 18144 15564
rect 18099 15524 18144 15552
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 18288 15524 18705 15552
rect 18288 15512 18294 15524
rect 18693 15521 18705 15524
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15521 18935 15555
rect 18877 15515 18935 15521
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 18892 15484 18920 15515
rect 18966 15512 18972 15564
rect 19024 15552 19030 15564
rect 19242 15552 19248 15564
rect 19024 15524 19069 15552
rect 19203 15524 19248 15552
rect 19024 15512 19030 15524
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 19518 15552 19524 15564
rect 19475 15524 19524 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 19058 15484 19064 15496
rect 17451 15456 18920 15484
rect 19019 15456 19064 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 19058 15444 19064 15456
rect 19116 15484 19122 15496
rect 19794 15484 19800 15496
rect 19116 15456 19800 15484
rect 19116 15444 19122 15456
rect 19794 15444 19800 15456
rect 19852 15444 19858 15496
rect 20180 15484 20208 15592
rect 20272 15561 20300 15660
rect 22094 15648 22100 15700
rect 22152 15688 22158 15700
rect 23566 15688 23572 15700
rect 22152 15660 22197 15688
rect 23527 15660 23572 15688
rect 22152 15648 22158 15660
rect 23566 15648 23572 15660
rect 23624 15648 23630 15700
rect 24946 15648 24952 15700
rect 25004 15688 25010 15700
rect 25777 15691 25835 15697
rect 25777 15688 25789 15691
rect 25004 15660 25789 15688
rect 25004 15648 25010 15660
rect 25777 15657 25789 15660
rect 25823 15657 25835 15691
rect 27706 15688 27712 15700
rect 27667 15660 27712 15688
rect 25777 15651 25835 15657
rect 27706 15648 27712 15660
rect 27764 15648 27770 15700
rect 30558 15648 30564 15700
rect 30616 15688 30622 15700
rect 31018 15688 31024 15700
rect 31076 15697 31082 15700
rect 31076 15691 31095 15697
rect 30616 15660 31024 15688
rect 30616 15648 30622 15660
rect 31018 15648 31024 15660
rect 31083 15657 31095 15691
rect 31076 15651 31095 15657
rect 31076 15648 31082 15651
rect 22278 15629 22284 15632
rect 22265 15623 22284 15629
rect 22265 15589 22277 15623
rect 22265 15583 22284 15589
rect 22278 15580 22284 15583
rect 22336 15580 22342 15632
rect 22370 15580 22376 15632
rect 22428 15620 22434 15632
rect 22465 15623 22523 15629
rect 22465 15620 22477 15623
rect 22428 15592 22477 15620
rect 22428 15580 22434 15592
rect 22465 15589 22477 15592
rect 22511 15589 22523 15623
rect 26329 15623 26387 15629
rect 26329 15620 26341 15623
rect 22465 15583 22523 15589
rect 22563 15592 26341 15620
rect 20257 15555 20315 15561
rect 20257 15521 20269 15555
rect 20303 15521 20315 15555
rect 20622 15552 20628 15564
rect 20583 15524 20628 15552
rect 20257 15515 20315 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 21174 15552 21180 15564
rect 21135 15524 21180 15552
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 22563 15552 22591 15592
rect 26329 15589 26341 15592
rect 26375 15589 26387 15623
rect 28166 15620 28172 15632
rect 26329 15583 26387 15589
rect 27356 15592 28172 15620
rect 23106 15552 23112 15564
rect 21284 15524 22591 15552
rect 22756 15524 23112 15552
rect 21284 15484 21312 15524
rect 20180 15456 21312 15484
rect 22462 15444 22468 15496
rect 22520 15484 22526 15496
rect 22756 15484 22784 15524
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 23201 15555 23259 15561
rect 23201 15521 23213 15555
rect 23247 15521 23259 15555
rect 23201 15515 23259 15521
rect 23385 15555 23443 15561
rect 23385 15521 23397 15555
rect 23431 15552 23443 15555
rect 23934 15552 23940 15564
rect 23431 15524 23940 15552
rect 23431 15521 23443 15524
rect 23385 15515 23443 15521
rect 22520 15456 22784 15484
rect 23216 15484 23244 15515
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 24302 15512 24308 15564
rect 24360 15552 24366 15564
rect 24489 15555 24547 15561
rect 24489 15552 24501 15555
rect 24360 15524 24501 15552
rect 24360 15512 24366 15524
rect 24489 15521 24501 15524
rect 24535 15521 24547 15555
rect 24489 15515 24547 15521
rect 26510 15512 26516 15564
rect 26568 15552 26574 15564
rect 27356 15561 27384 15592
rect 28166 15580 28172 15592
rect 28224 15580 28230 15632
rect 30837 15623 30895 15629
rect 30837 15589 30849 15623
rect 30883 15620 30895 15623
rect 30926 15620 30932 15632
rect 30883 15592 30932 15620
rect 30883 15589 30895 15592
rect 30837 15583 30895 15589
rect 30926 15580 30932 15592
rect 30984 15580 30990 15632
rect 26973 15555 27031 15561
rect 26973 15552 26985 15555
rect 26568 15524 26985 15552
rect 26568 15512 26574 15524
rect 26973 15521 26985 15524
rect 27019 15521 27031 15555
rect 27157 15555 27215 15561
rect 27157 15552 27169 15555
rect 26973 15515 27031 15521
rect 27080 15524 27169 15552
rect 23658 15484 23664 15496
rect 23216 15456 23664 15484
rect 22520 15444 22526 15456
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 24762 15484 24768 15496
rect 24723 15456 24768 15484
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 26602 15444 26608 15496
rect 26660 15484 26666 15496
rect 27080 15484 27108 15524
rect 27157 15521 27169 15524
rect 27203 15521 27215 15555
rect 27157 15515 27215 15521
rect 27341 15555 27399 15561
rect 27341 15521 27353 15555
rect 27387 15521 27399 15555
rect 27341 15515 27399 15521
rect 27430 15512 27436 15564
rect 27488 15552 27494 15564
rect 27525 15555 27583 15561
rect 27525 15552 27537 15555
rect 27488 15524 27537 15552
rect 27488 15512 27494 15524
rect 27525 15521 27537 15524
rect 27571 15521 27583 15555
rect 28353 15555 28411 15561
rect 28353 15552 28365 15555
rect 27525 15515 27583 15521
rect 27632 15524 28365 15552
rect 27246 15484 27252 15496
rect 26660 15456 27108 15484
rect 27207 15456 27252 15484
rect 26660 15444 26666 15456
rect 27246 15444 27252 15456
rect 27304 15444 27310 15496
rect 17586 15416 17592 15428
rect 15528 15388 15884 15416
rect 15948 15388 17592 15416
rect 15528 15376 15534 15388
rect 9582 15348 9588 15360
rect 9324 15320 9588 15348
rect 8665 15311 8723 15317
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 12158 15308 12164 15360
rect 12216 15348 12222 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 12216 15320 12909 15348
rect 12216 15308 12222 15320
rect 12897 15317 12909 15320
rect 12943 15348 12955 15351
rect 13538 15348 13544 15360
rect 12943 15320 13544 15348
rect 12943 15317 12955 15320
rect 12897 15311 12955 15317
rect 13538 15308 13544 15320
rect 13596 15348 13602 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13596 15320 13737 15348
rect 13596 15308 13602 15320
rect 13725 15317 13737 15320
rect 13771 15348 13783 15351
rect 13998 15348 14004 15360
rect 13771 15320 14004 15348
rect 13771 15317 13783 15320
rect 13725 15311 13783 15317
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 15378 15348 15384 15360
rect 15160 15320 15384 15348
rect 15160 15308 15166 15320
rect 15378 15308 15384 15320
rect 15436 15348 15442 15360
rect 15948 15348 15976 15388
rect 17586 15376 17592 15388
rect 17644 15416 17650 15428
rect 17957 15419 18015 15425
rect 17957 15416 17969 15419
rect 17644 15388 17969 15416
rect 17644 15376 17650 15388
rect 17957 15385 17969 15388
rect 18003 15416 18015 15419
rect 18966 15416 18972 15428
rect 18003 15388 18972 15416
rect 18003 15385 18015 15388
rect 17957 15379 18015 15385
rect 18966 15376 18972 15388
rect 19024 15376 19030 15428
rect 20254 15416 20260 15428
rect 20215 15388 20260 15416
rect 20254 15376 20260 15388
rect 20312 15376 20318 15428
rect 24670 15376 24676 15428
rect 24728 15416 24734 15428
rect 27632 15416 27660 15524
rect 28353 15521 28365 15524
rect 28399 15552 28411 15555
rect 29178 15552 29184 15564
rect 28399 15524 29184 15552
rect 28399 15521 28411 15524
rect 28353 15515 28411 15521
rect 29178 15512 29184 15524
rect 29236 15512 29242 15564
rect 29270 15512 29276 15564
rect 29328 15552 29334 15564
rect 29328 15524 29373 15552
rect 29328 15512 29334 15524
rect 29546 15484 29552 15496
rect 29507 15456 29552 15484
rect 29546 15444 29552 15456
rect 29604 15444 29610 15496
rect 24728 15388 27660 15416
rect 24728 15376 24734 15388
rect 28350 15376 28356 15428
rect 28408 15416 28414 15428
rect 28408 15388 31754 15416
rect 28408 15376 28414 15388
rect 15436 15320 15976 15348
rect 15436 15308 15442 15320
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 19978 15348 19984 15360
rect 16908 15320 19984 15348
rect 16908 15308 16914 15320
rect 19978 15308 19984 15320
rect 20036 15348 20042 15360
rect 20530 15348 20536 15360
rect 20036 15320 20536 15348
rect 20036 15308 20042 15320
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 22281 15351 22339 15357
rect 22281 15317 22293 15351
rect 22327 15348 22339 15351
rect 22462 15348 22468 15360
rect 22327 15320 22468 15348
rect 22327 15317 22339 15320
rect 22281 15311 22339 15317
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 23934 15308 23940 15360
rect 23992 15348 23998 15360
rect 24854 15348 24860 15360
rect 23992 15320 24860 15348
rect 23992 15308 23998 15320
rect 24854 15308 24860 15320
rect 24912 15308 24918 15360
rect 30834 15308 30840 15360
rect 30892 15348 30898 15360
rect 31021 15351 31079 15357
rect 31021 15348 31033 15351
rect 30892 15320 31033 15348
rect 30892 15308 30898 15320
rect 31021 15317 31033 15320
rect 31067 15317 31079 15351
rect 31202 15348 31208 15360
rect 31163 15320 31208 15348
rect 31021 15311 31079 15317
rect 31202 15308 31208 15320
rect 31260 15308 31266 15360
rect 31726 15348 31754 15388
rect 32320 15348 33120 15362
rect 31726 15320 33120 15348
rect 32320 15306 33120 15320
rect 1104 15258 32016 15280
rect 1104 15206 6102 15258
rect 6154 15206 6166 15258
rect 6218 15206 6230 15258
rect 6282 15206 6294 15258
rect 6346 15206 6358 15258
rect 6410 15206 16405 15258
rect 16457 15206 16469 15258
rect 16521 15206 16533 15258
rect 16585 15206 16597 15258
rect 16649 15206 16661 15258
rect 16713 15206 26709 15258
rect 26761 15206 26773 15258
rect 26825 15206 26837 15258
rect 26889 15206 26901 15258
rect 26953 15206 26965 15258
rect 27017 15206 32016 15258
rect 1104 15184 32016 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 1670 15144 1676 15156
rect 1627 15116 1676 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 1670 15104 1676 15116
rect 1728 15144 1734 15156
rect 4065 15147 4123 15153
rect 4065 15144 4077 15147
rect 1728 15116 4077 15144
rect 1728 15104 1734 15116
rect 4065 15113 4077 15116
rect 4111 15144 4123 15147
rect 4522 15144 4528 15156
rect 4111 15116 4528 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 4706 15104 4712 15156
rect 4764 15144 4770 15156
rect 7834 15144 7840 15156
rect 4764 15116 6684 15144
rect 4764 15104 4770 15116
rect 5994 15076 6000 15088
rect 2884 15048 6000 15076
rect 2884 15017 2912 15048
rect 5994 15036 6000 15048
rect 6052 15036 6058 15088
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 5534 15008 5540 15020
rect 5495 14980 5540 15008
rect 2869 14971 2927 14977
rect 5534 14968 5540 14980
rect 5592 14968 5598 15020
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6656 15008 6684 15116
rect 7116 15116 7840 15144
rect 6730 15036 6736 15088
rect 6788 15076 6794 15088
rect 7116 15085 7144 15116
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 8389 15147 8447 15153
rect 8389 15113 8401 15147
rect 8435 15144 8447 15147
rect 8846 15144 8852 15156
rect 8435 15116 8852 15144
rect 8435 15113 8447 15116
rect 8389 15107 8447 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9677 15147 9735 15153
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 10318 15144 10324 15156
rect 9723 15116 10324 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 11698 15104 11704 15156
rect 11756 15144 11762 15156
rect 12023 15147 12081 15153
rect 12023 15144 12035 15147
rect 11756 15116 12035 15144
rect 11756 15104 11762 15116
rect 12023 15113 12035 15116
rect 12069 15144 12081 15147
rect 12894 15144 12900 15156
rect 12069 15116 12900 15144
rect 12069 15113 12081 15116
rect 12023 15107 12081 15113
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 13446 15144 13452 15156
rect 13407 15116 13452 15144
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 14458 15104 14464 15156
rect 14516 15144 14522 15156
rect 15194 15144 15200 15156
rect 14516 15116 15200 15144
rect 14516 15104 14522 15116
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 15654 15144 15660 15156
rect 15615 15116 15660 15144
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 18049 15147 18107 15153
rect 16040 15116 16620 15144
rect 7101 15079 7159 15085
rect 7101 15076 7113 15079
rect 6788 15048 7113 15076
rect 6788 15036 6794 15048
rect 7101 15045 7113 15048
rect 7147 15045 7159 15079
rect 7101 15039 7159 15045
rect 7193 15079 7251 15085
rect 7193 15045 7205 15079
rect 7239 15076 7251 15079
rect 10042 15076 10048 15088
rect 7239 15048 10048 15076
rect 7239 15045 7251 15048
rect 7193 15039 7251 15045
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 13265 15079 13323 15085
rect 13265 15045 13277 15079
rect 13311 15076 13323 15079
rect 16040 15076 16068 15116
rect 13311 15048 16068 15076
rect 13311 15045 13323 15048
rect 13265 15039 13323 15045
rect 16206 15036 16212 15088
rect 16264 15076 16270 15088
rect 16485 15079 16543 15085
rect 16485 15076 16497 15079
rect 16264 15048 16497 15076
rect 16264 15036 16270 15048
rect 16485 15045 16497 15048
rect 16531 15045 16543 15079
rect 16592 15076 16620 15116
rect 18049 15113 18061 15147
rect 18095 15144 18107 15147
rect 18138 15144 18144 15156
rect 18095 15116 18144 15144
rect 18095 15113 18107 15116
rect 18049 15107 18107 15113
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 18509 15147 18567 15153
rect 18509 15113 18521 15147
rect 18555 15144 18567 15147
rect 18598 15144 18604 15156
rect 18555 15116 18604 15144
rect 18555 15113 18567 15116
rect 18509 15107 18567 15113
rect 18322 15076 18328 15088
rect 16592 15048 18328 15076
rect 16485 15039 16543 15045
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 18524 15076 18552 15107
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15144 18751 15147
rect 19610 15144 19616 15156
rect 18739 15116 19616 15144
rect 18739 15113 18751 15116
rect 18693 15107 18751 15113
rect 19610 15104 19616 15116
rect 19668 15104 19674 15156
rect 19978 15144 19984 15156
rect 19812 15116 19984 15144
rect 19242 15076 19248 15088
rect 18524 15048 19248 15076
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 19334 15036 19340 15088
rect 19392 15076 19398 15088
rect 19812 15076 19840 15116
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 20257 15147 20315 15153
rect 20257 15144 20269 15147
rect 20220 15116 20269 15144
rect 20220 15104 20226 15116
rect 20257 15113 20269 15116
rect 20303 15113 20315 15147
rect 20257 15107 20315 15113
rect 20441 15147 20499 15153
rect 20441 15113 20453 15147
rect 20487 15144 20499 15147
rect 20622 15144 20628 15156
rect 20487 15116 20628 15144
rect 20487 15113 20499 15116
rect 20441 15107 20499 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 22922 15104 22928 15156
rect 22980 15144 22986 15156
rect 23109 15147 23167 15153
rect 23109 15144 23121 15147
rect 22980 15116 23121 15144
rect 22980 15104 22986 15116
rect 23109 15113 23121 15116
rect 23155 15113 23167 15147
rect 23109 15107 23167 15113
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 23845 15147 23903 15153
rect 23845 15144 23857 15147
rect 23808 15116 23857 15144
rect 23808 15104 23814 15116
rect 23845 15113 23857 15116
rect 23891 15113 23903 15147
rect 23845 15107 23903 15113
rect 24302 15104 24308 15156
rect 24360 15144 24366 15156
rect 24489 15147 24547 15153
rect 24489 15144 24501 15147
rect 24360 15116 24501 15144
rect 24360 15104 24366 15116
rect 24489 15113 24501 15116
rect 24535 15113 24547 15147
rect 24489 15107 24547 15113
rect 24854 15104 24860 15156
rect 24912 15144 24918 15156
rect 25041 15147 25099 15153
rect 25041 15144 25053 15147
rect 24912 15116 25053 15144
rect 24912 15104 24918 15116
rect 25041 15113 25053 15116
rect 25087 15113 25099 15147
rect 25774 15144 25780 15156
rect 25735 15116 25780 15144
rect 25041 15107 25099 15113
rect 25774 15104 25780 15116
rect 25832 15104 25838 15156
rect 27062 15104 27068 15156
rect 27120 15144 27126 15156
rect 27617 15147 27675 15153
rect 27617 15144 27629 15147
rect 27120 15116 27629 15144
rect 27120 15104 27126 15116
rect 27617 15113 27629 15116
rect 27663 15113 27675 15147
rect 28350 15144 28356 15156
rect 28311 15116 28356 15144
rect 27617 15107 27675 15113
rect 19392 15048 19840 15076
rect 19889 15079 19947 15085
rect 19392 15036 19398 15048
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20346 15076 20352 15088
rect 19935 15048 20352 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 23658 15036 23664 15088
rect 23716 15036 23722 15088
rect 24578 15036 24584 15088
rect 24636 15076 24642 15088
rect 24946 15076 24952 15088
rect 24636 15048 24952 15076
rect 24636 15036 24642 15048
rect 24946 15036 24952 15048
rect 25004 15036 25010 15088
rect 27632 15076 27660 15107
rect 28350 15104 28356 15116
rect 28408 15104 28414 15156
rect 29641 15147 29699 15153
rect 29641 15113 29653 15147
rect 29687 15144 29699 15147
rect 30006 15144 30012 15156
rect 29687 15116 30012 15144
rect 29687 15113 29699 15116
rect 29641 15107 29699 15113
rect 30006 15104 30012 15116
rect 30064 15104 30070 15156
rect 28718 15076 28724 15088
rect 25056 15048 27108 15076
rect 27632 15048 28724 15076
rect 7282 15008 7288 15020
rect 6656 14980 7144 15008
rect 7243 14980 7288 15008
rect 6181 14971 6239 14977
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2593 14943 2651 14949
rect 2593 14940 2605 14943
rect 2280 14912 2605 14940
rect 2280 14900 2286 14912
rect 2593 14909 2605 14912
rect 2639 14909 2651 14943
rect 4798 14940 4804 14952
rect 4759 14912 4804 14940
rect 2593 14903 2651 14909
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 5074 14940 5080 14952
rect 5035 14912 5080 14940
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 5810 14940 5816 14952
rect 5771 14912 5816 14940
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 1762 14832 1768 14884
rect 1820 14872 1826 14884
rect 3234 14872 3240 14884
rect 1820 14844 3240 14872
rect 1820 14832 1826 14844
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 3881 14875 3939 14881
rect 3881 14841 3893 14875
rect 3927 14872 3939 14875
rect 5258 14872 5264 14884
rect 3927 14844 5264 14872
rect 3927 14841 3939 14844
rect 3881 14835 3939 14841
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 6196 14872 6224 14971
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14909 7067 14943
rect 7116 14940 7144 14980
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 7637 14980 8064 15008
rect 7637 14940 7665 14980
rect 7742 14940 7748 14952
rect 7116 14912 7665 14940
rect 7703 14912 7748 14940
rect 7009 14903 7067 14909
rect 7024 14872 7052 14903
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 8036 14949 8064 14980
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8720 14980 8953 15008
rect 8720 14968 8726 14980
rect 8941 14977 8953 14980
rect 8987 15008 8999 15011
rect 8987 14980 9260 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14940 8171 14943
rect 8202 14940 8208 14952
rect 8159 14912 8208 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 7190 14872 7196 14884
rect 6196 14844 6960 14872
rect 7024 14844 7196 14872
rect 2406 14764 2412 14816
rect 2464 14804 2470 14816
rect 2590 14804 2596 14816
rect 2464 14776 2596 14804
rect 2464 14764 2470 14776
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 4081 14807 4139 14813
rect 4081 14804 4093 14807
rect 3844 14776 4093 14804
rect 3844 14764 3850 14776
rect 4081 14773 4093 14776
rect 4127 14773 4139 14807
rect 4246 14804 4252 14816
rect 4207 14776 4252 14804
rect 4081 14767 4139 14773
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 6932 14804 6960 14844
rect 7190 14832 7196 14844
rect 7248 14832 7254 14884
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 7944 14872 7972 14903
rect 7616 14844 7972 14872
rect 8036 14872 8064 14903
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 9232 14940 9260 14980
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 9824 14980 19840 15008
rect 9824 14968 9830 14980
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 9232 14912 9505 14940
rect 9493 14909 9505 14912
rect 9539 14940 9551 14943
rect 9674 14940 9680 14952
rect 9539 14912 9680 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 10192 14912 10241 14940
rect 10192 14900 10198 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 11054 14940 11060 14952
rect 10551 14912 11060 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14909 11851 14943
rect 13538 14940 13544 14952
rect 13499 14912 13544 14940
rect 11793 14903 11851 14909
rect 8036 14844 8156 14872
rect 7616 14832 7622 14844
rect 8018 14804 8024 14816
rect 6932 14776 8024 14804
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8128 14804 8156 14844
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 9766 14872 9772 14884
rect 8812 14844 9772 14872
rect 8812 14832 8818 14844
rect 9766 14832 9772 14844
rect 9824 14832 9830 14884
rect 10778 14832 10784 14884
rect 10836 14872 10842 14884
rect 11808 14872 11836 14903
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 14516 14912 16313 14940
rect 14516 14900 14522 14912
rect 16301 14909 16313 14912
rect 16347 14940 16359 14943
rect 17034 14940 17040 14952
rect 16347 14912 17040 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14909 17187 14943
rect 18138 14940 18144 14952
rect 18099 14912 18144 14940
rect 17129 14903 17187 14909
rect 14185 14875 14243 14881
rect 14185 14872 14197 14875
rect 10836 14844 14197 14872
rect 10836 14832 10842 14844
rect 14185 14841 14197 14844
rect 14231 14872 14243 14875
rect 15562 14872 15568 14884
rect 14231 14844 15568 14872
rect 14231 14841 14243 14844
rect 14185 14835 14243 14841
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 15654 14832 15660 14884
rect 15712 14872 15718 14884
rect 15930 14872 15936 14884
rect 15712 14844 15936 14872
rect 15712 14832 15718 14844
rect 15930 14832 15936 14844
rect 15988 14872 15994 14884
rect 15988 14844 16712 14872
rect 15988 14832 15994 14844
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 8128 14776 13277 14804
rect 13265 14773 13277 14776
rect 13311 14773 13323 14807
rect 13265 14767 13323 14773
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 14645 14807 14703 14813
rect 14645 14804 14657 14807
rect 13872 14776 14657 14804
rect 13872 14764 13878 14776
rect 14645 14773 14657 14776
rect 14691 14773 14703 14807
rect 14645 14767 14703 14773
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16298 14804 16304 14816
rect 15804 14776 16304 14804
rect 15804 14764 15810 14776
rect 16298 14764 16304 14776
rect 16356 14764 16362 14816
rect 16684 14804 16712 14844
rect 16758 14832 16764 14884
rect 16816 14872 16822 14884
rect 17144 14872 17172 14903
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 18380 14912 18552 14940
rect 18380 14900 18386 14912
rect 16816 14844 17172 14872
rect 17405 14875 17463 14881
rect 16816 14832 16822 14844
rect 17405 14841 17417 14875
rect 17451 14872 17463 14875
rect 18414 14872 18420 14884
rect 17451 14844 18420 14872
rect 17451 14841 17463 14844
rect 17405 14835 17463 14841
rect 18414 14832 18420 14844
rect 18472 14832 18478 14884
rect 18524 14872 18552 14912
rect 18966 14900 18972 14952
rect 19024 14940 19030 14952
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 19024 14912 19257 14940
rect 19024 14900 19030 14912
rect 19245 14909 19257 14912
rect 19291 14909 19303 14943
rect 19245 14903 19303 14909
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 19392 14912 19441 14940
rect 19392 14900 19398 14912
rect 19429 14909 19441 14912
rect 19475 14909 19487 14943
rect 19812 14940 19840 14980
rect 20806 14968 20812 15020
rect 20864 15008 20870 15020
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 20864 14980 21189 15008
rect 20864 14968 20870 14980
rect 21177 14977 21189 14980
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 22830 14968 22836 15020
rect 22888 15008 22894 15020
rect 23676 15008 23704 15036
rect 22888 14980 24624 15008
rect 22888 14968 22894 14980
rect 19812 14912 23060 14940
rect 19429 14903 19487 14909
rect 19610 14872 19616 14884
rect 18524 14844 19616 14872
rect 19610 14832 19616 14844
rect 19668 14832 19674 14884
rect 20162 14832 20168 14884
rect 20220 14872 20226 14884
rect 21450 14881 21456 14884
rect 20257 14875 20315 14881
rect 20257 14872 20269 14875
rect 20220 14844 20269 14872
rect 20220 14832 20226 14844
rect 20257 14841 20269 14844
rect 20303 14841 20315 14875
rect 20257 14835 20315 14841
rect 21444 14835 21456 14881
rect 21508 14872 21514 14884
rect 21508 14844 21544 14872
rect 21450 14832 21456 14835
rect 21508 14832 21514 14844
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 16684 14776 18061 14804
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 18049 14767 18107 14773
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 18509 14807 18567 14813
rect 18509 14804 18521 14807
rect 18288 14776 18521 14804
rect 18288 14764 18294 14776
rect 18509 14773 18521 14776
rect 18555 14773 18567 14807
rect 18509 14767 18567 14773
rect 19337 14807 19395 14813
rect 19337 14773 19349 14807
rect 19383 14804 19395 14807
rect 19886 14804 19892 14816
rect 19383 14776 19892 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 22462 14804 22468 14816
rect 20036 14776 22468 14804
rect 20036 14764 20042 14776
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 22557 14807 22615 14813
rect 22557 14773 22569 14807
rect 22603 14804 22615 14807
rect 22646 14804 22652 14816
rect 22603 14776 22652 14804
rect 22603 14773 22615 14776
rect 22557 14767 22615 14773
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 23032 14804 23060 14912
rect 23106 14900 23112 14952
rect 23164 14940 23170 14952
rect 23201 14943 23259 14949
rect 23201 14940 23213 14943
rect 23164 14912 23213 14940
rect 23164 14900 23170 14912
rect 23201 14909 23213 14912
rect 23247 14909 23259 14943
rect 23201 14903 23259 14909
rect 23661 14943 23719 14949
rect 23661 14909 23673 14943
rect 23707 14940 23719 14943
rect 23750 14940 23756 14952
rect 23707 14912 23756 14940
rect 23707 14909 23719 14912
rect 23661 14903 23719 14909
rect 23750 14900 23756 14912
rect 23808 14900 23814 14952
rect 23845 14943 23903 14949
rect 23845 14909 23857 14943
rect 23891 14942 23903 14943
rect 23891 14914 23980 14942
rect 23891 14909 23903 14914
rect 23845 14903 23903 14909
rect 23952 14872 23980 14914
rect 24026 14900 24032 14952
rect 24084 14940 24090 14952
rect 24596 14949 24624 14980
rect 24670 14968 24676 15020
rect 24728 15008 24734 15020
rect 25056 15008 25084 15048
rect 26602 15008 26608 15020
rect 24728 14980 25084 15008
rect 25976 14980 26608 15008
rect 24728 14968 24734 14980
rect 25976 14949 26004 14980
rect 26602 14968 26608 14980
rect 26660 14968 26666 15020
rect 24397 14943 24455 14949
rect 24397 14940 24409 14943
rect 24084 14912 24409 14940
rect 24084 14900 24090 14912
rect 24397 14909 24409 14912
rect 24443 14909 24455 14943
rect 24397 14903 24455 14909
rect 24581 14943 24639 14949
rect 24581 14909 24593 14943
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 25961 14943 26019 14949
rect 25961 14909 25973 14943
rect 26007 14909 26019 14943
rect 26142 14940 26148 14952
rect 26103 14912 26148 14940
rect 25961 14903 26019 14909
rect 26142 14900 26148 14912
rect 26200 14900 26206 14952
rect 26237 14943 26295 14949
rect 26237 14909 26249 14943
rect 26283 14909 26295 14943
rect 26237 14903 26295 14909
rect 24762 14872 24768 14884
rect 23952 14844 24768 14872
rect 24762 14832 24768 14844
rect 24820 14832 24826 14884
rect 24854 14804 24860 14816
rect 23032 14776 24860 14804
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 25958 14764 25964 14816
rect 26016 14804 26022 14816
rect 26252 14804 26280 14903
rect 26326 14900 26332 14952
rect 26384 14940 26390 14952
rect 26384 14912 26429 14940
rect 26384 14900 26390 14912
rect 26510 14900 26516 14952
rect 26568 14940 26574 14952
rect 26568 14912 26613 14940
rect 26568 14900 26574 14912
rect 27080 14813 27108 15048
rect 28718 15036 28724 15048
rect 28776 15036 28782 15088
rect 28813 15079 28871 15085
rect 28813 15045 28825 15079
rect 28859 15045 28871 15079
rect 28813 15039 28871 15045
rect 28169 14943 28227 14949
rect 28169 14909 28181 14943
rect 28215 14940 28227 14943
rect 28828 14940 28856 15039
rect 28215 14912 28856 14940
rect 28997 14943 29055 14949
rect 28215 14909 28227 14912
rect 28169 14903 28227 14909
rect 28997 14909 29009 14943
rect 29043 14909 29055 14943
rect 28997 14903 29055 14909
rect 29012 14872 29040 14903
rect 29730 14900 29736 14952
rect 29788 14940 29794 14952
rect 31021 14943 31079 14949
rect 31021 14940 31033 14943
rect 29788 14912 31033 14940
rect 29788 14900 29794 14912
rect 31021 14909 31033 14912
rect 31067 14909 31079 14943
rect 31021 14903 31079 14909
rect 30282 14872 30288 14884
rect 29012 14844 30288 14872
rect 30282 14832 30288 14844
rect 30340 14832 30346 14884
rect 30374 14832 30380 14884
rect 30432 14872 30438 14884
rect 30754 14875 30812 14881
rect 30754 14872 30766 14875
rect 30432 14844 30766 14872
rect 30432 14832 30438 14844
rect 30754 14841 30766 14844
rect 30800 14841 30812 14875
rect 30754 14835 30812 14841
rect 26016 14776 26280 14804
rect 27065 14807 27123 14813
rect 26016 14764 26022 14776
rect 27065 14773 27077 14807
rect 27111 14804 27123 14807
rect 30558 14804 30564 14816
rect 27111 14776 30564 14804
rect 27111 14773 27123 14776
rect 27065 14767 27123 14773
rect 30558 14764 30564 14776
rect 30616 14764 30622 14816
rect 1104 14714 32016 14736
rect 1104 14662 11253 14714
rect 11305 14662 11317 14714
rect 11369 14662 11381 14714
rect 11433 14662 11445 14714
rect 11497 14662 11509 14714
rect 11561 14662 21557 14714
rect 21609 14662 21621 14714
rect 21673 14662 21685 14714
rect 21737 14662 21749 14714
rect 21801 14662 21813 14714
rect 21865 14662 32016 14714
rect 1104 14640 32016 14662
rect 2590 14560 2596 14612
rect 2648 14600 2654 14612
rect 2774 14600 2780 14612
rect 2648 14572 2780 14600
rect 2648 14560 2654 14572
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 3789 14603 3847 14609
rect 3292 14572 3372 14600
rect 3292 14560 3298 14572
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 2866 14532 2872 14544
rect 2188 14504 2872 14532
rect 2188 14492 2194 14504
rect 2866 14492 2872 14504
rect 2924 14532 2930 14544
rect 3344 14532 3372 14572
rect 3789 14569 3801 14603
rect 3835 14600 3847 14603
rect 5626 14600 5632 14612
rect 3835 14572 5632 14600
rect 3835 14569 3847 14572
rect 3789 14563 3847 14569
rect 5626 14560 5632 14572
rect 5684 14560 5690 14612
rect 7650 14600 7656 14612
rect 7611 14572 7656 14600
rect 7650 14560 7656 14572
rect 7708 14600 7714 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 7708 14572 8493 14600
rect 7708 14560 7714 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 8938 14600 8944 14612
rect 8899 14572 8944 14600
rect 8481 14563 8539 14569
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 10134 14600 10140 14612
rect 10095 14572 10140 14600
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10594 14600 10600 14612
rect 10555 14572 10600 14600
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12250 14600 12256 14612
rect 12207 14572 12256 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12250 14560 12256 14572
rect 12308 14600 12314 14612
rect 12618 14600 12624 14612
rect 12308 14572 12624 14600
rect 12308 14560 12314 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 19058 14600 19064 14612
rect 15804 14572 19064 14600
rect 15804 14560 15810 14572
rect 19058 14560 19064 14572
rect 19116 14560 19122 14612
rect 19153 14603 19211 14609
rect 19153 14569 19165 14603
rect 19199 14600 19211 14603
rect 19242 14600 19248 14612
rect 19199 14572 19248 14600
rect 19199 14569 19211 14572
rect 19153 14563 19211 14569
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19978 14600 19984 14612
rect 19352 14572 19984 14600
rect 4154 14532 4160 14544
rect 2924 14504 3280 14532
rect 3344 14504 4160 14532
rect 2924 14492 2930 14504
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14464 2375 14467
rect 2774 14464 2780 14476
rect 2363 14436 2780 14464
rect 2363 14433 2375 14436
rect 2317 14427 2375 14433
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 3053 14467 3111 14473
rect 3053 14433 3065 14467
rect 3099 14464 3111 14467
rect 3145 14467 3203 14473
rect 3145 14464 3157 14467
rect 3099 14436 3157 14464
rect 3099 14433 3111 14436
rect 3053 14427 3111 14433
rect 3145 14433 3157 14436
rect 3191 14433 3203 14467
rect 3252 14464 3280 14504
rect 3528 14473 3556 14504
rect 4154 14492 4160 14504
rect 4212 14532 4218 14544
rect 4433 14535 4491 14541
rect 4212 14504 4384 14532
rect 4212 14492 4218 14504
rect 3329 14467 3387 14473
rect 3329 14464 3341 14467
rect 3252 14436 3341 14464
rect 3145 14427 3203 14433
rect 3329 14433 3341 14436
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 3513 14467 3571 14473
rect 3513 14433 3525 14467
rect 3559 14433 3571 14467
rect 4246 14464 4252 14476
rect 4207 14436 4252 14464
rect 3513 14427 3571 14433
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2593 14399 2651 14405
rect 2593 14396 2605 14399
rect 2464 14368 2605 14396
rect 2464 14356 2470 14368
rect 2593 14365 2605 14368
rect 2639 14365 2651 14399
rect 3436 14396 3464 14427
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 4356 14464 4384 14504
rect 4433 14501 4445 14535
rect 4479 14532 4491 14535
rect 5074 14532 5080 14544
rect 4479 14504 5080 14532
rect 4479 14501 4491 14504
rect 4433 14495 4491 14501
rect 5074 14492 5080 14504
rect 5132 14492 5138 14544
rect 5994 14532 6000 14544
rect 5644 14504 6000 14532
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 4356 14436 4537 14464
rect 4525 14433 4537 14436
rect 4571 14433 4583 14467
rect 4982 14464 4988 14476
rect 4943 14436 4988 14464
rect 4525 14427 4583 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5258 14424 5264 14476
rect 5316 14464 5322 14476
rect 5644 14473 5672 14504
rect 5994 14492 6000 14504
rect 6052 14492 6058 14544
rect 6564 14504 7788 14532
rect 6564 14473 6592 14504
rect 5629 14467 5687 14473
rect 5629 14464 5641 14467
rect 5316 14436 5641 14464
rect 5316 14424 5322 14436
rect 5629 14433 5641 14436
rect 5675 14433 5687 14467
rect 5629 14427 5687 14433
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14464 5871 14467
rect 6549 14467 6607 14473
rect 5859 14436 6500 14464
rect 5859 14433 5871 14436
rect 5813 14427 5871 14433
rect 6472 14408 6500 14436
rect 6549 14433 6561 14467
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 6696 14436 6745 14464
rect 6696 14424 6702 14436
rect 6733 14433 6745 14436
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 3878 14396 3884 14408
rect 3436 14368 3884 14396
rect 2593 14359 2651 14365
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4338 14396 4344 14408
rect 4120 14368 4344 14396
rect 4120 14356 4126 14368
rect 4338 14356 4344 14368
rect 4396 14396 4402 14408
rect 4801 14399 4859 14405
rect 4801 14396 4813 14399
rect 4396 14368 4813 14396
rect 4396 14356 4402 14368
rect 4801 14365 4813 14368
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 3053 14331 3111 14337
rect 3053 14297 3065 14331
rect 3099 14328 3111 14331
rect 4816 14328 4844 14359
rect 5074 14356 5080 14408
rect 5132 14396 5138 14408
rect 5350 14396 5356 14408
rect 5132 14368 5356 14396
rect 5132 14356 5138 14368
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 6454 14356 6460 14408
rect 6512 14396 6518 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6512 14368 6837 14396
rect 6512 14356 6518 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6932 14396 6960 14427
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7101 14467 7159 14473
rect 7101 14464 7113 14467
rect 7064 14436 7113 14464
rect 7064 14424 7070 14436
rect 7101 14433 7113 14436
rect 7147 14433 7159 14467
rect 7558 14464 7564 14476
rect 7519 14436 7564 14464
rect 7101 14427 7159 14433
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 7760 14473 7788 14504
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 7892 14504 9444 14532
rect 7892 14492 7898 14504
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14464 7803 14467
rect 8110 14464 8116 14476
rect 7791 14436 8116 14464
rect 7791 14433 7803 14436
rect 7745 14427 7803 14433
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 9416 14473 9444 14504
rect 12066 14492 12072 14544
rect 12124 14532 12130 14544
rect 14366 14532 14372 14544
rect 12124 14504 14372 14532
rect 12124 14492 12130 14504
rect 13096 14473 13124 14504
rect 14366 14492 14372 14504
rect 14424 14492 14430 14544
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 15252 14504 15700 14532
rect 15252 14492 15258 14504
rect 15672 14486 15700 14504
rect 16850 14492 16856 14544
rect 16908 14532 16914 14544
rect 18046 14541 18052 14544
rect 17037 14535 17095 14541
rect 17037 14532 17049 14535
rect 16908 14504 17049 14532
rect 16908 14492 16914 14504
rect 17037 14501 17049 14504
rect 17083 14501 17095 14535
rect 17037 14495 17095 14501
rect 18040 14495 18052 14541
rect 18104 14532 18110 14544
rect 18104 14504 18140 14532
rect 18046 14492 18052 14495
rect 18104 14492 18110 14504
rect 13354 14473 13360 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8536 14436 8585 14464
rect 8536 14424 8542 14436
rect 8573 14433 8585 14436
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 9401 14467 9459 14473
rect 9401 14433 9413 14467
rect 9447 14433 9459 14467
rect 9401 14427 9459 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 13081 14467 13139 14473
rect 13081 14433 13093 14467
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 13348 14427 13360 14473
rect 13412 14464 13418 14476
rect 13412 14436 13448 14464
rect 6932 14368 7144 14396
rect 6825 14359 6883 14365
rect 7116 14340 7144 14368
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 8202 14396 8208 14408
rect 7432 14368 8208 14396
rect 7432 14356 7438 14368
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14365 8447 14399
rect 8588 14396 8616 14427
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 8588 14368 9505 14396
rect 8389 14359 8447 14365
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 5810 14328 5816 14340
rect 3099 14300 4292 14328
rect 4816 14300 5816 14328
rect 3099 14297 3111 14300
rect 3053 14291 3111 14297
rect 4264 14272 4292 14300
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 6730 14328 6736 14340
rect 6288 14300 6736 14328
rect 4246 14220 4252 14272
rect 4304 14220 4310 14272
rect 4522 14220 4528 14272
rect 4580 14260 4586 14272
rect 5534 14260 5540 14272
rect 4580 14232 5540 14260
rect 4580 14220 4586 14232
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 6288 14260 6316 14300
rect 6730 14288 6736 14300
rect 6788 14288 6794 14340
rect 7098 14288 7104 14340
rect 7156 14288 7162 14340
rect 8404 14328 8432 14359
rect 8754 14328 8760 14340
rect 8404 14300 8760 14328
rect 8754 14288 8760 14300
rect 8812 14288 8818 14340
rect 5684 14232 6316 14260
rect 6365 14263 6423 14269
rect 5684 14220 5690 14232
rect 6365 14229 6377 14263
rect 6411 14260 6423 14263
rect 6454 14260 6460 14272
rect 6411 14232 6460 14260
rect 6411 14229 6423 14232
rect 6365 14223 6423 14229
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 9600 14260 9628 14427
rect 13354 14424 13360 14427
rect 13412 14424 13418 14436
rect 14642 14424 14648 14476
rect 14700 14464 14706 14476
rect 14921 14467 14979 14473
rect 14921 14464 14933 14467
rect 14700 14436 14933 14464
rect 14700 14424 14706 14436
rect 14921 14433 14933 14436
rect 14967 14433 14979 14467
rect 15102 14464 15108 14476
rect 15063 14436 15108 14464
rect 14921 14427 14979 14433
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 15286 14464 15292 14476
rect 15247 14436 15292 14464
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 15672 14464 15884 14486
rect 19352 14464 19380 14572
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 21177 14603 21235 14609
rect 21177 14569 21189 14603
rect 21223 14569 21235 14603
rect 21177 14563 21235 14569
rect 20806 14532 20812 14544
rect 19812 14504 20812 14532
rect 15528 14436 15573 14464
rect 15672 14458 19380 14464
rect 15856 14436 19380 14458
rect 15528 14424 15534 14436
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 19812 14473 19840 14504
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 19576 14436 19809 14464
rect 19576 14424 19582 14436
rect 19797 14433 19809 14436
rect 19843 14433 19855 14467
rect 19797 14427 19855 14433
rect 19886 14424 19892 14476
rect 19944 14464 19950 14476
rect 20053 14467 20111 14473
rect 20053 14464 20065 14467
rect 19944 14436 20065 14464
rect 19944 14424 19950 14436
rect 20053 14433 20065 14436
rect 20099 14433 20111 14467
rect 21192 14464 21220 14563
rect 22462 14560 22468 14612
rect 22520 14600 22526 14612
rect 24026 14600 24032 14612
rect 22520 14572 23612 14600
rect 23987 14572 24032 14600
rect 22520 14560 22526 14572
rect 23474 14532 23480 14544
rect 22664 14504 23480 14532
rect 22664 14473 22692 14504
rect 23474 14492 23480 14504
rect 23532 14492 23538 14544
rect 23584 14532 23612 14572
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 24670 14560 24676 14612
rect 24728 14560 24734 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 27617 14603 27675 14609
rect 27617 14600 27629 14603
rect 24912 14572 27629 14600
rect 24912 14560 24918 14572
rect 27617 14569 27629 14572
rect 27663 14569 27675 14603
rect 28442 14600 28448 14612
rect 28355 14572 28448 14600
rect 27617 14563 27675 14569
rect 28442 14560 28448 14572
rect 28500 14600 28506 14612
rect 28718 14600 28724 14612
rect 28500 14572 28724 14600
rect 28500 14560 28506 14572
rect 28718 14560 28724 14572
rect 28776 14560 28782 14612
rect 30374 14600 30380 14612
rect 30335 14572 30380 14600
rect 30374 14560 30380 14572
rect 30432 14560 30438 14612
rect 31297 14603 31355 14609
rect 31297 14569 31309 14603
rect 31343 14600 31355 14603
rect 31478 14600 31484 14612
rect 31343 14572 31484 14600
rect 31343 14569 31355 14572
rect 31297 14563 31355 14569
rect 31478 14560 31484 14572
rect 31536 14560 31542 14612
rect 24688 14532 24716 14560
rect 23584 14504 24716 14532
rect 25130 14492 25136 14544
rect 25188 14532 25194 14544
rect 26142 14532 26148 14544
rect 25188 14504 26148 14532
rect 25188 14492 25194 14504
rect 26142 14492 26148 14504
rect 26200 14492 26206 14544
rect 21981 14467 22039 14473
rect 21981 14464 21993 14467
rect 21192 14436 21993 14464
rect 20053 14427 20111 14433
rect 21981 14433 21993 14436
rect 22027 14464 22039 14467
rect 22649 14467 22707 14473
rect 22027 14433 22048 14464
rect 21981 14427 22048 14433
rect 22649 14433 22661 14467
rect 22695 14433 22707 14467
rect 22649 14427 22707 14433
rect 22916 14467 22974 14473
rect 22916 14433 22928 14467
rect 22962 14464 22974 14467
rect 23382 14464 23388 14476
rect 22962 14436 23388 14464
rect 22962 14433 22974 14436
rect 22916 14427 22974 14433
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14396 15255 14399
rect 15378 14396 15384 14408
rect 15243 14368 15384 14396
rect 15243 14365 15255 14368
rect 15197 14359 15255 14365
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14396 16727 14399
rect 16758 14396 16764 14408
rect 16715 14368 16764 14396
rect 16715 14365 16727 14368
rect 16669 14359 16727 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 17770 14396 17776 14408
rect 17731 14368 17776 14396
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 22020 14396 22048 14427
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 24489 14467 24547 14473
rect 24489 14433 24501 14467
rect 24535 14464 24547 14467
rect 24578 14464 24584 14476
rect 24535 14436 24584 14464
rect 24535 14433 24547 14436
rect 24489 14427 24547 14433
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14464 24731 14467
rect 24946 14464 24952 14476
rect 24719 14436 24952 14464
rect 24719 14433 24731 14436
rect 24673 14427 24731 14433
rect 24946 14424 24952 14436
rect 25004 14424 25010 14476
rect 25041 14467 25099 14473
rect 25041 14433 25053 14467
rect 25087 14464 25099 14467
rect 25314 14464 25320 14476
rect 25087 14436 25320 14464
rect 25087 14433 25099 14436
rect 25041 14427 25099 14433
rect 25314 14424 25320 14436
rect 25372 14424 25378 14476
rect 25590 14424 25596 14476
rect 25648 14464 25654 14476
rect 25685 14467 25743 14473
rect 25685 14464 25697 14467
rect 25648 14436 25697 14464
rect 25648 14424 25654 14436
rect 25685 14433 25697 14436
rect 25731 14433 25743 14467
rect 25685 14427 25743 14433
rect 25869 14467 25927 14473
rect 25869 14433 25881 14467
rect 25915 14433 25927 14467
rect 25869 14427 25927 14433
rect 24762 14396 24768 14408
rect 22020 14368 22692 14396
rect 24675 14368 24768 14396
rect 14090 14288 14096 14340
rect 14148 14328 14154 14340
rect 14461 14331 14519 14337
rect 14461 14328 14473 14331
rect 14148 14300 14473 14328
rect 14148 14288 14154 14300
rect 14461 14297 14473 14300
rect 14507 14328 14519 14331
rect 17402 14328 17408 14340
rect 14507 14300 17408 14328
rect 14507 14297 14519 14300
rect 14461 14291 14519 14297
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 19518 14328 19524 14340
rect 18708 14300 19524 14328
rect 7984 14232 9628 14260
rect 11609 14263 11667 14269
rect 7984 14220 7990 14232
rect 11609 14229 11621 14263
rect 11655 14260 11667 14263
rect 12250 14260 12256 14272
rect 11655 14232 12256 14260
rect 11655 14229 11667 14232
rect 11609 14223 11667 14229
rect 12250 14220 12256 14232
rect 12308 14260 12314 14272
rect 13998 14260 14004 14272
rect 12308 14232 14004 14260
rect 12308 14220 12314 14232
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 16850 14260 16856 14272
rect 14976 14232 16856 14260
rect 14976 14220 14982 14232
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 17037 14263 17095 14269
rect 17037 14229 17049 14263
rect 17083 14260 17095 14263
rect 17126 14260 17132 14272
rect 17083 14232 17132 14260
rect 17083 14229 17095 14232
rect 17037 14223 17095 14229
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 17221 14263 17279 14269
rect 17221 14229 17233 14263
rect 17267 14260 17279 14263
rect 17954 14260 17960 14272
rect 17267 14232 17960 14260
rect 17267 14229 17279 14232
rect 17221 14223 17279 14229
rect 17954 14220 17960 14232
rect 18012 14220 18018 14272
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18708 14260 18736 14300
rect 19518 14288 19524 14300
rect 19576 14288 19582 14340
rect 18104 14232 18736 14260
rect 18104 14220 18110 14232
rect 19058 14220 19064 14272
rect 19116 14260 19122 14272
rect 21174 14260 21180 14272
rect 19116 14232 21180 14260
rect 19116 14220 19122 14232
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 21913 14263 21971 14269
rect 21913 14260 21925 14263
rect 21692 14232 21925 14260
rect 21692 14220 21698 14232
rect 21913 14229 21925 14232
rect 21959 14229 21971 14263
rect 22664 14260 22692 14368
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 24857 14399 24915 14405
rect 24857 14365 24869 14399
rect 24903 14396 24915 14399
rect 25130 14396 25136 14408
rect 24903 14368 25136 14396
rect 24903 14365 24915 14368
rect 24857 14359 24915 14365
rect 25130 14356 25136 14368
rect 25188 14356 25194 14408
rect 25332 14396 25360 14424
rect 25884 14396 25912 14427
rect 25958 14424 25964 14476
rect 26016 14464 26022 14476
rect 26237 14467 26295 14473
rect 26016 14436 26061 14464
rect 26016 14424 26022 14436
rect 26237 14433 26249 14467
rect 26283 14464 26295 14467
rect 26326 14464 26332 14476
rect 26283 14436 26332 14464
rect 26283 14433 26295 14436
rect 26237 14427 26295 14433
rect 26326 14424 26332 14436
rect 26384 14464 26390 14476
rect 26973 14467 27031 14473
rect 26973 14464 26985 14467
rect 26384 14436 26985 14464
rect 26384 14424 26390 14436
rect 26973 14433 26985 14436
rect 27019 14464 27031 14467
rect 27154 14464 27160 14476
rect 27019 14436 27160 14464
rect 27019 14433 27031 14436
rect 26973 14427 27031 14433
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 28460 14473 28488 14560
rect 29546 14532 29552 14544
rect 28736 14504 29552 14532
rect 28445 14467 28503 14473
rect 28445 14433 28457 14467
rect 28491 14433 28503 14467
rect 28626 14464 28632 14476
rect 28587 14436 28632 14464
rect 28445 14427 28503 14433
rect 28626 14424 28632 14436
rect 28684 14424 28690 14476
rect 28736 14473 28764 14504
rect 29546 14492 29552 14504
rect 29604 14532 29610 14544
rect 29604 14504 29960 14532
rect 29604 14492 29610 14504
rect 28721 14467 28779 14473
rect 28721 14433 28733 14467
rect 28767 14433 28779 14467
rect 28997 14467 29055 14473
rect 28997 14464 29009 14467
rect 28721 14427 28779 14433
rect 28920 14436 29009 14464
rect 25332 14368 25912 14396
rect 24780 14328 24808 14356
rect 25976 14328 26004 14424
rect 26053 14399 26111 14405
rect 26053 14365 26065 14399
rect 26099 14396 26111 14399
rect 26142 14396 26148 14408
rect 26099 14368 26148 14396
rect 26099 14365 26111 14368
rect 26053 14359 26111 14365
rect 26142 14356 26148 14368
rect 26200 14356 26206 14408
rect 28166 14356 28172 14408
rect 28224 14396 28230 14408
rect 28813 14399 28871 14405
rect 28813 14396 28825 14399
rect 28224 14368 28825 14396
rect 28224 14356 28230 14368
rect 28813 14365 28825 14368
rect 28859 14365 28871 14399
rect 28813 14359 28871 14365
rect 26510 14328 26516 14340
rect 24780 14300 26004 14328
rect 26252 14300 26516 14328
rect 22922 14260 22928 14272
rect 22664 14232 22928 14260
rect 21913 14223 21971 14229
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 23290 14220 23296 14272
rect 23348 14260 23354 14272
rect 24854 14260 24860 14272
rect 23348 14232 24860 14260
rect 23348 14220 23354 14232
rect 24854 14220 24860 14232
rect 24912 14220 24918 14272
rect 25222 14260 25228 14272
rect 25183 14232 25228 14260
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 25590 14220 25596 14272
rect 25648 14260 25654 14272
rect 26252 14260 26280 14300
rect 26510 14288 26516 14300
rect 26568 14288 26574 14340
rect 28442 14288 28448 14340
rect 28500 14328 28506 14340
rect 28920 14328 28948 14436
rect 28997 14433 29009 14436
rect 29043 14433 29055 14467
rect 29638 14464 29644 14476
rect 29599 14436 29644 14464
rect 28997 14427 29055 14433
rect 29638 14424 29644 14436
rect 29696 14424 29702 14476
rect 29822 14464 29828 14476
rect 29783 14436 29828 14464
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 29932 14405 29960 14504
rect 30006 14492 30012 14544
rect 30064 14532 30070 14544
rect 30064 14504 30236 14532
rect 30064 14492 30070 14504
rect 30208 14473 30236 14504
rect 30193 14467 30251 14473
rect 30193 14433 30205 14467
rect 30239 14433 30251 14467
rect 30193 14427 30251 14433
rect 30466 14424 30472 14476
rect 30524 14464 30530 14476
rect 31110 14464 31116 14476
rect 30524 14436 31116 14464
rect 30524 14424 30530 14436
rect 31110 14424 31116 14436
rect 31168 14424 31174 14476
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14365 29975 14399
rect 29917 14359 29975 14365
rect 30009 14399 30067 14405
rect 30009 14365 30021 14399
rect 30055 14396 30067 14399
rect 30098 14396 30104 14408
rect 30055 14368 30104 14396
rect 30055 14365 30067 14368
rect 30009 14359 30067 14365
rect 28500 14300 28948 14328
rect 28500 14288 28506 14300
rect 29932 14272 29960 14359
rect 30098 14356 30104 14368
rect 30156 14356 30162 14408
rect 30742 14356 30748 14408
rect 30800 14396 30806 14408
rect 30837 14399 30895 14405
rect 30837 14396 30849 14399
rect 30800 14368 30849 14396
rect 30800 14356 30806 14368
rect 30837 14365 30849 14368
rect 30883 14365 30895 14399
rect 30837 14359 30895 14365
rect 30929 14399 30987 14405
rect 30929 14365 30941 14399
rect 30975 14396 30987 14399
rect 31202 14396 31208 14408
rect 30975 14368 31208 14396
rect 30975 14365 30987 14368
rect 30929 14359 30987 14365
rect 31202 14356 31208 14368
rect 31260 14356 31266 14408
rect 26418 14260 26424 14272
rect 25648 14232 26280 14260
rect 26379 14232 26424 14260
rect 25648 14220 25654 14232
rect 26418 14220 26424 14232
rect 26476 14220 26482 14272
rect 27062 14260 27068 14272
rect 27023 14232 27068 14260
rect 27062 14220 27068 14232
rect 27120 14220 27126 14272
rect 29178 14260 29184 14272
rect 29139 14232 29184 14260
rect 29178 14220 29184 14232
rect 29236 14220 29242 14272
rect 29914 14220 29920 14272
rect 29972 14220 29978 14272
rect 1104 14170 32016 14192
rect 1104 14118 6102 14170
rect 6154 14118 6166 14170
rect 6218 14118 6230 14170
rect 6282 14118 6294 14170
rect 6346 14118 6358 14170
rect 6410 14118 16405 14170
rect 16457 14118 16469 14170
rect 16521 14118 16533 14170
rect 16585 14118 16597 14170
rect 16649 14118 16661 14170
rect 16713 14118 26709 14170
rect 26761 14118 26773 14170
rect 26825 14118 26837 14170
rect 26889 14118 26901 14170
rect 26953 14118 26965 14170
rect 27017 14118 32016 14170
rect 1104 14096 32016 14118
rect 1489 14059 1547 14065
rect 1489 14025 1501 14059
rect 1535 14056 1547 14059
rect 1762 14056 1768 14068
rect 1535 14028 1768 14056
rect 1535 14025 1547 14028
rect 1489 14019 1547 14025
rect 1762 14016 1768 14028
rect 1820 14056 1826 14068
rect 2038 14056 2044 14068
rect 1820 14028 2044 14056
rect 1820 14016 1826 14028
rect 2038 14016 2044 14028
rect 2096 14016 2102 14068
rect 2406 14016 2412 14068
rect 2464 14056 2470 14068
rect 3145 14059 3203 14065
rect 3145 14056 3157 14059
rect 2464 14028 3157 14056
rect 2464 14016 2470 14028
rect 3145 14025 3157 14028
rect 3191 14025 3203 14059
rect 4433 14059 4491 14065
rect 3145 14019 3203 14025
rect 3988 14028 4200 14056
rect 2130 13948 2136 14000
rect 2188 13948 2194 14000
rect 2958 13948 2964 14000
rect 3016 13988 3022 14000
rect 3878 13988 3884 14000
rect 3016 13960 3884 13988
rect 3016 13948 3022 13960
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 2148 13861 2176 13948
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13920 2375 13923
rect 3326 13920 3332 13932
rect 2363 13892 3332 13920
rect 2363 13889 2375 13892
rect 2317 13883 2375 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13821 2191 13855
rect 2133 13815 2191 13821
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2409 13855 2467 13861
rect 2409 13852 2421 13855
rect 2280 13824 2421 13852
rect 2280 13812 2286 13824
rect 2409 13821 2421 13824
rect 2455 13821 2467 13855
rect 2409 13815 2467 13821
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13821 2559 13855
rect 2501 13815 2559 13821
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 2774 13852 2780 13864
rect 2731 13824 2780 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 1394 13744 1400 13796
rect 1452 13784 1458 13796
rect 2516 13784 2544 13815
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 3789 13855 3847 13861
rect 3789 13821 3801 13855
rect 3835 13852 3847 13855
rect 3878 13852 3884 13864
rect 3835 13824 3884 13852
rect 3835 13821 3847 13824
rect 3789 13815 3847 13821
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 3988 13861 4016 14028
rect 4172 13988 4200 14028
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 4890 14056 4896 14068
rect 4479 14028 4896 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 6788 14028 7205 14056
rect 6788 14016 6794 14028
rect 7193 14025 7205 14028
rect 7239 14056 7251 14059
rect 8110 14056 8116 14068
rect 7239 14028 8116 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8260 14028 9045 14056
rect 8260 14016 8266 14028
rect 9033 14025 9045 14028
rect 9079 14025 9091 14059
rect 9033 14019 9091 14025
rect 9600 14028 10565 14056
rect 4522 13988 4528 14000
rect 4172 13960 4528 13988
rect 4522 13948 4528 13960
rect 4580 13948 4586 14000
rect 7098 13948 7104 14000
rect 7156 13948 7162 14000
rect 7745 13991 7803 13997
rect 7745 13957 7757 13991
rect 7791 13988 7803 13991
rect 7926 13988 7932 14000
rect 7791 13960 7932 13988
rect 7791 13957 7803 13960
rect 7745 13951 7803 13957
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 9600 13988 9628 14028
rect 8076 13960 9628 13988
rect 10537 13988 10565 14028
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 11425 14059 11483 14065
rect 11425 14056 11437 14059
rect 10652 14028 11437 14056
rect 10652 14016 10658 14028
rect 11425 14025 11437 14028
rect 11471 14025 11483 14059
rect 11425 14019 11483 14025
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 13412 14028 13553 14056
rect 13412 14016 13418 14028
rect 13541 14025 13553 14028
rect 13587 14025 13599 14059
rect 13541 14019 13599 14025
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 16114 14056 16120 14068
rect 14424 14028 16120 14056
rect 14424 14016 14430 14028
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16850 14016 16856 14068
rect 16908 14056 16914 14068
rect 19702 14056 19708 14068
rect 16908 14028 19708 14056
rect 16908 14016 16914 14028
rect 19702 14016 19708 14028
rect 19760 14016 19766 14068
rect 20898 14016 20904 14068
rect 20956 14056 20962 14068
rect 21266 14056 21272 14068
rect 20956 14028 21272 14056
rect 20956 14016 20962 14028
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 21361 14059 21419 14065
rect 21361 14025 21373 14059
rect 21407 14056 21419 14059
rect 21450 14056 21456 14068
rect 21407 14028 21456 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 21450 14016 21456 14028
rect 21508 14016 21514 14068
rect 21910 14016 21916 14068
rect 21968 14056 21974 14068
rect 23014 14056 23020 14068
rect 21968 14028 23020 14056
rect 21968 14016 21974 14028
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 23382 14056 23388 14068
rect 23343 14028 23388 14056
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 25682 14056 25688 14068
rect 24596 14028 25688 14056
rect 16574 13988 16580 14000
rect 10537 13960 16580 13988
rect 8076 13948 8082 13960
rect 16574 13948 16580 13960
rect 16632 13988 16638 14000
rect 21634 13988 21640 14000
rect 16632 13960 16988 13988
rect 21595 13960 21640 13988
rect 16632 13948 16638 13960
rect 5626 13920 5632 13932
rect 4096 13892 5632 13920
rect 4096 13861 4124 13892
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 7116 13920 7144 13948
rect 8297 13923 8355 13929
rect 8297 13920 8309 13923
rect 7116 13892 8309 13920
rect 8297 13889 8309 13892
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 10744 13892 11989 13920
rect 10744 13880 10750 13892
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 12952 13892 13185 13920
rect 12952 13880 12958 13892
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 13998 13920 14004 13932
rect 13173 13883 13231 13889
rect 13280 13892 14004 13920
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 4065 13855 4124 13861
rect 4065 13821 4077 13855
rect 4111 13821 4124 13855
rect 4177 13855 4235 13861
rect 4177 13854 4189 13855
rect 4172 13824 4189 13854
rect 4065 13815 4124 13821
rect 4177 13821 4189 13824
rect 4223 13854 4235 13855
rect 4223 13852 4292 13854
rect 4223 13826 4384 13852
rect 4223 13821 4235 13826
rect 4264 13824 4384 13826
rect 4177 13815 4235 13821
rect 4096 13784 4124 13815
rect 1452 13756 2544 13784
rect 3804 13756 4124 13784
rect 1452 13744 1458 13756
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 3804 13716 3832 13756
rect 2464 13688 3832 13716
rect 2464 13676 2470 13688
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 4062 13716 4068 13728
rect 3936 13688 4068 13716
rect 3936 13676 3942 13688
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4154 13676 4160 13728
rect 4212 13716 4218 13728
rect 4356 13716 4384 13824
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 5813 13855 5871 13861
rect 5813 13852 5825 13855
rect 5500 13824 5825 13852
rect 5500 13812 5506 13824
rect 5813 13821 5825 13824
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 6080 13855 6138 13861
rect 6080 13821 6092 13855
rect 6126 13852 6138 13855
rect 6454 13852 6460 13864
rect 6126 13824 6460 13852
rect 6126 13821 6138 13824
rect 6080 13815 6138 13821
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 6914 13852 6920 13864
rect 6696 13824 6920 13852
rect 6696 13812 6702 13824
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7558 13852 7564 13864
rect 7156 13824 7564 13852
rect 7156 13812 7162 13824
rect 7558 13812 7564 13824
rect 7616 13852 7622 13864
rect 7653 13855 7711 13861
rect 7653 13852 7665 13855
rect 7616 13824 7665 13852
rect 7616 13812 7622 13824
rect 7653 13821 7665 13824
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 8941 13855 8999 13861
rect 8941 13852 8953 13855
rect 8812 13824 8953 13852
rect 8812 13812 8818 13824
rect 8941 13821 8953 13824
rect 8987 13821 8999 13855
rect 9582 13852 9588 13864
rect 9543 13824 9588 13852
rect 8941 13815 8999 13821
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 9784 13824 11008 13852
rect 4798 13744 4804 13796
rect 4856 13784 4862 13796
rect 5074 13784 5080 13796
rect 4856 13756 5080 13784
rect 4856 13744 4862 13756
rect 5074 13744 5080 13756
rect 5132 13744 5138 13796
rect 5258 13784 5264 13796
rect 5219 13756 5264 13784
rect 5258 13744 5264 13756
rect 5316 13744 5322 13796
rect 8662 13744 8668 13796
rect 8720 13784 8726 13796
rect 9784 13784 9812 13824
rect 9858 13793 9864 13796
rect 8720 13756 9812 13784
rect 8720 13744 8726 13756
rect 9852 13747 9864 13793
rect 9916 13784 9922 13796
rect 10980 13784 11008 13824
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 11112 13824 12817 13852
rect 11112 13812 11118 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12986 13852 12992 13864
rect 12947 13824 12992 13852
rect 12805 13815 12863 13821
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13280 13852 13308 13892
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 14642 13880 14648 13932
rect 14700 13920 14706 13932
rect 15102 13920 15108 13932
rect 14700 13892 15108 13920
rect 14700 13880 14706 13892
rect 15102 13880 15108 13892
rect 15160 13920 15166 13932
rect 15381 13923 15439 13929
rect 15381 13920 15393 13923
rect 15160 13892 15393 13920
rect 15160 13880 15166 13892
rect 15381 13889 15393 13892
rect 15427 13889 15439 13923
rect 16390 13920 16396 13932
rect 15381 13883 15439 13889
rect 15589 13892 16396 13920
rect 13127 13824 13308 13852
rect 13357 13855 13415 13861
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 14090 13852 14096 13864
rect 13403 13824 14096 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15589 13852 15617 13892
rect 16390 13880 16396 13892
rect 16448 13920 16454 13932
rect 16666 13920 16672 13932
rect 16448 13892 16672 13920
rect 16448 13880 16454 13892
rect 15252 13824 15617 13852
rect 15657 13855 15715 13861
rect 15252 13812 15258 13824
rect 15657 13821 15669 13855
rect 15703 13852 15715 13855
rect 15746 13852 15752 13864
rect 15703 13824 15752 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 16592 13863 16620 13892
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 16850 13920 16856 13932
rect 16811 13892 16856 13920
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 16960 13929 16988 13960
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 22094 13948 22100 14000
rect 22152 13988 22158 14000
rect 24596 13988 24624 14028
rect 25682 14016 25688 14028
rect 25740 14016 25746 14068
rect 27154 14056 27160 14068
rect 25792 14028 26740 14056
rect 27115 14028 27160 14056
rect 24762 13988 24768 14000
rect 22152 13960 24624 13988
rect 24688 13960 24768 13988
rect 22152 13948 22158 13960
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13889 17003 13923
rect 16945 13883 17003 13889
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13920 18291 13923
rect 18322 13920 18328 13932
rect 18279 13892 18328 13920
rect 18279 13889 18291 13892
rect 18233 13883 18291 13889
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 19518 13920 19524 13932
rect 19479 13892 19524 13920
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 24688 13929 24716 13960
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 24854 13948 24860 14000
rect 24912 13988 24918 14000
rect 25792 13988 25820 14028
rect 24912 13960 25820 13988
rect 26712 13988 26740 14028
rect 27154 14016 27160 14028
rect 27212 14016 27218 14068
rect 27522 14016 27528 14068
rect 27580 14056 27586 14068
rect 29549 14059 29607 14065
rect 29549 14056 29561 14059
rect 27580 14028 29561 14056
rect 27580 14016 27586 14028
rect 29549 14025 29561 14028
rect 29595 14025 29607 14059
rect 30742 14056 30748 14068
rect 30703 14028 30748 14056
rect 29549 14019 29607 14025
rect 30742 14016 30748 14028
rect 30800 14016 30806 14068
rect 28534 13988 28540 14000
rect 26712 13960 28540 13988
rect 24912 13948 24918 13960
rect 28534 13948 28540 13960
rect 28592 13948 28598 14000
rect 29822 13948 29828 14000
rect 29880 13988 29886 14000
rect 30190 13988 30196 14000
rect 29880 13960 30196 13988
rect 29880 13948 29886 13960
rect 30190 13948 30196 13960
rect 30248 13988 30254 14000
rect 30834 13988 30840 14000
rect 30248 13960 30840 13988
rect 30248 13948 30254 13960
rect 30834 13948 30840 13960
rect 30892 13948 30898 14000
rect 21729 13923 21787 13929
rect 21729 13920 21741 13923
rect 20548 13892 21741 13920
rect 16577 13857 16635 13863
rect 16577 13823 16589 13857
rect 16623 13823 16635 13857
rect 17129 13855 17187 13861
rect 16749 13849 16807 13855
rect 17129 13852 17141 13855
rect 16749 13846 16761 13849
rect 16577 13817 16635 13823
rect 16684 13818 16761 13846
rect 13262 13784 13268 13796
rect 9916 13756 9952 13784
rect 10980 13756 13268 13784
rect 9858 13744 9864 13747
rect 9916 13744 9922 13756
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 14185 13787 14243 13793
rect 14185 13753 14197 13787
rect 14231 13784 14243 13787
rect 14642 13784 14648 13796
rect 14231 13756 14648 13784
rect 14231 13753 14243 13756
rect 14185 13747 14243 13753
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 16482 13744 16488 13796
rect 16540 13784 16546 13796
rect 16684 13784 16712 13818
rect 16749 13815 16761 13818
rect 16795 13815 16807 13849
rect 16749 13809 16807 13815
rect 17127 13821 17141 13852
rect 17175 13821 17187 13855
rect 17127 13815 17187 13821
rect 17313 13855 17371 13861
rect 17313 13821 17325 13855
rect 17359 13852 17371 13855
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17359 13824 17785 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 17773 13821 17785 13824
rect 17819 13821 17831 13855
rect 17954 13852 17960 13864
rect 17915 13824 17960 13852
rect 17773 13815 17831 13821
rect 16540 13756 16712 13784
rect 17127 13784 17155 13815
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 18046 13812 18052 13864
rect 18104 13852 18110 13864
rect 20548 13852 20576 13892
rect 21729 13889 21741 13892
rect 21775 13889 21787 13923
rect 24673 13923 24731 13929
rect 21729 13883 21787 13889
rect 22664 13892 24624 13920
rect 22664 13864 22692 13892
rect 18104 13824 20576 13852
rect 21545 13855 21603 13861
rect 18104 13812 18110 13824
rect 21545 13821 21557 13855
rect 21591 13821 21603 13855
rect 21818 13852 21824 13864
rect 21779 13824 21824 13852
rect 21545 13815 21603 13821
rect 17218 13784 17224 13796
rect 17127 13756 17224 13784
rect 16540 13744 16546 13756
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 18325 13787 18383 13793
rect 18325 13753 18337 13787
rect 18371 13784 18383 13787
rect 18414 13784 18420 13796
rect 18371 13756 18420 13784
rect 18371 13753 18383 13756
rect 18325 13747 18383 13753
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 19788 13787 19846 13793
rect 19788 13753 19800 13787
rect 19834 13784 19846 13787
rect 19978 13784 19984 13796
rect 19834 13756 19984 13784
rect 19834 13753 19846 13756
rect 19788 13747 19846 13753
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 21450 13744 21456 13796
rect 21508 13784 21514 13796
rect 21560 13784 21588 13815
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13852 22063 13855
rect 22465 13855 22523 13861
rect 22465 13852 22477 13855
rect 22051 13824 22477 13852
rect 22051 13821 22063 13824
rect 22005 13815 22063 13821
rect 22465 13821 22477 13824
rect 22511 13821 22523 13855
rect 22646 13852 22652 13864
rect 22607 13824 22652 13852
rect 22465 13815 22523 13821
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 22830 13852 22836 13864
rect 22791 13824 22836 13852
rect 22830 13812 22836 13824
rect 22888 13812 22894 13864
rect 22922 13812 22928 13864
rect 22980 13852 22986 13864
rect 22980 13824 23025 13852
rect 22980 13812 22986 13824
rect 23106 13812 23112 13864
rect 23164 13852 23170 13864
rect 24596 13861 24624 13892
rect 24673 13889 24685 13923
rect 24719 13889 24731 13923
rect 25130 13920 25136 13932
rect 24673 13883 24731 13889
rect 24780 13892 25136 13920
rect 24780 13861 24808 13892
rect 25130 13880 25136 13892
rect 25188 13880 25194 13932
rect 28994 13920 29000 13932
rect 28092 13892 29000 13920
rect 23569 13855 23627 13861
rect 23569 13852 23581 13855
rect 23164 13824 23581 13852
rect 23164 13812 23170 13824
rect 23569 13821 23581 13824
rect 23615 13821 23627 13855
rect 23569 13815 23627 13821
rect 24397 13855 24455 13861
rect 24397 13821 24409 13855
rect 24443 13852 24455 13855
rect 24581 13855 24639 13861
rect 24443 13824 24532 13852
rect 24443 13821 24455 13824
rect 24397 13815 24455 13821
rect 22554 13784 22560 13796
rect 21508 13756 22560 13784
rect 21508 13744 21514 13756
rect 22554 13744 22560 13756
rect 22612 13744 22618 13796
rect 24504 13784 24532 13824
rect 24581 13821 24593 13855
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 24765 13855 24823 13861
rect 24765 13821 24777 13855
rect 24811 13821 24823 13855
rect 24946 13852 24952 13864
rect 24907 13824 24952 13852
rect 24765 13815 24823 13821
rect 24946 13812 24952 13824
rect 25004 13812 25010 13864
rect 25590 13852 25596 13864
rect 25056 13824 25596 13852
rect 25056 13784 25084 13824
rect 25590 13812 25596 13824
rect 25648 13812 25654 13864
rect 25777 13855 25835 13861
rect 25777 13821 25789 13855
rect 25823 13852 25835 13855
rect 25866 13852 25872 13864
rect 25823 13824 25872 13852
rect 25823 13821 25835 13824
rect 25777 13815 25835 13821
rect 25866 13812 25872 13824
rect 25924 13812 25930 13864
rect 26044 13855 26102 13861
rect 26044 13821 26056 13855
rect 26090 13852 26102 13855
rect 26418 13852 26424 13864
rect 26090 13824 26424 13852
rect 26090 13821 26102 13824
rect 26044 13815 26102 13821
rect 26418 13812 26424 13824
rect 26476 13812 26482 13864
rect 28092 13861 28120 13892
rect 28994 13880 29000 13892
rect 29052 13880 29058 13932
rect 30926 13880 30932 13932
rect 30984 13920 30990 13932
rect 31021 13923 31079 13929
rect 31021 13920 31033 13923
rect 30984 13892 31033 13920
rect 30984 13880 30990 13892
rect 31021 13889 31033 13892
rect 31067 13889 31079 13923
rect 31021 13883 31079 13889
rect 28077 13855 28135 13861
rect 28077 13821 28089 13855
rect 28123 13821 28135 13855
rect 28077 13815 28135 13821
rect 28166 13812 28172 13864
rect 28224 13852 28230 13864
rect 28261 13855 28319 13861
rect 28261 13852 28273 13855
rect 28224 13824 28273 13852
rect 28224 13812 28230 13824
rect 28261 13821 28273 13824
rect 28307 13821 28319 13855
rect 28261 13815 28319 13821
rect 28353 13855 28411 13861
rect 28353 13821 28365 13855
rect 28399 13821 28411 13855
rect 28353 13815 28411 13821
rect 24504 13756 25084 13784
rect 27246 13744 27252 13796
rect 27304 13784 27310 13796
rect 28368 13784 28396 13815
rect 28442 13812 28448 13864
rect 28500 13852 28506 13864
rect 28629 13855 28687 13861
rect 28500 13824 28545 13852
rect 28500 13812 28506 13824
rect 28629 13821 28641 13855
rect 28675 13852 28687 13855
rect 28718 13852 28724 13864
rect 28675 13824 28724 13852
rect 28675 13821 28687 13824
rect 28629 13815 28687 13821
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 30101 13855 30159 13861
rect 30101 13821 30113 13855
rect 30147 13852 30159 13855
rect 30374 13852 30380 13864
rect 30147 13824 30380 13852
rect 30147 13821 30159 13824
rect 30101 13815 30159 13821
rect 30374 13812 30380 13824
rect 30432 13812 30438 13864
rect 30466 13812 30472 13864
rect 30524 13852 30530 13864
rect 30650 13852 30656 13864
rect 30524 13824 30656 13852
rect 30524 13812 30530 13824
rect 30650 13812 30656 13824
rect 30708 13852 30714 13864
rect 30745 13855 30803 13861
rect 30745 13852 30757 13855
rect 30708 13824 30757 13852
rect 30708 13812 30714 13824
rect 30745 13821 30757 13824
rect 30791 13821 30803 13855
rect 30745 13815 30803 13821
rect 27304 13756 28396 13784
rect 30300 13756 30972 13784
rect 27304 13744 27310 13756
rect 4212 13688 4384 13716
rect 5169 13719 5227 13725
rect 4212 13676 4218 13688
rect 5169 13685 5181 13719
rect 5215 13716 5227 13719
rect 5994 13716 6000 13728
rect 5215 13688 6000 13716
rect 5215 13685 5227 13688
rect 5169 13679 5227 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 10410 13716 10416 13728
rect 10008 13688 10416 13716
rect 10008 13676 10014 13688
rect 10410 13676 10416 13688
rect 10468 13716 10474 13728
rect 10965 13719 11023 13725
rect 10965 13716 10977 13719
rect 10468 13688 10977 13716
rect 10468 13676 10474 13688
rect 10965 13685 10977 13688
rect 11011 13685 11023 13719
rect 10965 13679 11023 13685
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13446 13716 13452 13728
rect 12768 13688 13452 13716
rect 12768 13676 12774 13688
rect 13446 13676 13452 13688
rect 13504 13716 13510 13728
rect 18230 13716 18236 13728
rect 13504 13688 18236 13716
rect 13504 13676 13510 13688
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 20530 13676 20536 13728
rect 20588 13716 20594 13728
rect 24762 13716 24768 13728
rect 20588 13688 24768 13716
rect 20588 13676 20594 13688
rect 24762 13676 24768 13688
rect 24820 13676 24826 13728
rect 25130 13716 25136 13728
rect 25091 13688 25136 13716
rect 25130 13676 25136 13688
rect 25188 13676 25194 13728
rect 25682 13676 25688 13728
rect 25740 13716 25746 13728
rect 27430 13716 27436 13728
rect 25740 13688 27436 13716
rect 25740 13676 25746 13688
rect 27430 13676 27436 13688
rect 27488 13676 27494 13728
rect 27890 13716 27896 13728
rect 27851 13688 27896 13716
rect 27890 13676 27896 13688
rect 27948 13676 27954 13728
rect 30300 13725 30328 13756
rect 30285 13719 30343 13725
rect 30285 13685 30297 13719
rect 30331 13685 30343 13719
rect 30944 13716 30972 13756
rect 30944 13688 32352 13716
rect 30285 13679 30343 13685
rect 1104 13626 32016 13648
rect 1104 13574 11253 13626
rect 11305 13574 11317 13626
rect 11369 13574 11381 13626
rect 11433 13574 11445 13626
rect 11497 13574 11509 13626
rect 11561 13574 21557 13626
rect 21609 13574 21621 13626
rect 21673 13574 21685 13626
rect 21737 13574 21749 13626
rect 21801 13574 21813 13626
rect 21865 13574 32016 13626
rect 1104 13552 32016 13574
rect 1394 13512 1400 13524
rect 1355 13484 1400 13512
rect 1394 13472 1400 13484
rect 1452 13512 1458 13524
rect 4062 13512 4068 13524
rect 1452 13484 4068 13512
rect 1452 13472 1458 13484
rect 1670 13404 1676 13456
rect 1728 13444 1734 13456
rect 2406 13444 2412 13456
rect 1728 13416 2412 13444
rect 1728 13404 1734 13416
rect 2406 13404 2412 13416
rect 2464 13404 2470 13456
rect 2532 13447 2590 13453
rect 2532 13413 2544 13447
rect 2578 13444 2590 13447
rect 3237 13447 3295 13453
rect 3237 13444 3249 13447
rect 2578 13416 3249 13444
rect 2578 13413 2590 13416
rect 2532 13407 2590 13413
rect 3237 13413 3249 13416
rect 3283 13413 3295 13447
rect 3237 13407 3295 13413
rect 2682 13336 2688 13388
rect 2740 13376 2746 13388
rect 3436 13385 3464 13484
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 4304 13484 5181 13512
rect 4304 13472 4310 13484
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 5258 13472 5264 13524
rect 5316 13512 5322 13524
rect 5718 13512 5724 13524
rect 5316 13484 5724 13512
rect 5316 13472 5322 13484
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 5868 13484 5913 13512
rect 5868 13472 5874 13484
rect 7742 13472 7748 13524
rect 7800 13512 7806 13524
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 7800 13484 7849 13512
rect 7800 13472 7806 13484
rect 7837 13481 7849 13484
rect 7883 13481 7895 13515
rect 7837 13475 7895 13481
rect 9769 13515 9827 13521
rect 9769 13481 9781 13515
rect 9815 13512 9827 13515
rect 9858 13512 9864 13524
rect 9815 13484 9864 13512
rect 9815 13481 9827 13484
rect 9769 13475 9827 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10318 13472 10324 13524
rect 10376 13472 10382 13524
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13906 13512 13912 13524
rect 13587 13484 13912 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 14737 13515 14795 13521
rect 14737 13481 14749 13515
rect 14783 13512 14795 13515
rect 15470 13512 15476 13524
rect 14783 13484 15476 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 17865 13515 17923 13521
rect 16632 13484 17724 13512
rect 16632 13472 16638 13484
rect 3878 13444 3884 13456
rect 3804 13416 3884 13444
rect 3804 13385 3832 13416
rect 3878 13404 3884 13416
rect 3936 13404 3942 13456
rect 4080 13444 4108 13472
rect 6638 13444 6644 13456
rect 4080 13416 5120 13444
rect 6551 13416 6644 13444
rect 3985 13389 4043 13395
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2740 13348 2789 13376
rect 2740 13336 2746 13348
rect 2777 13345 2789 13348
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13345 3479 13379
rect 3421 13339 3479 13345
rect 3789 13379 3847 13385
rect 3789 13345 3801 13379
rect 3835 13345 3847 13379
rect 3985 13376 3997 13389
rect 3789 13339 3847 13345
rect 3896 13355 3997 13376
rect 4031 13355 4043 13389
rect 5092 13388 5120 13416
rect 3896 13349 4043 13355
rect 3896 13348 4016 13349
rect 0 13308 800 13322
rect 3896 13320 3924 13348
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4617 13379 4675 13385
rect 4617 13376 4629 13379
rect 4304 13348 4629 13376
rect 4304 13336 4310 13348
rect 4617 13345 4629 13348
rect 4663 13345 4675 13379
rect 5074 13376 5080 13388
rect 4987 13348 5080 13376
rect 4617 13339 4675 13345
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 6564 13385 6592 13416
rect 6638 13404 6644 13416
rect 6696 13444 6702 13456
rect 6822 13444 6828 13456
rect 6696 13416 6828 13444
rect 6696 13404 6702 13416
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 8757 13447 8815 13453
rect 8757 13413 8769 13447
rect 8803 13444 8815 13447
rect 9309 13447 9367 13453
rect 9309 13444 9321 13447
rect 8803 13416 9321 13444
rect 8803 13413 8815 13416
rect 8757 13407 8815 13413
rect 9309 13413 9321 13416
rect 9355 13444 9367 13447
rect 10336 13444 10364 13472
rect 13449 13447 13507 13453
rect 9355 13416 10548 13444
rect 9355 13413 9367 13416
rect 9309 13407 9367 13413
rect 6549 13379 6607 13385
rect 6549 13345 6561 13379
rect 6595 13345 6607 13379
rect 6730 13376 6736 13388
rect 6691 13348 6736 13376
rect 6549 13339 6607 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7929 13379 7987 13385
rect 7156 13348 7201 13376
rect 7156 13336 7162 13348
rect 7929 13345 7941 13379
rect 7975 13376 7987 13379
rect 8110 13376 8116 13388
rect 7975 13348 8116 13376
rect 7975 13345 7987 13348
rect 7929 13339 7987 13345
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 9950 13376 9956 13388
rect 9911 13348 9956 13376
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10318 13376 10324 13388
rect 10279 13348 10324 13376
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 10520 13385 10548 13416
rect 13449 13413 13461 13447
rect 13495 13444 13507 13447
rect 14642 13444 14648 13456
rect 13495 13416 14648 13444
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 15654 13404 15660 13456
rect 15712 13444 15718 13456
rect 15850 13447 15908 13453
rect 15850 13444 15862 13447
rect 15712 13416 15862 13444
rect 15712 13404 15718 13416
rect 15850 13413 15862 13416
rect 15896 13413 15908 13447
rect 15850 13407 15908 13413
rect 15959 13416 16252 13444
rect 10505 13379 10563 13385
rect 10505 13345 10517 13379
rect 10551 13376 10563 13379
rect 10686 13376 10692 13388
rect 10551 13348 10692 13376
rect 10551 13345 10563 13348
rect 10505 13339 10563 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 11773 13379 11831 13385
rect 11773 13376 11785 13379
rect 11664 13348 11785 13376
rect 11664 13336 11670 13348
rect 11773 13345 11785 13348
rect 11819 13345 11831 13379
rect 11773 13339 11831 13345
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 13538 13376 13544 13388
rect 13136 13348 13544 13376
rect 13136 13336 13142 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 14277 13379 14335 13385
rect 14277 13345 14289 13379
rect 14323 13376 14335 13379
rect 14826 13376 14832 13388
rect 14323 13348 14832 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 1394 13308 1400 13320
rect 0 13280 1400 13308
rect 0 13266 800 13280
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3605 13311 3663 13317
rect 3605 13308 3617 13311
rect 3384 13280 3617 13308
rect 3384 13268 3390 13280
rect 3605 13277 3617 13280
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 3697 13311 3755 13317
rect 3697 13277 3709 13311
rect 3743 13277 3755 13311
rect 3697 13271 3755 13277
rect 3712 13240 3740 13271
rect 3878 13268 3884 13320
rect 3936 13268 3942 13320
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5166 13308 5172 13320
rect 4764 13280 5172 13308
rect 4764 13268 4770 13280
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6564 13280 6837 13308
rect 6564 13252 6592 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 10137 13311 10195 13317
rect 6972 13280 7017 13308
rect 6972 13268 6978 13280
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13308 10287 13311
rect 10594 13308 10600 13320
rect 10275 13280 10600 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 3160 13212 3740 13240
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 2130 13172 2136 13184
rect 1912 13144 2136 13172
rect 1912 13132 1918 13144
rect 2130 13132 2136 13144
rect 2188 13172 2194 13184
rect 3160 13172 3188 13212
rect 4062 13200 4068 13252
rect 4120 13240 4126 13252
rect 5442 13240 5448 13252
rect 4120 13212 5448 13240
rect 4120 13200 4126 13212
rect 5442 13200 5448 13212
rect 5500 13200 5506 13252
rect 6546 13200 6552 13252
rect 6604 13200 6610 13252
rect 10152 13240 10180 13271
rect 10594 13268 10600 13280
rect 10652 13308 10658 13320
rect 11054 13308 11060 13320
rect 10652 13280 11060 13308
rect 10652 13268 10658 13280
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 11146 13240 11152 13252
rect 10152 13212 11152 13240
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 4522 13172 4528 13184
rect 2188 13144 3188 13172
rect 4483 13144 4528 13172
rect 2188 13132 2194 13144
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 5166 13132 5172 13184
rect 5224 13172 5230 13184
rect 5350 13172 5356 13184
rect 5224 13144 5356 13172
rect 5224 13132 5230 13144
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5718 13132 5724 13184
rect 5776 13172 5782 13184
rect 5902 13172 5908 13184
rect 5776 13144 5908 13172
rect 5776 13132 5782 13144
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 7282 13172 7288 13184
rect 7243 13144 7288 13172
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 11532 13172 11560 13271
rect 12894 13240 12900 13252
rect 12807 13212 12900 13240
rect 12894 13200 12900 13212
rect 12952 13240 12958 13252
rect 14292 13240 14320 13339
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15959 13376 15987 13416
rect 16114 13376 16120 13388
rect 15344 13348 15987 13376
rect 16075 13348 16120 13376
rect 15344 13336 15350 13348
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 16224 13308 16252 13416
rect 16482 13404 16488 13456
rect 16540 13444 16546 13456
rect 16942 13444 16948 13456
rect 16540 13416 16948 13444
rect 16540 13404 16546 13416
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 17586 13444 17592 13456
rect 17144 13416 17592 13444
rect 16390 13336 16396 13388
rect 16448 13376 16454 13388
rect 17144 13385 17172 13416
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 16448 13348 16865 13376
rect 16448 13336 16454 13348
rect 16853 13345 16865 13348
rect 16899 13345 16911 13379
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 16853 13339 16911 13345
rect 16951 13348 17049 13376
rect 16951 13308 16979 13348
rect 17037 13345 17049 13348
rect 17083 13345 17095 13379
rect 17037 13339 17095 13345
rect 17126 13379 17184 13385
rect 17126 13345 17138 13379
rect 17172 13345 17184 13379
rect 17126 13339 17184 13345
rect 17230 13336 17236 13388
rect 17288 13378 17294 13388
rect 17405 13379 17463 13385
rect 17288 13350 17331 13378
rect 17288 13336 17294 13350
rect 17405 13345 17417 13379
rect 17451 13345 17463 13379
rect 17696 13376 17724 13484
rect 17865 13481 17877 13515
rect 17911 13512 17923 13515
rect 18138 13512 18144 13524
rect 17911 13484 18144 13512
rect 17911 13481 17923 13484
rect 17865 13475 17923 13481
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 19610 13472 19616 13524
rect 19668 13512 19674 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 19668 13484 20269 13512
rect 19668 13472 19674 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 20257 13475 20315 13481
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 22278 13512 22284 13524
rect 21232 13484 22284 13512
rect 21232 13472 21238 13484
rect 21836 13456 21864 13484
rect 22278 13472 22284 13484
rect 22336 13512 22342 13524
rect 22389 13515 22447 13521
rect 22389 13512 22401 13515
rect 22336 13484 22401 13512
rect 22336 13472 22342 13484
rect 22389 13481 22401 13484
rect 22435 13481 22447 13515
rect 22389 13475 22447 13481
rect 22557 13515 22615 13521
rect 22557 13481 22569 13515
rect 22603 13512 22615 13515
rect 23106 13512 23112 13524
rect 22603 13484 23112 13512
rect 22603 13481 22615 13484
rect 22557 13475 22615 13481
rect 23106 13472 23112 13484
rect 23164 13472 23170 13524
rect 23569 13515 23627 13521
rect 23569 13481 23581 13515
rect 23615 13512 23627 13515
rect 23750 13512 23756 13524
rect 23615 13484 23756 13512
rect 23615 13481 23627 13484
rect 23569 13475 23627 13481
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 18978 13447 19036 13453
rect 18978 13444 18990 13447
rect 18840 13416 18990 13444
rect 18840 13404 18846 13416
rect 18978 13413 18990 13416
rect 19024 13413 19036 13447
rect 20162 13444 20168 13456
rect 18978 13407 19036 13413
rect 19076 13416 20168 13444
rect 19076 13376 19104 13416
rect 20162 13404 20168 13416
rect 20220 13404 20226 13456
rect 21358 13404 21364 13456
rect 21416 13444 21422 13456
rect 21542 13444 21548 13456
rect 21416 13416 21548 13444
rect 21416 13404 21422 13416
rect 21542 13404 21548 13416
rect 21600 13404 21606 13456
rect 21818 13404 21824 13456
rect 21876 13404 21882 13456
rect 22189 13447 22247 13453
rect 22189 13413 22201 13447
rect 22235 13444 22247 13447
rect 22235 13416 22416 13444
rect 22235 13413 22247 13416
rect 22189 13407 22247 13413
rect 22388 13388 22416 13416
rect 17696 13348 19104 13376
rect 19245 13379 19303 13385
rect 17405 13339 17463 13345
rect 19245 13345 19257 13379
rect 19291 13376 19303 13379
rect 19518 13376 19524 13388
rect 19291 13348 19524 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 17420 13308 17448 13339
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 19702 13336 19708 13388
rect 19760 13336 19766 13388
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 22094 13376 22100 13388
rect 20772 13348 22100 13376
rect 20772 13336 20778 13348
rect 22094 13336 22100 13348
rect 22152 13336 22158 13388
rect 22370 13336 22376 13388
rect 22428 13336 22434 13388
rect 16224 13280 16979 13308
rect 17328 13280 17448 13308
rect 19720 13308 19748 13336
rect 22462 13308 22468 13320
rect 19720 13280 22468 13308
rect 12952 13212 14320 13240
rect 12952 13200 12958 13212
rect 16114 13200 16120 13252
rect 16172 13240 16178 13252
rect 16390 13240 16396 13252
rect 16172 13212 16396 13240
rect 16172 13200 16178 13212
rect 16390 13200 16396 13212
rect 16448 13200 16454 13252
rect 17328 13240 17356 13280
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 16592 13212 17356 13240
rect 11882 13172 11888 13184
rect 11532 13144 11888 13172
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 14182 13172 14188 13184
rect 14143 13144 14188 13172
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 15102 13132 15108 13184
rect 15160 13172 15166 13184
rect 16592 13172 16620 13212
rect 17402 13200 17408 13252
rect 17460 13240 17466 13252
rect 18046 13240 18052 13252
rect 17460 13212 18052 13240
rect 17460 13200 17466 13212
rect 18046 13200 18052 13212
rect 18104 13200 18110 13252
rect 19334 13200 19340 13252
rect 19392 13240 19398 13252
rect 19705 13243 19763 13249
rect 19705 13240 19717 13243
rect 19392 13212 19717 13240
rect 19392 13200 19398 13212
rect 19705 13209 19717 13212
rect 19751 13240 19763 13243
rect 23584 13240 23612 13475
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 24029 13515 24087 13521
rect 24029 13481 24041 13515
rect 24075 13512 24087 13515
rect 24946 13512 24952 13524
rect 24075 13484 24952 13512
rect 24075 13481 24087 13484
rect 24029 13475 24087 13481
rect 24946 13472 24952 13484
rect 25004 13512 25010 13524
rect 25004 13484 25912 13512
rect 25004 13472 25010 13484
rect 23658 13404 23664 13456
rect 23716 13444 23722 13456
rect 23716 13416 25452 13444
rect 23716 13404 23722 13416
rect 25130 13336 25136 13388
rect 25188 13385 25194 13388
rect 25424 13385 25452 13416
rect 25884 13385 25912 13484
rect 30374 13472 30380 13524
rect 30432 13512 30438 13524
rect 30558 13512 30564 13524
rect 30432 13484 30564 13512
rect 30432 13472 30438 13484
rect 30558 13472 30564 13484
rect 30616 13472 30622 13524
rect 25958 13404 25964 13456
rect 26016 13444 26022 13456
rect 26016 13416 27292 13444
rect 26016 13404 26022 13416
rect 25188 13376 25200 13385
rect 25409 13379 25467 13385
rect 25188 13348 25233 13376
rect 25188 13339 25200 13348
rect 25409 13345 25421 13379
rect 25455 13345 25467 13379
rect 25409 13339 25467 13345
rect 25869 13379 25927 13385
rect 25869 13345 25881 13379
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 25188 13336 25194 13339
rect 27062 13336 27068 13388
rect 27120 13376 27126 13388
rect 27264 13385 27292 13416
rect 29178 13404 29184 13456
rect 29236 13444 29242 13456
rect 29466 13447 29524 13453
rect 29466 13444 29478 13447
rect 29236 13416 29478 13444
rect 29236 13404 29242 13416
rect 29466 13413 29478 13416
rect 29512 13413 29524 13447
rect 32324 13444 32352 13688
rect 29466 13407 29524 13413
rect 29564 13416 30604 13444
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 27120 13348 27169 13376
rect 27120 13336 27126 13348
rect 27157 13345 27169 13348
rect 27203 13345 27215 13379
rect 27157 13339 27215 13345
rect 27249 13379 27307 13385
rect 27249 13345 27261 13379
rect 27295 13376 27307 13379
rect 29564 13376 29592 13416
rect 29730 13376 29736 13388
rect 27295 13348 29592 13376
rect 29691 13348 29736 13376
rect 27295 13345 27307 13348
rect 27249 13339 27307 13345
rect 29730 13336 29736 13348
rect 29788 13336 29794 13388
rect 30576 13385 30604 13416
rect 32232 13416 32352 13444
rect 30561 13379 30619 13385
rect 30561 13345 30573 13379
rect 30607 13376 30619 13379
rect 31202 13376 31208 13388
rect 30607 13348 31208 13376
rect 30607 13345 30619 13348
rect 30561 13339 30619 13345
rect 31202 13336 31208 13348
rect 31260 13336 31266 13388
rect 26602 13268 26608 13320
rect 26660 13308 26666 13320
rect 26973 13311 27031 13317
rect 26973 13308 26985 13311
rect 26660 13280 26985 13308
rect 26660 13268 26666 13280
rect 26973 13277 26985 13280
rect 27019 13277 27031 13311
rect 30834 13308 30840 13320
rect 30795 13280 30840 13308
rect 26973 13271 27031 13277
rect 30834 13268 30840 13280
rect 30892 13268 30898 13320
rect 32232 13308 32260 13416
rect 32320 13308 33120 13322
rect 32232 13280 33120 13308
rect 32320 13266 33120 13280
rect 27709 13243 27767 13249
rect 27709 13240 27721 13243
rect 19751 13212 23612 13240
rect 25801 13212 27721 13240
rect 19751 13209 19763 13212
rect 19705 13203 19763 13209
rect 15160 13144 16620 13172
rect 16669 13175 16727 13181
rect 15160 13132 15166 13144
rect 16669 13141 16681 13175
rect 16715 13172 16727 13175
rect 16758 13172 16764 13184
rect 16715 13144 16764 13172
rect 16715 13141 16727 13144
rect 16669 13135 16727 13141
rect 16758 13132 16764 13144
rect 16816 13132 16822 13184
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 20714 13172 20720 13184
rect 18196 13144 20720 13172
rect 18196 13132 18202 13144
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 21269 13175 21327 13181
rect 21269 13141 21281 13175
rect 21315 13172 21327 13175
rect 21450 13172 21456 13184
rect 21315 13144 21456 13172
rect 21315 13141 21327 13144
rect 21269 13135 21327 13141
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 21542 13132 21548 13184
rect 21600 13172 21606 13184
rect 22278 13172 22284 13184
rect 21600 13144 22284 13172
rect 21600 13132 21606 13144
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 22373 13175 22431 13181
rect 22373 13141 22385 13175
rect 22419 13172 22431 13175
rect 22922 13172 22928 13184
rect 22419 13144 22928 13172
rect 22419 13141 22431 13144
rect 22373 13135 22431 13141
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 24762 13132 24768 13184
rect 24820 13172 24826 13184
rect 25801 13172 25829 13212
rect 27709 13209 27721 13212
rect 27755 13240 27767 13243
rect 27755 13212 28856 13240
rect 27755 13209 27767 13212
rect 27709 13203 27767 13209
rect 25958 13172 25964 13184
rect 24820 13144 25829 13172
rect 25919 13144 25964 13172
rect 24820 13132 24826 13144
rect 25958 13132 25964 13144
rect 26016 13132 26022 13184
rect 27062 13172 27068 13184
rect 27023 13144 27068 13172
rect 27062 13132 27068 13144
rect 27120 13132 27126 13184
rect 28353 13175 28411 13181
rect 28353 13141 28365 13175
rect 28399 13172 28411 13175
rect 28442 13172 28448 13184
rect 28399 13144 28448 13172
rect 28399 13141 28411 13144
rect 28353 13135 28411 13141
rect 28442 13132 28448 13144
rect 28500 13132 28506 13184
rect 28828 13172 28856 13212
rect 30282 13200 30288 13252
rect 30340 13240 30346 13252
rect 30653 13243 30711 13249
rect 30653 13240 30665 13243
rect 30340 13212 30665 13240
rect 30340 13200 30346 13212
rect 30653 13209 30665 13212
rect 30699 13209 30711 13243
rect 30653 13203 30711 13209
rect 30098 13172 30104 13184
rect 28828 13144 30104 13172
rect 30098 13132 30104 13144
rect 30156 13132 30162 13184
rect 30742 13172 30748 13184
rect 30703 13144 30748 13172
rect 30742 13132 30748 13144
rect 30800 13132 30806 13184
rect 1104 13082 32016 13104
rect 1104 13030 6102 13082
rect 6154 13030 6166 13082
rect 6218 13030 6230 13082
rect 6282 13030 6294 13082
rect 6346 13030 6358 13082
rect 6410 13030 16405 13082
rect 16457 13030 16469 13082
rect 16521 13030 16533 13082
rect 16585 13030 16597 13082
rect 16649 13030 16661 13082
rect 16713 13030 26709 13082
rect 26761 13030 26773 13082
rect 26825 13030 26837 13082
rect 26889 13030 26901 13082
rect 26953 13030 26965 13082
rect 27017 13030 32016 13082
rect 1104 13008 32016 13030
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3878 12968 3884 12980
rect 2832 12940 3884 12968
rect 2832 12928 2838 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4982 12928 4988 12980
rect 5040 12968 5046 12980
rect 5077 12971 5135 12977
rect 5077 12968 5089 12971
rect 5040 12940 5089 12968
rect 5040 12928 5046 12940
rect 5077 12937 5089 12940
rect 5123 12937 5135 12971
rect 5077 12931 5135 12937
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 6089 12971 6147 12977
rect 6089 12968 6101 12971
rect 5776 12940 6101 12968
rect 5776 12928 5782 12940
rect 6089 12937 6101 12940
rect 6135 12937 6147 12971
rect 10318 12968 10324 12980
rect 10279 12940 10324 12968
rect 6089 12931 6147 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11606 12968 11612 12980
rect 11563 12940 11612 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 15657 12971 15715 12977
rect 13280 12940 15617 12968
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3237 12903 3295 12909
rect 3237 12900 3249 12903
rect 2924 12872 3249 12900
rect 2924 12860 2930 12872
rect 3237 12869 3249 12872
rect 3283 12900 3295 12903
rect 4246 12900 4252 12912
rect 3283 12872 4252 12900
rect 3283 12869 3295 12872
rect 3237 12863 3295 12869
rect 4246 12860 4252 12872
rect 4304 12860 4310 12912
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 6972 12872 7052 12900
rect 6972 12860 6978 12872
rect 4264 12832 4292 12860
rect 4264 12804 4936 12832
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 2682 12764 2688 12776
rect 1903 12736 2688 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 2682 12724 2688 12736
rect 2740 12764 2746 12776
rect 4062 12764 4068 12776
rect 2740 12736 4068 12764
rect 2740 12724 2746 12736
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 4908 12773 4936 12804
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 5905 12835 5963 12841
rect 5905 12832 5917 12835
rect 5040 12804 5917 12832
rect 5040 12792 5046 12804
rect 5905 12801 5917 12804
rect 5951 12801 5963 12835
rect 5905 12795 5963 12801
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 7024 12841 7052 12872
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 13280 12909 13308 12940
rect 13265 12903 13323 12909
rect 13265 12900 13277 12903
rect 12584 12872 13277 12900
rect 12584 12860 12590 12872
rect 13265 12869 13277 12872
rect 13311 12869 13323 12903
rect 15286 12900 15292 12912
rect 13265 12863 13323 12869
rect 14660 12872 15292 12900
rect 7009 12835 7067 12841
rect 6604 12804 6960 12832
rect 6604 12792 6610 12804
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4304 12736 4445 12764
rect 4304 12724 4310 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 4893 12767 4951 12773
rect 4893 12733 4905 12767
rect 4939 12733 4951 12767
rect 5074 12764 5080 12776
rect 5035 12736 5080 12764
rect 4893 12727 4951 12733
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 6181 12767 6239 12773
rect 6181 12733 6193 12767
rect 6227 12764 6239 12767
rect 6454 12764 6460 12776
rect 6227 12736 6460 12764
rect 6227 12733 6239 12736
rect 6181 12727 6239 12733
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 6638 12764 6644 12776
rect 6599 12736 6644 12764
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 6932 12773 6960 12804
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 7009 12795 7067 12801
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 12894 12832 12900 12844
rect 11348 12804 12900 12832
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 6917 12727 6975 12733
rect 1946 12656 1952 12708
rect 2004 12696 2010 12708
rect 2102 12699 2160 12705
rect 2102 12696 2114 12699
rect 2004 12668 2114 12696
rect 2004 12656 2010 12668
rect 2102 12665 2114 12668
rect 2148 12665 2160 12699
rect 2102 12659 2160 12665
rect 2590 12656 2596 12708
rect 2648 12696 2654 12708
rect 3878 12696 3884 12708
rect 2648 12668 3884 12696
rect 2648 12656 2654 12668
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 4341 12699 4399 12705
rect 4341 12665 4353 12699
rect 4387 12696 4399 12699
rect 5534 12696 5540 12708
rect 4387 12668 5540 12696
rect 4387 12665 4399 12668
rect 4341 12659 4399 12665
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 5718 12656 5724 12708
rect 5776 12696 5782 12708
rect 6656 12696 6684 12724
rect 5776 12668 6684 12696
rect 6840 12696 6868 12727
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7834 12764 7840 12776
rect 7795 12736 7840 12764
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12764 8999 12767
rect 9582 12764 9588 12776
rect 8987 12736 9588 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 10781 12767 10839 12773
rect 10781 12764 10793 12767
rect 10744 12736 10793 12764
rect 10744 12724 10750 12736
rect 10781 12733 10793 12736
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10928 12736 10977 12764
rect 10928 12724 10934 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 7098 12696 7104 12708
rect 6840 12668 7104 12696
rect 5776 12656 5782 12668
rect 7098 12656 7104 12668
rect 7156 12696 7162 12708
rect 7650 12696 7656 12708
rect 7156 12668 7656 12696
rect 7156 12656 7162 12668
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 9208 12699 9266 12705
rect 9208 12665 9220 12699
rect 9254 12696 9266 12699
rect 10980 12696 11008 12727
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11348 12773 11376 12804
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 14660 12841 14688 12872
rect 15286 12860 15292 12872
rect 15344 12860 15350 12912
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12832 14795 12835
rect 15378 12832 15384 12844
rect 14783 12804 15384 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 11333 12767 11391 12773
rect 11112 12736 11157 12764
rect 11112 12724 11118 12736
rect 11333 12733 11345 12767
rect 11379 12733 11391 12767
rect 12342 12764 12348 12776
rect 12303 12736 12348 12764
rect 11333 12727 11391 12733
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12764 12679 12767
rect 14182 12764 14188 12776
rect 12667 12736 14188 12764
rect 12667 12733 12679 12736
rect 12621 12727 12679 12733
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14461 12767 14519 12773
rect 14461 12733 14473 12767
rect 14507 12733 14519 12767
rect 14461 12727 14519 12733
rect 12710 12696 12716 12708
rect 9254 12668 9628 12696
rect 10980 12668 12716 12696
rect 9254 12665 9266 12668
rect 9208 12659 9266 12665
rect 9600 12640 9628 12668
rect 12710 12656 12716 12668
rect 12768 12656 12774 12708
rect 13081 12699 13139 12705
rect 13081 12665 13093 12699
rect 13127 12696 13139 12699
rect 13262 12696 13268 12708
rect 13127 12668 13268 12696
rect 13127 12665 13139 12668
rect 13081 12659 13139 12665
rect 13262 12656 13268 12668
rect 13320 12656 13326 12708
rect 14476 12696 14504 12727
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 15013 12767 15071 12773
rect 14884 12736 14929 12764
rect 14884 12724 14890 12736
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 15102 12764 15108 12776
rect 15059 12736 15108 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15470 12696 15476 12708
rect 14476 12668 15476 12696
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 15589 12696 15617 12940
rect 15657 12937 15669 12971
rect 15703 12968 15715 12971
rect 16114 12968 16120 12980
rect 15703 12940 16120 12968
rect 15703 12937 15715 12940
rect 15657 12931 15715 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 17770 12968 17776 12980
rect 17052 12940 17776 12968
rect 17052 12841 17080 12940
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18046 12928 18052 12980
rect 18104 12968 18110 12980
rect 19978 12968 19984 12980
rect 18104 12940 19546 12968
rect 19939 12940 19984 12968
rect 18104 12928 18110 12940
rect 19518 12900 19546 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 21913 12971 21971 12977
rect 21913 12937 21925 12971
rect 21959 12937 21971 12971
rect 21913 12931 21971 12937
rect 22097 12971 22155 12977
rect 22097 12937 22109 12971
rect 22143 12968 22155 12971
rect 22738 12968 22744 12980
rect 22143 12940 22744 12968
rect 22143 12937 22155 12940
rect 22097 12931 22155 12937
rect 19518 12872 19748 12900
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 17037 12795 17095 12801
rect 17144 12804 17601 12832
rect 16758 12724 16764 12776
rect 16816 12773 16822 12776
rect 16816 12764 16828 12773
rect 16816 12736 16861 12764
rect 16816 12727 16828 12736
rect 16816 12724 16822 12727
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17144 12764 17172 12804
rect 17589 12801 17601 12804
rect 17635 12801 17647 12835
rect 19518 12832 19524 12844
rect 19479 12804 19524 12832
rect 17589 12795 17647 12801
rect 19518 12792 19524 12804
rect 19576 12792 19582 12844
rect 19720 12832 19748 12872
rect 20806 12860 20812 12912
rect 20864 12900 20870 12912
rect 21266 12900 21272 12912
rect 20864 12872 21272 12900
rect 20864 12860 20870 12872
rect 21266 12860 21272 12872
rect 21324 12860 21330 12912
rect 21928 12900 21956 12931
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 23658 12968 23664 12980
rect 23571 12940 23664 12968
rect 23658 12928 23664 12940
rect 23716 12968 23722 12980
rect 24210 12968 24216 12980
rect 23716 12940 24216 12968
rect 23716 12928 23722 12940
rect 24210 12928 24216 12940
rect 24268 12928 24274 12980
rect 28994 12968 29000 12980
rect 27632 12940 28580 12968
rect 28955 12940 29000 12968
rect 22554 12900 22560 12912
rect 21928 12872 22560 12900
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 27632 12900 27660 12940
rect 22848 12872 27660 12900
rect 28552 12900 28580 12940
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 30282 12928 30288 12980
rect 30340 12968 30346 12980
rect 31021 12971 31079 12977
rect 31021 12968 31033 12971
rect 30340 12940 31033 12968
rect 30340 12928 30346 12940
rect 31021 12937 31033 12940
rect 31067 12937 31079 12971
rect 31021 12931 31079 12937
rect 29086 12900 29092 12912
rect 28552 12872 29092 12900
rect 20717 12835 20775 12841
rect 20717 12832 20729 12835
rect 19720 12804 20729 12832
rect 20717 12801 20729 12804
rect 20763 12832 20775 12835
rect 22738 12832 22744 12844
rect 20763 12804 22744 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 17000 12736 17172 12764
rect 17000 12724 17006 12736
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 17402 12764 17408 12776
rect 17276 12736 17408 12764
rect 17276 12724 17282 12736
rect 17402 12724 17408 12736
rect 17460 12764 17466 12776
rect 17497 12767 17555 12773
rect 17497 12764 17509 12767
rect 17460 12736 17509 12764
rect 17460 12724 17466 12736
rect 17497 12733 17509 12736
rect 17543 12733 17555 12767
rect 18138 12764 18144 12776
rect 17497 12727 17555 12733
rect 17788 12736 18144 12764
rect 17788 12696 17816 12736
rect 18138 12724 18144 12736
rect 18196 12724 18202 12776
rect 19150 12724 19156 12776
rect 19208 12764 19214 12776
rect 19245 12767 19303 12773
rect 19245 12764 19257 12767
rect 19208 12736 19257 12764
rect 19208 12724 19214 12736
rect 19245 12733 19257 12736
rect 19291 12733 19303 12767
rect 19429 12767 19487 12773
rect 19429 12764 19441 12767
rect 19245 12727 19303 12733
rect 19352 12736 19441 12764
rect 15589 12668 17816 12696
rect 17954 12656 17960 12708
rect 18012 12696 18018 12708
rect 19352 12696 19380 12736
rect 19429 12733 19441 12736
rect 19475 12733 19487 12767
rect 19610 12764 19616 12776
rect 19571 12736 19616 12764
rect 19429 12727 19487 12733
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20806 12764 20812 12776
rect 19843 12736 20812 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 21910 12764 21916 12776
rect 21192 12736 21916 12764
rect 19702 12696 19708 12708
rect 18012 12668 19288 12696
rect 19352 12668 19708 12696
rect 18012 12656 18018 12668
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5132 12600 5917 12628
rect 5132 12588 5138 12600
rect 5905 12597 5917 12600
rect 5951 12597 5963 12631
rect 5905 12591 5963 12597
rect 7377 12631 7435 12637
rect 7377 12597 7389 12631
rect 7423 12628 7435 12631
rect 7466 12628 7472 12640
rect 7423 12600 7472 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 7926 12628 7932 12640
rect 7887 12600 7932 12628
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 9582 12588 9588 12640
rect 9640 12588 9646 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10318 12628 10324 12640
rect 9824 12600 10324 12628
rect 9824 12588 9830 12600
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 14277 12631 14335 12637
rect 14277 12597 14289 12631
rect 14323 12628 14335 12631
rect 14366 12628 14372 12640
rect 14323 12600 14372 12628
rect 14323 12597 14335 12600
rect 14277 12591 14335 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 18046 12628 18052 12640
rect 14700 12600 18052 12628
rect 14700 12588 14706 12600
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18230 12628 18236 12640
rect 18191 12600 18236 12628
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 19260 12628 19288 12668
rect 19702 12656 19708 12668
rect 19760 12656 19766 12708
rect 21192 12640 21220 12736
rect 21910 12724 21916 12736
rect 21968 12724 21974 12776
rect 22462 12724 22468 12776
rect 22520 12764 22526 12776
rect 22557 12767 22615 12773
rect 22557 12764 22569 12767
rect 22520 12736 22569 12764
rect 22520 12724 22526 12736
rect 22557 12733 22569 12736
rect 22603 12764 22615 12767
rect 22646 12764 22652 12776
rect 22603 12736 22652 12764
rect 22603 12733 22615 12736
rect 22557 12727 22615 12733
rect 22646 12724 22652 12736
rect 22704 12764 22710 12776
rect 22848 12764 22876 12872
rect 29086 12860 29092 12872
rect 29144 12860 29150 12912
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25130 12832 25136 12844
rect 25087 12804 25136 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25130 12792 25136 12804
rect 25188 12832 25194 12844
rect 25498 12832 25504 12844
rect 25188 12804 25504 12832
rect 25188 12792 25194 12804
rect 25498 12792 25504 12804
rect 25556 12792 25562 12844
rect 27246 12832 27252 12844
rect 26896 12804 27252 12832
rect 22704 12736 22876 12764
rect 23017 12767 23075 12773
rect 22704 12724 22710 12736
rect 23017 12733 23029 12767
rect 23063 12733 23075 12767
rect 24486 12764 24492 12776
rect 24447 12736 24492 12764
rect 23017 12727 23075 12733
rect 21729 12699 21787 12705
rect 21729 12665 21741 12699
rect 21775 12696 21787 12699
rect 22186 12696 22192 12708
rect 21775 12668 22192 12696
rect 21775 12665 21787 12668
rect 21729 12659 21787 12665
rect 22186 12656 22192 12668
rect 22244 12696 22250 12708
rect 22370 12696 22376 12708
rect 22244 12668 22376 12696
rect 22244 12656 22250 12668
rect 22370 12656 22376 12668
rect 22428 12656 22434 12708
rect 22922 12656 22928 12708
rect 22980 12696 22986 12708
rect 23032 12696 23060 12727
rect 24486 12724 24492 12736
rect 24544 12724 24550 12776
rect 25682 12724 25688 12776
rect 25740 12764 25746 12776
rect 26896 12773 26924 12804
rect 27246 12792 27252 12804
rect 27304 12792 27310 12844
rect 30006 12832 30012 12844
rect 29967 12804 30012 12832
rect 30006 12792 30012 12804
rect 30064 12792 30070 12844
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 25740 12736 25789 12764
rect 25740 12724 25746 12736
rect 25777 12733 25789 12736
rect 25823 12733 25835 12767
rect 25777 12727 25835 12733
rect 26881 12767 26939 12773
rect 26881 12733 26893 12767
rect 26927 12733 26939 12767
rect 27062 12764 27068 12776
rect 27023 12736 27068 12764
rect 26881 12727 26939 12733
rect 27062 12724 27068 12736
rect 27120 12724 27126 12776
rect 27157 12767 27215 12773
rect 27157 12733 27169 12767
rect 27203 12764 27215 12767
rect 27338 12764 27344 12776
rect 27203 12736 27344 12764
rect 27203 12733 27215 12736
rect 27157 12727 27215 12733
rect 27338 12724 27344 12736
rect 27396 12724 27402 12776
rect 27617 12767 27675 12773
rect 27617 12733 27629 12767
rect 27663 12764 27675 12767
rect 29546 12764 29552 12776
rect 27663 12736 29552 12764
rect 27663 12733 27675 12736
rect 27617 12727 27675 12733
rect 22980 12668 23060 12696
rect 22980 12656 22986 12668
rect 25406 12656 25412 12708
rect 25464 12696 25470 12708
rect 25866 12696 25872 12708
rect 25464 12668 25872 12696
rect 25464 12656 25470 12668
rect 25866 12656 25872 12668
rect 25924 12656 25930 12708
rect 26050 12656 26056 12708
rect 26108 12696 26114 12708
rect 27632 12696 27660 12727
rect 29546 12724 29552 12736
rect 29604 12724 29610 12776
rect 29638 12724 29644 12776
rect 29696 12764 29702 12776
rect 29825 12767 29883 12773
rect 29696 12736 29741 12764
rect 29696 12724 29702 12736
rect 29825 12733 29837 12767
rect 29871 12733 29883 12767
rect 29825 12727 29883 12733
rect 27890 12705 27896 12708
rect 27884 12696 27896 12705
rect 26108 12668 27660 12696
rect 27851 12668 27896 12696
rect 26108 12656 26114 12668
rect 27884 12659 27896 12668
rect 27890 12656 27896 12659
rect 27948 12656 27954 12708
rect 29840 12696 29868 12727
rect 29914 12724 29920 12776
rect 29972 12764 29978 12776
rect 30190 12764 30196 12776
rect 29972 12736 30017 12764
rect 30151 12736 30196 12764
rect 29972 12724 29978 12736
rect 30190 12724 30196 12736
rect 30248 12764 30254 12776
rect 30374 12764 30380 12776
rect 30248 12736 30380 12764
rect 30248 12724 30254 12736
rect 30374 12724 30380 12736
rect 30432 12724 30438 12776
rect 30834 12724 30840 12776
rect 30892 12724 30898 12776
rect 30852 12696 30880 12724
rect 31205 12699 31263 12705
rect 31205 12696 31217 12699
rect 29840 12668 31217 12696
rect 31205 12665 31217 12668
rect 31251 12665 31263 12699
rect 31205 12659 31263 12665
rect 20714 12628 20720 12640
rect 19260 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21174 12628 21180 12640
rect 21135 12600 21180 12628
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 21910 12588 21916 12640
rect 21968 12637 21974 12640
rect 21968 12631 21987 12637
rect 21975 12597 21987 12631
rect 21968 12591 21987 12597
rect 21968 12588 21974 12591
rect 25682 12588 25688 12640
rect 25740 12628 25746 12640
rect 25961 12631 26019 12637
rect 25961 12628 25973 12631
rect 25740 12600 25973 12628
rect 25740 12588 25746 12600
rect 25961 12597 25973 12600
rect 26007 12597 26019 12631
rect 25961 12591 26019 12597
rect 26697 12631 26755 12637
rect 26697 12597 26709 12631
rect 26743 12628 26755 12631
rect 27522 12628 27528 12640
rect 26743 12600 27528 12628
rect 26743 12597 26755 12600
rect 26697 12591 26755 12597
rect 27522 12588 27528 12600
rect 27580 12588 27586 12640
rect 30190 12588 30196 12640
rect 30248 12628 30254 12640
rect 30377 12631 30435 12637
rect 30377 12628 30389 12631
rect 30248 12600 30389 12628
rect 30248 12588 30254 12600
rect 30377 12597 30389 12600
rect 30423 12597 30435 12631
rect 30834 12628 30840 12640
rect 30795 12600 30840 12628
rect 30377 12591 30435 12597
rect 30834 12588 30840 12600
rect 30892 12588 30898 12640
rect 31018 12637 31024 12640
rect 30995 12631 31024 12637
rect 30995 12597 31007 12631
rect 30995 12591 31024 12597
rect 31018 12588 31024 12591
rect 31076 12588 31082 12640
rect 1104 12538 32016 12560
rect 1104 12486 11253 12538
rect 11305 12486 11317 12538
rect 11369 12486 11381 12538
rect 11433 12486 11445 12538
rect 11497 12486 11509 12538
rect 11561 12486 21557 12538
rect 21609 12486 21621 12538
rect 21673 12486 21685 12538
rect 21737 12486 21749 12538
rect 21801 12486 21813 12538
rect 21865 12486 32016 12538
rect 1104 12464 32016 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 2593 12427 2651 12433
rect 2593 12424 2605 12427
rect 1820 12396 2605 12424
rect 1820 12384 1826 12396
rect 2593 12393 2605 12396
rect 2639 12393 2651 12427
rect 2593 12387 2651 12393
rect 3237 12427 3295 12433
rect 3237 12393 3249 12427
rect 3283 12424 3295 12427
rect 3602 12424 3608 12436
rect 3283 12396 3608 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 3786 12424 3792 12436
rect 3747 12396 3792 12424
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 9033 12427 9091 12433
rect 9033 12393 9045 12427
rect 9079 12424 9091 12427
rect 10042 12424 10048 12436
rect 9079 12396 10048 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 4154 12356 4160 12368
rect 3712 12328 4160 12356
rect 1394 12288 1400 12300
rect 1307 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12288 1458 12300
rect 2682 12288 2688 12300
rect 1452 12260 2688 12288
rect 1452 12248 1458 12260
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 3712 12297 3740 12328
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 5258 12316 5264 12368
rect 5316 12356 5322 12368
rect 7926 12356 7932 12368
rect 5316 12328 5672 12356
rect 5316 12316 5322 12328
rect 5644 12300 5672 12328
rect 5736 12328 7932 12356
rect 3697 12291 3755 12297
rect 3697 12257 3709 12291
rect 3743 12257 3755 12291
rect 3697 12251 3755 12257
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12288 3939 12291
rect 4522 12288 4528 12300
rect 3927 12260 4528 12288
rect 3927 12257 3939 12260
rect 3881 12251 3939 12257
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 5074 12288 5080 12300
rect 4755 12260 5080 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5350 12288 5356 12300
rect 5311 12260 5356 12288
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 5736 12297 5764 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6696 12260 7021 12288
rect 6696 12248 6702 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7009 12251 7067 12257
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 8205 12291 8263 12297
rect 8205 12288 8217 12291
rect 7248 12260 8217 12288
rect 7248 12248 7254 12260
rect 8205 12257 8217 12260
rect 8251 12257 8263 12291
rect 8205 12251 8263 12257
rect 8389 12291 8447 12297
rect 8389 12257 8401 12291
rect 8435 12288 8447 12291
rect 8754 12288 8760 12300
rect 8435 12260 8760 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4028 12192 4905 12220
rect 4028 12180 4034 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 5810 12220 5816 12232
rect 5316 12192 5816 12220
rect 5316 12180 5322 12192
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12220 7343 12223
rect 7374 12220 7380 12232
rect 7331 12192 7380 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 7374 12180 7380 12192
rect 7432 12220 7438 12232
rect 9048 12220 9076 12387
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10686 12424 10692 12436
rect 10244 12396 10692 12424
rect 10244 12297 10272 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 11848 12396 12265 12424
rect 11848 12384 11854 12396
rect 12253 12393 12265 12396
rect 12299 12424 12311 12427
rect 12342 12424 12348 12436
rect 12299 12396 12348 12424
rect 12299 12393 12311 12396
rect 12253 12387 12311 12393
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 13262 12424 13268 12436
rect 13223 12396 13268 12424
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 15470 12424 15476 12436
rect 15431 12396 15476 12424
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 15930 12424 15936 12436
rect 15891 12396 15936 12424
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 18138 12424 18144 12436
rect 17696 12396 18144 12424
rect 10318 12316 10324 12368
rect 10376 12356 10382 12368
rect 11885 12359 11943 12365
rect 11885 12356 11897 12359
rect 10376 12328 11897 12356
rect 10376 12316 10382 12328
rect 11885 12325 11897 12328
rect 11931 12325 11943 12359
rect 11885 12319 11943 12325
rect 12101 12359 12159 12365
rect 12101 12325 12113 12359
rect 12147 12356 12159 12359
rect 12434 12356 12440 12368
rect 12147 12328 12440 12356
rect 12147 12325 12159 12328
rect 12101 12319 12159 12325
rect 12434 12316 12440 12328
rect 12492 12316 12498 12368
rect 13081 12359 13139 12365
rect 13081 12325 13093 12359
rect 13127 12356 13139 12359
rect 13354 12356 13360 12368
rect 13127 12328 13360 12356
rect 13127 12325 13139 12328
rect 13081 12319 13139 12325
rect 13354 12316 13360 12328
rect 13412 12316 13418 12368
rect 14366 12365 14372 12368
rect 14360 12356 14372 12365
rect 14327 12328 14372 12356
rect 14360 12319 14372 12328
rect 14366 12316 14372 12319
rect 14424 12316 14430 12368
rect 15488 12356 15516 12384
rect 17402 12356 17408 12368
rect 15488 12328 17408 12356
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12257 10287 12291
rect 10410 12288 10416 12300
rect 10371 12260 10416 12288
rect 10229 12251 10287 12257
rect 7432 12192 9076 12220
rect 10244 12220 10272 12251
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 10778 12288 10784 12300
rect 10739 12260 10784 12288
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 12710 12288 12716 12300
rect 12671 12260 12716 12288
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 17696 12297 17724 12396
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 19426 12424 19432 12436
rect 18432 12396 19432 12424
rect 18432 12368 18460 12396
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 19518 12396 21220 12424
rect 17954 12316 17960 12368
rect 18012 12356 18018 12368
rect 18012 12328 18276 12356
rect 18012 12316 18018 12328
rect 17681 12291 17739 12297
rect 14056 12260 17080 12288
rect 14056 12248 14062 12260
rect 10318 12220 10324 12232
rect 10244 12192 10324 12220
rect 7432 12180 7438 12192
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10686 12220 10692 12232
rect 10643 12192 10692 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 10686 12180 10692 12192
rect 10744 12220 10750 12232
rect 11146 12220 11152 12232
rect 10744 12192 11152 12220
rect 10744 12180 10750 12192
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 14090 12220 14096 12232
rect 14051 12192 14096 12220
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 16022 12220 16028 12232
rect 15528 12192 16028 12220
rect 15528 12180 15534 12192
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 17052 12220 17080 12260
rect 17681 12257 17693 12291
rect 17727 12257 17739 12291
rect 17862 12288 17868 12300
rect 17823 12260 17868 12288
rect 17681 12251 17739 12257
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 18046 12288 18052 12300
rect 18007 12260 18052 12288
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18248 12297 18276 12328
rect 18414 12316 18420 12368
rect 18472 12316 18478 12368
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 19518 12356 19546 12396
rect 20070 12356 20076 12368
rect 18748 12328 19546 12356
rect 19639 12328 20076 12356
rect 18748 12316 18754 12328
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 19150 12288 19156 12300
rect 18279 12260 19156 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 19639 12288 19667 12328
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 21192 12356 21220 12396
rect 21910 12384 21916 12436
rect 21968 12424 21974 12436
rect 23290 12424 23296 12436
rect 21968 12396 23296 12424
rect 21968 12384 21974 12396
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 23477 12427 23535 12433
rect 23477 12393 23489 12427
rect 23523 12424 23535 12427
rect 24486 12424 24492 12436
rect 23523 12396 24492 12424
rect 23523 12393 23535 12396
rect 23477 12387 23535 12393
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 24673 12427 24731 12433
rect 24673 12393 24685 12427
rect 24719 12424 24731 12427
rect 25314 12424 25320 12436
rect 24719 12396 25320 12424
rect 24719 12393 24731 12396
rect 24673 12387 24731 12393
rect 25314 12384 25320 12396
rect 25372 12384 25378 12436
rect 25406 12384 25412 12436
rect 25464 12424 25470 12436
rect 25866 12424 25872 12436
rect 25464 12396 25872 12424
rect 25464 12384 25470 12396
rect 25866 12384 25872 12396
rect 25924 12424 25930 12436
rect 27338 12424 27344 12436
rect 25924 12396 26188 12424
rect 27299 12396 27344 12424
rect 25924 12384 25930 12396
rect 24578 12356 24584 12368
rect 21192 12328 21496 12356
rect 19794 12288 19800 12300
rect 19352 12260 19667 12288
rect 19755 12260 19800 12288
rect 19352 12232 19380 12260
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 21468 12288 21496 12328
rect 21836 12328 24584 12356
rect 21836 12288 21864 12328
rect 24578 12316 24584 12328
rect 24636 12316 24642 12368
rect 25222 12316 25228 12368
rect 25280 12356 25286 12368
rect 25786 12359 25844 12365
rect 25786 12356 25798 12359
rect 25280 12328 25798 12356
rect 25280 12316 25286 12328
rect 25786 12325 25798 12328
rect 25832 12325 25844 12359
rect 25786 12319 25844 12325
rect 19904 12260 21036 12288
rect 21468 12260 21864 12288
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17052 12192 17969 12220
rect 17957 12189 17969 12192
rect 18003 12220 18015 12223
rect 18414 12220 18420 12232
rect 18003 12192 18420 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 19334 12180 19340 12232
rect 19392 12180 19398 12232
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19484 12192 19625 12220
rect 19484 12180 19490 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 5077 12155 5135 12161
rect 5077 12121 5089 12155
rect 5123 12152 5135 12155
rect 13906 12152 13912 12164
rect 5123 12124 13912 12152
rect 5123 12121 5135 12124
rect 5077 12115 5135 12121
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 15930 12112 15936 12164
rect 15988 12152 15994 12164
rect 19904 12152 19932 12260
rect 19978 12180 19984 12232
rect 20036 12220 20042 12232
rect 20806 12220 20812 12232
rect 20036 12192 20812 12220
rect 20036 12180 20042 12192
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 15988 12124 19932 12152
rect 15988 12112 15994 12124
rect 20162 12112 20168 12164
rect 20220 12152 20226 12164
rect 21008 12152 21036 12260
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22189 12291 22247 12297
rect 22189 12288 22201 12291
rect 22152 12260 22201 12288
rect 22152 12248 22158 12260
rect 22189 12257 22201 12260
rect 22235 12257 22247 12291
rect 22738 12288 22744 12300
rect 22651 12260 22744 12288
rect 22189 12251 22247 12257
rect 22738 12248 22744 12260
rect 22796 12288 22802 12300
rect 23658 12288 23664 12300
rect 22796 12260 23664 12288
rect 22796 12248 22802 12260
rect 23658 12248 23664 12260
rect 23716 12248 23722 12300
rect 26050 12288 26056 12300
rect 26011 12260 26056 12288
rect 26050 12248 26056 12260
rect 26108 12248 26114 12300
rect 26160 12288 26188 12396
rect 27338 12384 27344 12396
rect 27396 12384 27402 12436
rect 29365 12427 29423 12433
rect 29365 12393 29377 12427
rect 29411 12424 29423 12427
rect 30282 12424 30288 12436
rect 29411 12396 30288 12424
rect 29411 12393 29423 12396
rect 29365 12387 29423 12393
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 30374 12384 30380 12436
rect 30432 12424 30438 12436
rect 31297 12427 31355 12433
rect 31297 12424 31309 12427
rect 30432 12396 31309 12424
rect 30432 12384 30438 12396
rect 31297 12393 31309 12396
rect 31343 12393 31355 12427
rect 31297 12387 31355 12393
rect 26602 12316 26608 12368
rect 26660 12356 26666 12368
rect 26973 12359 27031 12365
rect 26973 12356 26985 12359
rect 26660 12328 26985 12356
rect 26660 12316 26666 12328
rect 26973 12325 26985 12328
rect 27019 12325 27031 12359
rect 26973 12319 27031 12325
rect 27189 12359 27247 12365
rect 27189 12325 27201 12359
rect 27235 12356 27247 12359
rect 27706 12356 27712 12368
rect 27235 12328 27712 12356
rect 27235 12325 27247 12328
rect 27189 12319 27247 12325
rect 27706 12316 27712 12328
rect 27764 12316 27770 12368
rect 30190 12365 30196 12368
rect 30184 12356 30196 12365
rect 30151 12328 30196 12356
rect 30184 12319 30196 12328
rect 30190 12316 30196 12319
rect 30248 12316 30254 12368
rect 27893 12291 27951 12297
rect 27893 12288 27905 12291
rect 26160 12260 27905 12288
rect 27893 12257 27905 12260
rect 27939 12257 27951 12291
rect 27893 12251 27951 12257
rect 28442 12248 28448 12300
rect 28500 12288 28506 12300
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 28500 12260 28549 12288
rect 28500 12248 28506 12260
rect 28537 12257 28549 12260
rect 28583 12257 28595 12291
rect 28537 12251 28595 12257
rect 29273 12291 29331 12297
rect 29273 12257 29285 12291
rect 29319 12288 29331 12291
rect 29730 12288 29736 12300
rect 29319 12260 29736 12288
rect 29319 12257 29331 12260
rect 29273 12251 29331 12257
rect 29730 12248 29736 12260
rect 29788 12248 29794 12300
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 21358 12220 21364 12232
rect 21315 12192 21364 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 21542 12180 21548 12232
rect 21600 12220 21606 12232
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21600 12192 21925 12220
rect 21600 12180 21606 12192
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 22922 12220 22928 12232
rect 22883 12192 22928 12220
rect 21913 12183 21971 12189
rect 22922 12180 22928 12192
rect 22980 12180 22986 12232
rect 23937 12223 23995 12229
rect 23937 12189 23949 12223
rect 23983 12220 23995 12223
rect 24762 12220 24768 12232
rect 23983 12192 24768 12220
rect 23983 12189 23995 12192
rect 23937 12183 23995 12189
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 28626 12220 28632 12232
rect 26206 12192 28632 12220
rect 21818 12152 21824 12164
rect 20220 12124 20944 12152
rect 21008 12124 21824 12152
rect 20220 12112 20226 12124
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4430 12084 4436 12096
rect 4212 12056 4436 12084
rect 4212 12044 4218 12056
rect 4430 12044 4436 12056
rect 4488 12044 4494 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 9398 12084 9404 12096
rect 9272 12056 9404 12084
rect 9272 12044 9278 12056
rect 9398 12044 9404 12056
rect 9456 12084 9462 12096
rect 9585 12087 9643 12093
rect 9585 12084 9597 12087
rect 9456 12056 9597 12084
rect 9456 12044 9462 12056
rect 9585 12053 9597 12056
rect 9631 12053 9643 12087
rect 9585 12047 9643 12053
rect 10965 12087 11023 12093
rect 10965 12053 10977 12087
rect 11011 12084 11023 12087
rect 11698 12084 11704 12096
rect 11011 12056 11704 12084
rect 11011 12053 11023 12056
rect 10965 12047 11023 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12250 12084 12256 12096
rect 12115 12056 12256 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 12952 12056 13093 12084
rect 12952 12044 12958 12056
rect 13081 12053 13093 12056
rect 13127 12053 13139 12087
rect 13081 12047 13139 12053
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16669 12087 16727 12093
rect 16669 12084 16681 12087
rect 16080 12056 16681 12084
rect 16080 12044 16086 12056
rect 16669 12053 16681 12056
rect 16715 12053 16727 12087
rect 16669 12047 16727 12053
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 17497 12087 17555 12093
rect 17497 12084 17509 12087
rect 17460 12056 17509 12084
rect 17460 12044 17466 12056
rect 17497 12053 17509 12056
rect 17543 12053 17555 12087
rect 18690 12084 18696 12096
rect 18651 12056 18696 12084
rect 17497 12047 17555 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 19886 12044 19892 12096
rect 19944 12084 19950 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19944 12056 19993 12084
rect 19944 12044 19950 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 20438 12084 20444 12096
rect 20399 12056 20444 12084
rect 19981 12047 20039 12053
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 20916 12084 20944 12124
rect 21818 12112 21824 12124
rect 21876 12112 21882 12164
rect 23768 12124 25185 12152
rect 23768 12084 23796 12124
rect 20916 12056 23796 12084
rect 23845 12087 23903 12093
rect 23845 12053 23857 12087
rect 23891 12084 23903 12087
rect 24394 12084 24400 12096
rect 23891 12056 24400 12084
rect 23891 12053 23903 12056
rect 23845 12047 23903 12053
rect 24394 12044 24400 12056
rect 24452 12044 24458 12096
rect 25157 12084 25185 12124
rect 26206 12084 26234 12192
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 29546 12180 29552 12232
rect 29604 12220 29610 12232
rect 29917 12223 29975 12229
rect 29917 12220 29929 12223
rect 29604 12192 29929 12220
rect 29604 12180 29610 12192
rect 29917 12189 29929 12192
rect 29963 12189 29975 12223
rect 29917 12183 29975 12189
rect 28350 12112 28356 12164
rect 28408 12152 28414 12164
rect 29638 12152 29644 12164
rect 28408 12124 29644 12152
rect 28408 12112 28414 12124
rect 29638 12112 29644 12124
rect 29696 12112 29702 12164
rect 27154 12084 27160 12096
rect 25157 12056 26234 12084
rect 27115 12056 27160 12084
rect 27154 12044 27160 12056
rect 27212 12044 27218 12096
rect 27890 12044 27896 12096
rect 27948 12084 27954 12096
rect 28445 12087 28503 12093
rect 28445 12084 28457 12087
rect 27948 12056 28457 12084
rect 27948 12044 27954 12056
rect 28445 12053 28457 12056
rect 28491 12053 28503 12087
rect 28445 12047 28503 12053
rect 1104 11994 32016 12016
rect 1104 11942 6102 11994
rect 6154 11942 6166 11994
rect 6218 11942 6230 11994
rect 6282 11942 6294 11994
rect 6346 11942 6358 11994
rect 6410 11942 16405 11994
rect 16457 11942 16469 11994
rect 16521 11942 16533 11994
rect 16585 11942 16597 11994
rect 16649 11942 16661 11994
rect 16713 11942 26709 11994
rect 26761 11942 26773 11994
rect 26825 11942 26837 11994
rect 26889 11942 26901 11994
rect 26953 11942 26965 11994
rect 27017 11942 32016 11994
rect 1104 11920 32016 11942
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 9490 11880 9496 11892
rect 4172 11852 9496 11880
rect 2774 11812 2780 11824
rect 1596 11784 2780 11812
rect 1596 11685 1624 11784
rect 2774 11772 2780 11784
rect 2832 11772 2838 11824
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2866 11744 2872 11756
rect 1995 11716 2872 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2866 11704 2872 11716
rect 2924 11744 2930 11756
rect 3326 11744 3332 11756
rect 2924 11716 3332 11744
rect 2924 11704 2930 11716
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11645 1639 11679
rect 1581 11639 1639 11645
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11645 1823 11679
rect 1765 11639 1823 11645
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2314 11676 2320 11688
rect 2179 11648 2320 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 1780 11608 1808 11639
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 2958 11676 2964 11688
rect 2823 11648 2964 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 4172 11685 4200 11852
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 13354 11880 13360 11892
rect 9640 11852 9685 11880
rect 13315 11852 13360 11880
rect 9640 11840 9646 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 14369 11883 14427 11889
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 14550 11880 14556 11892
rect 14415 11852 14556 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 16114 11880 16120 11892
rect 15896 11852 16120 11880
rect 15896 11840 15902 11852
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 19610 11880 19616 11892
rect 19536 11852 19616 11880
rect 5442 11812 5448 11824
rect 5403 11784 5448 11812
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 5534 11772 5540 11824
rect 5592 11772 5598 11824
rect 10226 11772 10232 11824
rect 10284 11812 10290 11824
rect 10502 11812 10508 11824
rect 10284 11784 10508 11812
rect 10284 11772 10290 11784
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 13906 11772 13912 11824
rect 13964 11812 13970 11824
rect 18598 11812 18604 11824
rect 13964 11784 18604 11812
rect 13964 11772 13970 11784
rect 18598 11772 18604 11784
rect 18656 11772 18662 11824
rect 5552 11744 5580 11772
rect 6086 11744 6092 11756
rect 5552 11716 6092 11744
rect 6086 11704 6092 11716
rect 6144 11744 6150 11756
rect 7006 11744 7012 11756
rect 6144 11716 6592 11744
rect 6144 11704 6150 11716
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4430 11636 4436 11688
rect 4488 11676 4494 11688
rect 6564 11685 6592 11716
rect 6656 11716 7012 11744
rect 6365 11679 6423 11685
rect 6365 11676 6377 11679
rect 4488 11648 6377 11676
rect 4488 11636 4494 11648
rect 6365 11645 6377 11648
rect 6411 11645 6423 11679
rect 6365 11639 6423 11645
rect 6549 11679 6607 11685
rect 6549 11645 6561 11679
rect 6595 11645 6607 11679
rect 6549 11639 6607 11645
rect 2038 11608 2044 11620
rect 1780 11580 2044 11608
rect 2038 11568 2044 11580
rect 2096 11608 2102 11620
rect 3878 11608 3884 11620
rect 2096 11580 3884 11608
rect 2096 11568 2102 11580
rect 3878 11568 3884 11580
rect 3936 11568 3942 11620
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 6656 11608 6684 11716
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 10468 11716 11161 11744
rect 10468 11704 10474 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 15252 11716 15577 11744
rect 15252 11704 15258 11716
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 19334 11744 19340 11756
rect 15565 11707 15623 11713
rect 16684 11716 19340 11744
rect 7282 11685 7288 11688
rect 7276 11639 7288 11685
rect 7340 11676 7346 11688
rect 9766 11676 9772 11688
rect 7340 11648 7376 11676
rect 9727 11648 9772 11676
rect 7282 11636 7288 11639
rect 7340 11636 7346 11648
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 9950 11676 9956 11688
rect 9911 11648 9956 11676
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11645 10195 11679
rect 10318 11676 10324 11688
rect 10279 11648 10324 11676
rect 10137 11639 10195 11645
rect 10060 11608 10088 11639
rect 5500 11580 6684 11608
rect 9048 11580 10088 11608
rect 10152 11608 10180 11639
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11676 11391 11679
rect 11790 11676 11796 11688
rect 11379 11648 11796 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 11974 11676 11980 11688
rect 11935 11648 11980 11676
rect 11974 11636 11980 11648
rect 12032 11676 12038 11688
rect 16684 11676 16712 11716
rect 19334 11704 19340 11716
rect 19392 11704 19398 11756
rect 19536 11744 19564 11852
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 20622 11880 20628 11892
rect 19812 11852 20628 11880
rect 19702 11772 19708 11824
rect 19760 11812 19766 11824
rect 19812 11812 19840 11852
rect 20622 11840 20628 11852
rect 20680 11880 20686 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20680 11852 20821 11880
rect 20680 11840 20686 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 20993 11883 21051 11889
rect 20993 11849 21005 11883
rect 21039 11880 21051 11883
rect 21542 11880 21548 11892
rect 21039 11852 21548 11880
rect 21039 11849 21051 11852
rect 20993 11843 21051 11849
rect 21542 11840 21548 11852
rect 21600 11840 21606 11892
rect 21913 11883 21971 11889
rect 21913 11849 21925 11883
rect 21959 11849 21971 11883
rect 21913 11843 21971 11849
rect 21266 11812 21272 11824
rect 19760 11784 19840 11812
rect 19760 11772 19766 11784
rect 19613 11747 19671 11753
rect 19613 11744 19625 11747
rect 19536 11716 19625 11744
rect 19613 11713 19625 11716
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 12032 11648 16712 11676
rect 16761 11679 16819 11685
rect 12032 11636 12038 11648
rect 16761 11645 16773 11679
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 17037 11679 17095 11685
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 17126 11676 17132 11688
rect 17083 11648 17132 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 10226 11608 10232 11620
rect 10152 11580 10232 11608
rect 5500 11568 5506 11580
rect 2317 11543 2375 11549
rect 2317 11509 2329 11543
rect 2363 11540 2375 11543
rect 2498 11540 2504 11552
rect 2363 11512 2504 11540
rect 2363 11509 2375 11512
rect 2317 11503 2375 11509
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 6454 11540 6460 11552
rect 6415 11512 6460 11540
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 7708 11512 8401 11540
rect 7708 11500 7714 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9048 11549 9076 11580
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8536 11512 9045 11540
rect 8536 11500 8542 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 10060 11540 10088 11580
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 12250 11617 12256 11620
rect 12244 11571 12256 11617
rect 12308 11608 12314 11620
rect 14921 11611 14979 11617
rect 12308 11580 12344 11608
rect 12250 11568 12256 11571
rect 12308 11568 12314 11580
rect 14921 11577 14933 11611
rect 14967 11608 14979 11611
rect 14967 11580 15700 11608
rect 14967 11577 14979 11580
rect 14921 11571 14979 11577
rect 10594 11540 10600 11552
rect 10060 11512 10600 11540
rect 9033 11503 9091 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 11517 11543 11575 11549
rect 11517 11509 11529 11543
rect 11563 11540 11575 11543
rect 11790 11540 11796 11552
rect 11563 11512 11796 11540
rect 11563 11509 11575 11512
rect 11517 11503 11575 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 15010 11540 15016 11552
rect 14971 11512 15016 11540
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15672 11540 15700 11580
rect 15746 11568 15752 11620
rect 15804 11608 15810 11620
rect 16776 11608 16804 11639
rect 17126 11636 17132 11648
rect 17184 11676 17190 11688
rect 17862 11676 17868 11688
rect 17184 11648 17868 11676
rect 17184 11636 17190 11648
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 19150 11636 19156 11688
rect 19208 11676 19214 11688
rect 19245 11679 19303 11685
rect 19245 11676 19257 11679
rect 19208 11648 19257 11676
rect 19208 11636 19214 11648
rect 19245 11645 19257 11648
rect 19291 11645 19303 11679
rect 19426 11676 19432 11688
rect 19387 11648 19432 11676
rect 19245 11639 19303 11645
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 19812 11685 19840 11784
rect 20456 11784 21272 11812
rect 20456 11685 20484 11784
rect 21266 11772 21272 11784
rect 21324 11812 21330 11824
rect 21928 11812 21956 11843
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 24394 11880 24400 11892
rect 22152 11852 22197 11880
rect 24355 11852 24400 11880
rect 22152 11840 22158 11852
rect 24394 11840 24400 11852
rect 24452 11840 24458 11892
rect 24486 11840 24492 11892
rect 24544 11880 24550 11892
rect 24581 11883 24639 11889
rect 24581 11880 24593 11883
rect 24544 11852 24593 11880
rect 24544 11840 24550 11852
rect 24581 11849 24593 11852
rect 24627 11880 24639 11883
rect 25406 11880 25412 11892
rect 24627 11852 25412 11880
rect 24627 11849 24639 11852
rect 24581 11843 24639 11849
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 29822 11880 29828 11892
rect 25884 11852 26280 11880
rect 25884 11812 25912 11852
rect 21324 11784 21956 11812
rect 23308 11784 25912 11812
rect 21324 11772 21330 11784
rect 20622 11704 20628 11756
rect 20680 11744 20686 11756
rect 21545 11747 21603 11753
rect 21545 11744 21557 11747
rect 20680 11716 21557 11744
rect 20680 11704 20686 11716
rect 21545 11713 21557 11716
rect 21591 11713 21603 11747
rect 21545 11707 21603 11713
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 23308 11753 23336 11784
rect 25958 11772 25964 11824
rect 26016 11812 26022 11824
rect 26053 11815 26111 11821
rect 26053 11812 26065 11815
rect 26016 11784 26065 11812
rect 26016 11772 26022 11784
rect 26053 11781 26065 11784
rect 26099 11781 26111 11815
rect 26053 11775 26111 11781
rect 23293 11747 23351 11753
rect 23293 11744 23305 11747
rect 22244 11716 23305 11744
rect 22244 11704 22250 11716
rect 23293 11713 23305 11716
rect 23339 11713 23351 11747
rect 23293 11707 23351 11713
rect 25314 11704 25320 11756
rect 25372 11744 25378 11756
rect 25774 11744 25780 11756
rect 25372 11716 25780 11744
rect 25372 11704 25378 11716
rect 25774 11704 25780 11716
rect 25832 11744 25838 11756
rect 25832 11716 26188 11744
rect 25832 11704 25838 11716
rect 19521 11679 19579 11685
rect 19521 11645 19533 11679
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 19797 11679 19855 11685
rect 19797 11645 19809 11679
rect 19843 11645 19855 11679
rect 19797 11639 19855 11645
rect 20441 11679 20499 11685
rect 20441 11645 20453 11679
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 16850 11608 16856 11620
rect 15804 11580 16856 11608
rect 15804 11568 15810 11580
rect 16850 11568 16856 11580
rect 16908 11608 16914 11620
rect 18230 11608 18236 11620
rect 16908 11580 18236 11608
rect 16908 11568 16914 11580
rect 18230 11568 18236 11580
rect 18288 11608 18294 11620
rect 18601 11611 18659 11617
rect 18601 11608 18613 11611
rect 18288 11580 18613 11608
rect 18288 11568 18294 11580
rect 18601 11577 18613 11580
rect 18647 11577 18659 11611
rect 18601 11571 18659 11577
rect 16022 11540 16028 11552
rect 15672 11512 16028 11540
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 17678 11540 17684 11552
rect 17000 11512 17684 11540
rect 17000 11500 17006 11512
rect 17678 11500 17684 11512
rect 17736 11540 17742 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17736 11512 18061 11540
rect 17736 11500 17742 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 19536 11540 19564 11639
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 22830 11676 22836 11688
rect 22520 11648 22836 11676
rect 22520 11636 22526 11648
rect 22830 11636 22836 11648
rect 22888 11676 22894 11688
rect 23017 11679 23075 11685
rect 23017 11676 23029 11679
rect 22888 11648 23029 11676
rect 22888 11636 22894 11648
rect 23017 11645 23029 11648
rect 23063 11645 23075 11679
rect 24946 11676 24952 11688
rect 24907 11648 24952 11676
rect 23017 11639 23075 11645
rect 24946 11636 24952 11648
rect 25004 11636 25010 11688
rect 25682 11676 25688 11688
rect 25643 11648 25688 11676
rect 25682 11636 25688 11648
rect 25740 11636 25746 11688
rect 25866 11676 25872 11688
rect 25827 11648 25872 11676
rect 25866 11636 25872 11648
rect 25924 11636 25930 11688
rect 26160 11685 26188 11716
rect 25961 11679 26019 11685
rect 25961 11645 25973 11679
rect 26007 11645 26019 11679
rect 25961 11639 26019 11645
rect 26145 11679 26203 11685
rect 26145 11645 26157 11679
rect 26191 11645 26203 11679
rect 26252 11676 26280 11852
rect 28552 11852 29828 11880
rect 28552 11753 28580 11852
rect 29822 11840 29828 11852
rect 29880 11840 29886 11892
rect 30742 11840 30748 11892
rect 30800 11880 30806 11892
rect 30929 11883 30987 11889
rect 30929 11880 30941 11883
rect 30800 11852 30941 11880
rect 30800 11840 30806 11852
rect 30929 11849 30941 11852
rect 30975 11849 30987 11883
rect 30929 11843 30987 11849
rect 28644 11784 29960 11812
rect 28644 11753 28672 11784
rect 28537 11747 28595 11753
rect 27632 11716 28488 11744
rect 26510 11676 26516 11688
rect 26252 11648 26516 11676
rect 26145 11639 26203 11645
rect 19812 11580 20116 11608
rect 19812 11552 19840 11580
rect 18472 11512 19564 11540
rect 18472 11500 18478 11512
rect 19794 11500 19800 11552
rect 19852 11500 19858 11552
rect 19978 11540 19984 11552
rect 19939 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20088 11540 20116 11580
rect 22922 11568 22928 11620
rect 22980 11608 22986 11620
rect 25976 11608 26004 11639
rect 26510 11636 26516 11648
rect 26568 11676 26574 11688
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 26568 11648 26985 11676
rect 26568 11636 26574 11648
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 27154 11676 27160 11688
rect 27115 11648 27160 11676
rect 26973 11639 27031 11645
rect 27154 11636 27160 11648
rect 27212 11636 27218 11688
rect 27338 11636 27344 11688
rect 27396 11676 27402 11688
rect 27632 11685 27660 11716
rect 28460 11688 28488 11716
rect 28537 11713 28549 11747
rect 28583 11713 28595 11747
rect 28537 11707 28595 11713
rect 28629 11747 28687 11753
rect 28629 11713 28641 11747
rect 28675 11713 28687 11747
rect 28629 11707 28687 11713
rect 28718 11704 28724 11756
rect 28776 11744 28782 11756
rect 29822 11744 29828 11756
rect 28776 11716 29592 11744
rect 29783 11716 29828 11744
rect 28776 11704 28782 11716
rect 27617 11679 27675 11685
rect 27617 11676 27629 11679
rect 27396 11648 27629 11676
rect 27396 11636 27402 11648
rect 27617 11645 27629 11648
rect 27663 11645 27675 11679
rect 27617 11639 27675 11645
rect 27801 11679 27859 11685
rect 27801 11645 27813 11679
rect 27847 11676 27859 11679
rect 27890 11676 27896 11688
rect 27847 11648 27896 11676
rect 27847 11645 27859 11648
rect 27801 11639 27859 11645
rect 27890 11636 27896 11648
rect 27948 11636 27954 11688
rect 28261 11679 28319 11685
rect 28261 11645 28273 11679
rect 28307 11676 28319 11679
rect 28350 11676 28356 11688
rect 28307 11648 28356 11676
rect 28307 11645 28319 11648
rect 28261 11639 28319 11645
rect 28350 11636 28356 11648
rect 28408 11636 28414 11688
rect 28442 11636 28448 11688
rect 28500 11676 28506 11688
rect 29564 11685 29592 11716
rect 29822 11704 29828 11716
rect 29880 11704 29886 11756
rect 29932 11753 29960 11784
rect 29917 11747 29975 11753
rect 29917 11713 29929 11747
rect 29963 11744 29975 11747
rect 30006 11744 30012 11756
rect 29963 11716 30012 11744
rect 29963 11713 29975 11716
rect 29917 11707 29975 11713
rect 30006 11704 30012 11716
rect 30064 11704 30070 11756
rect 30834 11744 30840 11756
rect 30795 11716 30840 11744
rect 30834 11704 30840 11716
rect 30892 11704 30898 11756
rect 28813 11679 28871 11685
rect 28500 11648 28545 11676
rect 28500 11636 28506 11648
rect 28813 11645 28825 11679
rect 28859 11678 28871 11679
rect 29549 11679 29607 11685
rect 28859 11676 28948 11678
rect 28859 11650 29040 11676
rect 28859 11645 28871 11650
rect 28920 11648 29040 11650
rect 28813 11639 28871 11645
rect 27522 11608 27528 11620
rect 22980 11580 27528 11608
rect 22980 11568 22986 11580
rect 27522 11568 27528 11580
rect 27580 11568 27586 11620
rect 29012 11608 29040 11648
rect 29549 11645 29561 11679
rect 29595 11645 29607 11679
rect 29730 11676 29736 11688
rect 29691 11648 29736 11676
rect 29549 11639 29607 11645
rect 29730 11636 29736 11648
rect 29788 11636 29794 11688
rect 30101 11679 30159 11685
rect 30101 11645 30113 11679
rect 30147 11676 30159 11679
rect 30926 11676 30932 11688
rect 30147 11648 30932 11676
rect 30147 11645 30159 11648
rect 30101 11639 30159 11645
rect 30926 11636 30932 11648
rect 30984 11636 30990 11688
rect 31110 11676 31116 11688
rect 31071 11648 31116 11676
rect 31110 11636 31116 11648
rect 31168 11636 31174 11688
rect 29748 11608 29776 11636
rect 29012 11580 29776 11608
rect 20818 11543 20876 11549
rect 20818 11540 20830 11543
rect 20088 11512 20830 11540
rect 20818 11509 20830 11512
rect 20864 11509 20876 11543
rect 21910 11540 21916 11552
rect 21871 11512 21916 11540
rect 20818 11503 20876 11509
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 24302 11500 24308 11552
rect 24360 11540 24366 11552
rect 24581 11543 24639 11549
rect 24581 11540 24593 11543
rect 24360 11512 24593 11540
rect 24360 11500 24366 11512
rect 24581 11509 24593 11512
rect 24627 11509 24639 11543
rect 24581 11503 24639 11509
rect 26329 11543 26387 11549
rect 26329 11509 26341 11543
rect 26375 11540 26387 11543
rect 26602 11540 26608 11552
rect 26375 11512 26608 11540
rect 26375 11509 26387 11512
rect 26329 11503 26387 11509
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 27062 11540 27068 11552
rect 27023 11512 27068 11540
rect 27062 11500 27068 11512
rect 27120 11500 27126 11552
rect 27614 11540 27620 11552
rect 27575 11512 27620 11540
rect 27614 11500 27620 11512
rect 27672 11500 27678 11552
rect 28997 11543 29055 11549
rect 28997 11509 29009 11543
rect 29043 11540 29055 11543
rect 29638 11540 29644 11552
rect 29043 11512 29644 11540
rect 29043 11509 29055 11512
rect 28997 11503 29055 11509
rect 29638 11500 29644 11512
rect 29696 11500 29702 11552
rect 30282 11540 30288 11552
rect 30243 11512 30288 11540
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 31110 11500 31116 11552
rect 31168 11540 31174 11552
rect 31297 11543 31355 11549
rect 31297 11540 31309 11543
rect 31168 11512 31309 11540
rect 31168 11500 31174 11512
rect 31297 11509 31309 11512
rect 31343 11509 31355 11543
rect 31297 11503 31355 11509
rect 1104 11450 32016 11472
rect 1104 11398 11253 11450
rect 11305 11398 11317 11450
rect 11369 11398 11381 11450
rect 11433 11398 11445 11450
rect 11497 11398 11509 11450
rect 11561 11398 21557 11450
rect 21609 11398 21621 11450
rect 21673 11398 21685 11450
rect 21737 11398 21749 11450
rect 21801 11398 21813 11450
rect 21865 11398 32016 11450
rect 1104 11376 32016 11398
rect 2958 11336 2964 11348
rect 1412 11308 2964 11336
rect 0 11268 800 11282
rect 1412 11268 1440 11308
rect 2958 11296 2964 11308
rect 3016 11336 3022 11348
rect 3326 11336 3332 11348
rect 3016 11308 3332 11336
rect 3016 11296 3022 11308
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4614 11336 4620 11348
rect 4120 11308 4620 11336
rect 4120 11296 4126 11308
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5074 11336 5080 11348
rect 4764 11308 5080 11336
rect 4764 11296 4770 11308
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 5350 11296 5356 11348
rect 5408 11336 5414 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 5408 11308 5457 11336
rect 5408 11296 5414 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5445 11299 5503 11305
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 5994 11336 6000 11348
rect 5868 11308 6000 11336
rect 5868 11296 5874 11308
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 8754 11336 8760 11348
rect 8715 11308 8760 11336
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 10042 11336 10048 11348
rect 9447 11308 10048 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12250 11336 12256 11348
rect 12207 11308 12256 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12618 11336 12624 11348
rect 12579 11308 12624 11336
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 15565 11339 15623 11345
rect 15565 11305 15577 11339
rect 15611 11336 15623 11339
rect 16022 11336 16028 11348
rect 15611 11308 16028 11336
rect 15611 11305 15623 11308
rect 15565 11299 15623 11305
rect 2866 11268 2872 11280
rect 0 11240 1440 11268
rect 2148 11240 2872 11268
rect 0 11226 800 11240
rect 1578 11160 1584 11212
rect 1636 11200 1642 11212
rect 1762 11200 1768 11212
rect 1636 11172 1768 11200
rect 1636 11160 1642 11172
rect 1762 11160 1768 11172
rect 1820 11200 1826 11212
rect 2148 11209 2176 11240
rect 2866 11228 2872 11240
rect 2924 11228 2930 11280
rect 3878 11268 3884 11280
rect 3160 11240 3884 11268
rect 1949 11203 2007 11209
rect 1949 11200 1961 11203
rect 1820 11172 1961 11200
rect 1820 11160 1826 11172
rect 1949 11169 1961 11172
rect 1995 11169 2007 11203
rect 1949 11163 2007 11169
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11169 2191 11203
rect 2314 11200 2320 11212
rect 2275 11172 2320 11200
rect 2133 11163 2191 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2774 11200 2780 11212
rect 2547 11172 2780 11200
rect 2547 11170 2575 11172
rect 2547 11169 2559 11170
rect 2501 11163 2559 11169
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 3160 11209 3188 11240
rect 3878 11228 3884 11240
rect 3936 11228 3942 11280
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 6454 11268 6460 11280
rect 4396 11240 4936 11268
rect 4396 11228 4402 11240
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11169 3203 11203
rect 3145 11163 3203 11169
rect 3234 11160 3240 11212
rect 3292 11200 3298 11212
rect 4908 11209 4936 11240
rect 5368 11240 6460 11268
rect 5368 11212 5396 11240
rect 6454 11228 6460 11240
rect 6512 11277 6518 11280
rect 6512 11271 6575 11277
rect 6512 11237 6529 11271
rect 6563 11237 6575 11271
rect 6730 11268 6736 11280
rect 6691 11240 6736 11268
rect 6512 11231 6575 11237
rect 6512 11228 6518 11231
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 7622 11271 7680 11277
rect 7622 11268 7634 11271
rect 7524 11240 7634 11268
rect 7524 11228 7530 11240
rect 7622 11237 7634 11240
rect 7668 11237 7680 11271
rect 12636 11268 12664 11296
rect 7622 11231 7680 11237
rect 10152 11240 12664 11268
rect 13449 11271 13507 11277
rect 3513 11203 3571 11209
rect 3513 11200 3525 11203
rect 3292 11172 3525 11200
rect 3292 11160 3298 11172
rect 3513 11169 3525 11172
rect 3559 11169 3571 11203
rect 3513 11163 3571 11169
rect 3697 11203 3755 11209
rect 3697 11169 3709 11203
rect 3743 11169 3755 11203
rect 3697 11163 3755 11169
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 1912 11104 2237 11132
rect 1912 11092 1918 11104
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 1762 11064 1768 11076
rect 1723 11036 1768 11064
rect 1762 11024 1768 11036
rect 1820 11024 1826 11076
rect 2792 11064 2820 11160
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 3329 11135 3387 11141
rect 3329 11132 3341 11135
rect 2924 11104 3341 11132
rect 2924 11092 2930 11104
rect 3329 11101 3341 11104
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3602 11132 3608 11144
rect 3467 11104 3608 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 3712 11064 3740 11163
rect 4706 11132 4712 11144
rect 4667 11104 4712 11132
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 4798 11092 4804 11144
rect 4856 11132 4862 11144
rect 4908 11132 4936 11163
rect 5350 11160 5356 11212
rect 5408 11160 5414 11212
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5491 11172 6592 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 4856 11104 4936 11132
rect 5077 11135 5135 11141
rect 4856 11092 4862 11104
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 6454 11132 6460 11144
rect 5123 11104 6460 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 2792 11036 3740 11064
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 4890 11064 4896 11076
rect 4396 11036 4896 11064
rect 4396 11024 4402 11036
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 2958 10996 2964 11008
rect 2919 10968 2964 10996
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 3878 10956 3884 11008
rect 3936 10996 3942 11008
rect 5092 10996 5120 11095
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6086 11064 6092 11076
rect 5920 11036 6092 11064
rect 5920 11008 5948 11036
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 6365 11067 6423 11073
rect 6365 11033 6377 11067
rect 6411 11064 6423 11067
rect 6564 11064 6592 11172
rect 7006 11160 7012 11212
rect 7064 11200 7070 11212
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 7064 11172 7389 11200
rect 7064 11160 7070 11172
rect 7377 11169 7389 11172
rect 7423 11169 7435 11203
rect 9214 11200 9220 11212
rect 9175 11172 9220 11200
rect 7377 11163 7435 11169
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 10152 11209 10180 11240
rect 13449 11237 13461 11271
rect 13495 11268 13507 11271
rect 14001 11271 14059 11277
rect 14001 11268 14013 11271
rect 13495 11240 14013 11268
rect 13495 11237 13507 11240
rect 13449 11231 13507 11237
rect 14001 11237 14013 11240
rect 14047 11268 14059 11271
rect 15580 11268 15608 11299
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16850 11336 16856 11348
rect 16811 11308 16856 11336
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 19058 11336 19064 11348
rect 17328 11308 19064 11336
rect 16942 11268 16948 11280
rect 14047 11240 15608 11268
rect 16903 11240 16948 11268
rect 14047 11237 14059 11240
rect 14001 11231 14059 11237
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 11790 11160 11796 11212
rect 11848 11200 11854 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11848 11172 11989 11200
rect 11848 11160 11854 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 11977 11163 12035 11169
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 13464 11200 13492 11231
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 12124 11172 13492 11200
rect 12124 11160 12130 11172
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14608 11172 14749 11200
rect 14608 11160 14614 11172
rect 14737 11169 14749 11172
rect 14783 11200 14795 11203
rect 14918 11200 14924 11212
rect 14783 11172 14924 11200
rect 14783 11169 14795 11172
rect 14737 11163 14795 11169
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 15930 11200 15936 11212
rect 15519 11172 15936 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 10410 11132 10416 11144
rect 10371 11104 10416 11132
rect 10410 11092 10416 11104
rect 10468 11132 10474 11144
rect 10686 11132 10692 11144
rect 10468 11104 10692 11132
rect 10468 11092 10474 11104
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 14056 11104 14197 11132
rect 14056 11092 14062 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 17328 11132 17356 11308
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 20717 11339 20775 11345
rect 20717 11336 20729 11339
rect 20680 11308 20729 11336
rect 20680 11296 20686 11308
rect 20717 11305 20729 11308
rect 20763 11305 20775 11339
rect 20717 11299 20775 11305
rect 22281 11339 22339 11345
rect 22281 11305 22293 11339
rect 22327 11336 22339 11339
rect 24118 11336 24124 11348
rect 22327 11308 24124 11336
rect 22327 11305 22339 11308
rect 22281 11299 22339 11305
rect 24118 11296 24124 11308
rect 24176 11296 24182 11348
rect 24302 11336 24308 11348
rect 24263 11308 24308 11336
rect 24302 11296 24308 11308
rect 24360 11296 24366 11348
rect 25866 11336 25872 11348
rect 25827 11308 25872 11336
rect 25866 11296 25872 11308
rect 25924 11296 25930 11348
rect 27154 11336 27160 11348
rect 27115 11308 27160 11336
rect 27154 11296 27160 11308
rect 27212 11296 27218 11348
rect 28442 11296 28448 11348
rect 28500 11336 28506 11348
rect 28994 11336 29000 11348
rect 28500 11308 29000 11336
rect 28500 11296 28506 11308
rect 28994 11296 29000 11308
rect 29052 11296 29058 11348
rect 30561 11339 30619 11345
rect 30561 11305 30573 11339
rect 30607 11336 30619 11339
rect 30650 11336 30656 11348
rect 30607 11308 30656 11336
rect 30607 11305 30619 11308
rect 30561 11299 30619 11305
rect 30650 11296 30656 11308
rect 30708 11296 30714 11348
rect 31297 11339 31355 11345
rect 31297 11305 31309 11339
rect 31343 11336 31355 11339
rect 31343 11308 31754 11336
rect 31343 11305 31355 11308
rect 31297 11299 31355 11305
rect 19604 11271 19662 11277
rect 17512 11240 19196 11268
rect 17512 11209 17540 11240
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11169 17555 11203
rect 17753 11203 17811 11209
rect 17753 11200 17765 11203
rect 17497 11163 17555 11169
rect 17604 11172 17765 11200
rect 14185 11095 14243 11101
rect 14844 11104 17356 11132
rect 14844 11064 14872 11104
rect 17402 11092 17408 11144
rect 17460 11132 17466 11144
rect 17604 11132 17632 11172
rect 17753 11169 17765 11172
rect 17799 11169 17811 11203
rect 17753 11163 17811 11169
rect 19168 11144 19196 11240
rect 19604 11237 19616 11271
rect 19650 11268 19662 11271
rect 19978 11268 19984 11280
rect 19650 11240 19984 11268
rect 19650 11237 19662 11240
rect 19604 11231 19662 11237
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 24995 11271 25053 11277
rect 24995 11268 25007 11271
rect 23532 11240 25007 11268
rect 23532 11228 23538 11240
rect 24995 11237 25007 11240
rect 25041 11237 25053 11271
rect 27890 11268 27896 11280
rect 24995 11231 25053 11237
rect 27448 11240 27896 11268
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 22094 11200 22100 11212
rect 21324 11172 22100 11200
rect 21324 11160 21330 11172
rect 22094 11160 22100 11172
rect 22152 11160 22158 11212
rect 23198 11209 23204 11212
rect 23192 11163 23204 11209
rect 23256 11200 23262 11212
rect 24762 11200 24768 11212
rect 23256 11172 23292 11200
rect 24723 11172 24768 11200
rect 23198 11160 23204 11163
rect 23256 11160 23262 11172
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 25406 11200 25412 11212
rect 25367 11172 25412 11200
rect 25406 11160 25412 11172
rect 25464 11160 25470 11212
rect 25774 11160 25780 11212
rect 25832 11200 25838 11212
rect 25869 11203 25927 11209
rect 25869 11200 25881 11203
rect 25832 11172 25881 11200
rect 25832 11160 25838 11172
rect 25869 11169 25881 11172
rect 25915 11169 25927 11203
rect 25869 11163 25927 11169
rect 25958 11160 25964 11212
rect 26016 11200 26022 11212
rect 26053 11203 26111 11209
rect 26053 11200 26065 11203
rect 26016 11172 26065 11200
rect 26016 11160 26022 11172
rect 26053 11169 26065 11172
rect 26099 11169 26111 11203
rect 27338 11200 27344 11212
rect 27299 11172 27344 11200
rect 26053 11163 26111 11169
rect 27338 11160 27344 11172
rect 27396 11160 27402 11212
rect 27448 11209 27476 11240
rect 27890 11228 27896 11240
rect 27948 11228 27954 11280
rect 28261 11271 28319 11277
rect 28261 11237 28273 11271
rect 28307 11268 28319 11271
rect 28902 11268 28908 11280
rect 28307 11240 28908 11268
rect 28307 11237 28319 11240
rect 28261 11231 28319 11237
rect 28902 11228 28908 11240
rect 28960 11228 28966 11280
rect 31726 11268 31754 11308
rect 32320 11268 33120 11282
rect 31726 11240 33120 11268
rect 32320 11226 33120 11240
rect 27433 11203 27491 11209
rect 27433 11169 27445 11203
rect 27479 11169 27491 11203
rect 27614 11200 27620 11212
rect 27575 11172 27620 11200
rect 27433 11163 27491 11169
rect 27614 11160 27620 11172
rect 27672 11160 27678 11212
rect 27801 11203 27859 11209
rect 27801 11169 27813 11203
rect 27847 11200 27859 11203
rect 30466 11200 30472 11212
rect 27847 11172 30472 11200
rect 27847 11169 27859 11172
rect 27801 11163 27859 11169
rect 17460 11104 17632 11132
rect 17460 11092 17466 11104
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19337 11135 19395 11141
rect 19337 11132 19349 11135
rect 19208 11104 19349 11132
rect 19208 11092 19214 11104
rect 19337 11101 19349 11104
rect 19383 11101 19395 11135
rect 19337 11095 19395 11101
rect 22738 11092 22744 11144
rect 22796 11132 22802 11144
rect 22925 11135 22983 11141
rect 22925 11132 22937 11135
rect 22796 11104 22937 11132
rect 22796 11092 22802 11104
rect 22925 11101 22937 11104
rect 22971 11101 22983 11135
rect 27522 11132 27528 11144
rect 27483 11104 27528 11132
rect 22925 11095 22983 11101
rect 27522 11092 27528 11104
rect 27580 11092 27586 11144
rect 6411 11036 6592 11064
rect 14200 11036 14872 11064
rect 6411 11033 6423 11036
rect 6365 11027 6423 11033
rect 14200 11008 14228 11036
rect 25682 11024 25688 11076
rect 25740 11064 25746 11076
rect 27816 11064 27844 11163
rect 30466 11160 30472 11172
rect 30524 11160 30530 11212
rect 31110 11200 31116 11212
rect 31071 11172 31116 11200
rect 31110 11160 31116 11172
rect 31168 11160 31174 11212
rect 25740 11036 27844 11064
rect 25740 11024 25746 11036
rect 3936 10968 5120 10996
rect 3936 10956 3942 10968
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6549 10999 6607 11005
rect 6549 10996 6561 10999
rect 6052 10968 6561 10996
rect 6052 10956 6058 10968
rect 6549 10965 6561 10968
rect 6595 10965 6607 10999
rect 6549 10959 6607 10965
rect 14182 10956 14188 11008
rect 14240 10956 14246 11008
rect 14829 10999 14887 11005
rect 14829 10965 14841 10999
rect 14875 10996 14887 10999
rect 15838 10996 15844 11008
rect 14875 10968 15844 10996
rect 14875 10965 14887 10968
rect 14829 10959 14887 10965
rect 15838 10956 15844 10968
rect 15896 10996 15902 11008
rect 17402 10996 17408 11008
rect 15896 10968 17408 10996
rect 15896 10956 15902 10968
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 18138 10956 18144 11008
rect 18196 10996 18202 11008
rect 18877 10999 18935 11005
rect 18877 10996 18889 10999
rect 18196 10968 18889 10996
rect 18196 10956 18202 10968
rect 18877 10965 18889 10968
rect 18923 10965 18935 10999
rect 18877 10959 18935 10965
rect 24946 10956 24952 11008
rect 25004 10996 25010 11008
rect 25041 10999 25099 11005
rect 25041 10996 25053 10999
rect 25004 10968 25053 10996
rect 25004 10956 25010 10968
rect 25041 10965 25053 10968
rect 25087 10965 25099 10999
rect 25041 10959 25099 10965
rect 25130 10956 25136 11008
rect 25188 10996 25194 11008
rect 28902 10996 28908 11008
rect 25188 10968 28908 10996
rect 25188 10956 25194 10968
rect 28902 10956 28908 10968
rect 28960 10956 28966 11008
rect 29546 10996 29552 11008
rect 29507 10968 29552 10996
rect 29546 10956 29552 10968
rect 29604 10956 29610 11008
rect 1104 10906 32016 10928
rect 1104 10854 6102 10906
rect 6154 10854 6166 10906
rect 6218 10854 6230 10906
rect 6282 10854 6294 10906
rect 6346 10854 6358 10906
rect 6410 10854 16405 10906
rect 16457 10854 16469 10906
rect 16521 10854 16533 10906
rect 16585 10854 16597 10906
rect 16649 10854 16661 10906
rect 16713 10854 26709 10906
rect 26761 10854 26773 10906
rect 26825 10854 26837 10906
rect 26889 10854 26901 10906
rect 26953 10854 26965 10906
rect 27017 10854 32016 10906
rect 1104 10832 32016 10854
rect 2682 10752 2688 10804
rect 2740 10792 2746 10804
rect 3602 10792 3608 10804
rect 2740 10764 3608 10792
rect 2740 10752 2746 10764
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 3970 10792 3976 10804
rect 3931 10764 3976 10792
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5092 10764 5641 10792
rect 5092 10724 5120 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 10226 10792 10232 10804
rect 5868 10764 6040 10792
rect 5868 10752 5874 10764
rect 5902 10724 5908 10736
rect 1964 10696 5120 10724
rect 1964 10597 1992 10696
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 2961 10659 3019 10665
rect 2961 10656 2973 10659
rect 2924 10628 2973 10656
rect 2924 10616 2930 10628
rect 2961 10625 2973 10628
rect 3007 10625 3019 10659
rect 2961 10619 3019 10625
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 3200 10628 3249 10656
rect 3200 10616 3206 10628
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3970 10656 3976 10668
rect 3237 10619 3295 10625
rect 3804 10628 3976 10656
rect 3804 10597 3832 10628
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10656 4123 10659
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4111 10628 4537 10656
rect 4111 10625 4123 10628
rect 4065 10619 4123 10625
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 3936 10560 3981 10588
rect 3936 10548 3942 10560
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 4781 10591 4839 10597
rect 4781 10588 4793 10591
rect 4672 10560 4793 10588
rect 4672 10548 4678 10560
rect 4781 10557 4793 10560
rect 4827 10557 4839 10591
rect 4781 10551 4839 10557
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 5006 10591 5064 10597
rect 5006 10557 5018 10591
rect 5052 10588 5064 10591
rect 5092 10588 5120 10696
rect 5184 10696 5908 10724
rect 5184 10597 5212 10696
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5810 10656 5816 10668
rect 5675 10628 5816 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5810 10616 5816 10628
rect 5868 10656 5874 10668
rect 6012 10665 6040 10764
rect 7852 10764 10232 10792
rect 5997 10659 6055 10665
rect 5868 10628 5948 10656
rect 5868 10616 5874 10628
rect 5052 10560 5120 10588
rect 5169 10591 5227 10597
rect 5052 10557 5064 10560
rect 5006 10551 5064 10557
rect 5169 10557 5181 10591
rect 5215 10557 5227 10591
rect 5718 10588 5724 10600
rect 5679 10560 5724 10588
rect 5169 10551 5227 10557
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 4430 10520 4436 10532
rect 1903 10492 4436 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 4908 10520 4936 10551
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 5920 10597 5948 10628
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6914 10656 6920 10668
rect 6135 10628 6920 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 6012 10588 6040 10619
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 6178 10588 6184 10600
rect 6012 10560 6184 10588
rect 5905 10551 5963 10557
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6273 10591 6331 10597
rect 6273 10557 6285 10591
rect 6319 10588 6331 10591
rect 6546 10588 6552 10600
rect 6319 10560 6552 10588
rect 6319 10557 6331 10560
rect 6273 10551 6331 10557
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7852 10597 7880 10764
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 10597 10795 10655 10801
rect 10597 10761 10609 10795
rect 10643 10792 10655 10795
rect 10778 10792 10784 10804
rect 10643 10764 10784 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 18690 10792 18696 10804
rect 13780 10764 18696 10792
rect 13780 10752 13786 10764
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 19429 10795 19487 10801
rect 19429 10761 19441 10795
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10792 19671 10795
rect 19794 10792 19800 10804
rect 19659 10764 19800 10792
rect 19659 10761 19671 10764
rect 19613 10755 19671 10761
rect 9950 10724 9956 10736
rect 8036 10696 9956 10724
rect 8036 10665 8064 10696
rect 9950 10684 9956 10696
rect 10008 10724 10014 10736
rect 10410 10724 10416 10736
rect 10008 10696 10416 10724
rect 10008 10684 10014 10696
rect 10410 10684 10416 10696
rect 10468 10684 10474 10736
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 18230 10724 18236 10736
rect 17552 10696 18236 10724
rect 17552 10684 17558 10696
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 19444 10724 19472 10755
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 20438 10792 20444 10804
rect 19904 10764 20444 10792
rect 19904 10724 19932 10764
rect 20438 10752 20444 10764
rect 20496 10792 20502 10804
rect 20990 10792 20996 10804
rect 20496 10764 20996 10792
rect 20496 10752 20502 10764
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 21453 10795 21511 10801
rect 21453 10761 21465 10795
rect 21499 10792 21511 10795
rect 21910 10792 21916 10804
rect 21499 10764 21916 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 21910 10752 21916 10764
rect 21968 10752 21974 10804
rect 24486 10792 24492 10804
rect 24447 10764 24492 10792
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 27982 10752 27988 10804
rect 28040 10792 28046 10804
rect 28537 10795 28595 10801
rect 28537 10792 28549 10795
rect 28040 10764 28549 10792
rect 28040 10752 28046 10764
rect 28537 10761 28549 10764
rect 28583 10761 28595 10795
rect 28537 10755 28595 10761
rect 29730 10752 29736 10804
rect 29788 10792 29794 10804
rect 30929 10795 30987 10801
rect 30929 10792 30941 10795
rect 29788 10764 30941 10792
rect 29788 10752 29794 10764
rect 30929 10761 30941 10764
rect 30975 10761 30987 10795
rect 30929 10755 30987 10761
rect 19444 10696 19932 10724
rect 21082 10684 21088 10736
rect 21140 10724 21146 10736
rect 21358 10724 21364 10736
rect 21140 10696 21364 10724
rect 21140 10684 21146 10696
rect 21358 10684 21364 10696
rect 21416 10724 21422 10736
rect 21416 10696 26087 10724
rect 21416 10684 21422 10696
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 10134 10656 10140 10668
rect 8021 10619 8079 10625
rect 8220 10628 10140 10656
rect 8220 10597 8248 10628
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 11992 10628 14136 10656
rect 7101 10591 7159 10597
rect 7101 10588 7113 10591
rect 6880 10560 7113 10588
rect 6880 10548 6886 10560
rect 7101 10557 7113 10560
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10557 8171 10591
rect 8113 10551 8171 10557
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8846 10588 8852 10600
rect 8435 10560 8852 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8128 10520 8156 10551
rect 8846 10548 8852 10560
rect 8904 10588 8910 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 8904 10560 9505 10588
rect 8904 10548 8910 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9732 10560 9781 10588
rect 9732 10548 9738 10560
rect 9769 10557 9781 10560
rect 9815 10588 9827 10591
rect 10410 10588 10416 10600
rect 9815 10560 10416 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 10410 10548 10416 10560
rect 10468 10548 10474 10600
rect 11698 10548 11704 10600
rect 11756 10597 11762 10600
rect 11756 10588 11768 10597
rect 11756 10560 11801 10588
rect 11756 10551 11768 10560
rect 11756 10548 11762 10551
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 11992 10597 12020 10628
rect 14108 10600 14136 10628
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 18325 10659 18383 10665
rect 18325 10656 18337 10659
rect 17184 10628 18337 10656
rect 17184 10616 17190 10628
rect 18325 10625 18337 10628
rect 18371 10656 18383 10659
rect 19610 10656 19616 10668
rect 18371 10628 19616 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 20070 10656 20076 10668
rect 20031 10628 20076 10656
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 22002 10616 22008 10668
rect 22060 10656 22066 10668
rect 25498 10656 25504 10668
rect 22060 10628 25504 10656
rect 22060 10616 22066 10628
rect 25498 10616 25504 10628
rect 25556 10616 25562 10668
rect 11977 10591 12035 10597
rect 11977 10588 11989 10591
rect 11940 10560 11989 10588
rect 11940 10548 11946 10560
rect 11977 10557 11989 10560
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 9306 10520 9312 10532
rect 4908 10492 5120 10520
rect 8128 10492 9312 10520
rect 5092 10464 5120 10492
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 12452 10520 12480 10551
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12621 10591 12679 10597
rect 12621 10588 12633 10591
rect 12584 10560 12633 10588
rect 12584 10548 12590 10560
rect 12621 10557 12633 10560
rect 12667 10557 12679 10591
rect 12621 10551 12679 10557
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 13906 10588 13912 10600
rect 13587 10560 13912 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 14090 10588 14096 10600
rect 14003 10560 14096 10588
rect 14090 10548 14096 10560
rect 14148 10588 14154 10600
rect 14734 10588 14740 10600
rect 14148 10560 14740 10588
rect 14148 10548 14154 10560
rect 14734 10548 14740 10560
rect 14792 10588 14798 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 14792 10560 16129 10588
rect 14792 10548 14798 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 17954 10588 17960 10600
rect 17915 10560 17960 10588
rect 16117 10551 16175 10557
rect 17954 10548 17960 10560
rect 18012 10548 18018 10600
rect 18138 10588 18144 10600
rect 18099 10560 18144 10588
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10588 18291 10591
rect 18414 10588 18420 10600
rect 18279 10560 18420 10588
rect 18279 10557 18291 10560
rect 18233 10551 18291 10557
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 19334 10588 19340 10600
rect 18555 10560 19340 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 19334 10548 19340 10560
rect 19392 10548 19398 10600
rect 20088 10588 20116 10616
rect 20088 10560 22094 10588
rect 12802 10520 12808 10532
rect 12452 10492 12808 10520
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 14182 10520 14188 10532
rect 13412 10492 14188 10520
rect 13412 10480 13418 10492
rect 14182 10480 14188 10492
rect 14240 10480 14246 10532
rect 14366 10529 14372 10532
rect 14360 10483 14372 10529
rect 14424 10520 14430 10532
rect 14424 10492 14460 10520
rect 14366 10480 14372 10483
rect 14424 10480 14430 10492
rect 14550 10480 14556 10532
rect 14608 10520 14614 10532
rect 16384 10523 16442 10529
rect 14608 10492 15516 10520
rect 14608 10480 14614 10492
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5902 10452 5908 10464
rect 5132 10424 5908 10452
rect 5132 10412 5138 10424
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6454 10452 6460 10464
rect 6415 10424 6460 10452
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 7006 10452 7012 10464
rect 6788 10424 7012 10452
rect 6788 10412 6794 10424
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7650 10452 7656 10464
rect 7611 10424 7656 10452
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 12529 10455 12587 10461
rect 12529 10421 12541 10455
rect 12575 10452 12587 10455
rect 12986 10452 12992 10464
rect 12575 10424 12992 10452
rect 12575 10421 12587 10424
rect 12529 10415 12587 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13449 10455 13507 10461
rect 13449 10421 13461 10455
rect 13495 10452 13507 10455
rect 15102 10452 15108 10464
rect 13495 10424 15108 10452
rect 13495 10421 13507 10424
rect 13449 10415 13507 10421
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 15488 10461 15516 10492
rect 16384 10489 16396 10523
rect 16430 10520 16442 10523
rect 16758 10520 16764 10532
rect 16430 10492 16764 10520
rect 16430 10489 16442 10492
rect 16384 10483 16442 10489
rect 16758 10480 16764 10492
rect 16816 10480 16822 10532
rect 18156 10520 18184 10548
rect 19245 10523 19303 10529
rect 19245 10520 19257 10523
rect 18156 10492 19257 10520
rect 19245 10489 19257 10492
rect 19291 10489 19303 10523
rect 19245 10483 19303 10489
rect 19461 10523 19519 10529
rect 19461 10489 19473 10523
rect 19507 10520 19519 10523
rect 19794 10520 19800 10532
rect 19507 10492 19800 10520
rect 19507 10489 19519 10492
rect 19461 10483 19519 10489
rect 19794 10480 19800 10492
rect 19852 10480 19858 10532
rect 20346 10529 20352 10532
rect 20340 10483 20352 10529
rect 20404 10520 20410 10532
rect 22066 10520 22094 10560
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22244 10560 22293 10588
rect 22244 10548 22250 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22462 10588 22468 10600
rect 22423 10560 22468 10588
rect 22281 10551 22339 10557
rect 22462 10548 22468 10560
rect 22520 10548 22526 10600
rect 22554 10548 22560 10600
rect 22612 10588 22618 10600
rect 23106 10588 23112 10600
rect 22612 10560 22657 10588
rect 23067 10560 23112 10588
rect 22612 10548 22618 10560
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 23293 10591 23351 10597
rect 23293 10557 23305 10591
rect 23339 10588 23351 10591
rect 23474 10588 23480 10600
rect 23339 10560 23480 10588
rect 23339 10557 23351 10560
rect 23293 10551 23351 10557
rect 23474 10548 23480 10560
rect 23532 10548 23538 10600
rect 24578 10548 24584 10600
rect 24636 10588 24642 10600
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24636 10560 25145 10588
rect 24636 10548 24642 10560
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 22738 10520 22744 10532
rect 20404 10492 20440 10520
rect 22066 10492 22744 10520
rect 20346 10480 20352 10483
rect 20404 10480 20410 10492
rect 22738 10480 22744 10492
rect 22796 10480 22802 10532
rect 24026 10480 24032 10532
rect 24084 10520 24090 10532
rect 24949 10523 25007 10529
rect 24949 10520 24961 10523
rect 24084 10492 24961 10520
rect 24084 10480 24090 10492
rect 24949 10489 24961 10492
rect 24995 10520 25007 10523
rect 25777 10523 25835 10529
rect 25777 10520 25789 10523
rect 24995 10492 25789 10520
rect 24995 10489 25007 10492
rect 24949 10483 25007 10489
rect 25777 10489 25789 10492
rect 25823 10489 25835 10523
rect 25958 10520 25964 10532
rect 25919 10492 25964 10520
rect 25777 10483 25835 10489
rect 25958 10480 25964 10492
rect 26016 10480 26022 10532
rect 26059 10520 26087 10696
rect 26510 10616 26516 10668
rect 26568 10656 26574 10668
rect 27249 10659 27307 10665
rect 26568 10628 26832 10656
rect 26568 10616 26574 10628
rect 26602 10588 26608 10600
rect 26563 10560 26608 10588
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 26804 10597 26832 10628
rect 27249 10625 27261 10659
rect 27295 10656 27307 10659
rect 28000 10656 28028 10752
rect 27295 10628 28028 10656
rect 27295 10625 27307 10628
rect 27249 10619 27307 10625
rect 26789 10591 26847 10597
rect 26789 10557 26801 10591
rect 26835 10557 26847 10591
rect 26789 10551 26847 10557
rect 27430 10548 27436 10600
rect 27488 10588 27494 10600
rect 27525 10591 27583 10597
rect 27525 10588 27537 10591
rect 27488 10560 27537 10588
rect 27488 10548 27494 10560
rect 27525 10557 27537 10560
rect 27571 10557 27583 10591
rect 29546 10588 29552 10600
rect 29507 10560 29552 10588
rect 27525 10551 27583 10557
rect 29546 10548 29552 10560
rect 29604 10548 29610 10600
rect 29638 10548 29644 10600
rect 29696 10588 29702 10600
rect 29805 10591 29863 10597
rect 29805 10588 29817 10591
rect 29696 10560 29817 10588
rect 29696 10548 29702 10560
rect 29805 10557 29817 10560
rect 29851 10557 29863 10591
rect 29805 10551 29863 10557
rect 28166 10520 28172 10532
rect 26059 10492 28172 10520
rect 28166 10480 28172 10492
rect 28224 10480 28230 10532
rect 15473 10455 15531 10461
rect 15473 10421 15485 10455
rect 15519 10421 15531 10455
rect 17494 10452 17500 10464
rect 17455 10424 17500 10452
rect 15473 10415 15531 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 18690 10452 18696 10464
rect 18651 10424 18696 10452
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 22097 10455 22155 10461
rect 22097 10421 22109 10455
rect 22143 10452 22155 10455
rect 22370 10452 22376 10464
rect 22143 10424 22376 10452
rect 22143 10421 22155 10424
rect 22097 10415 22155 10421
rect 22370 10412 22376 10424
rect 22428 10412 22434 10464
rect 23382 10412 23388 10464
rect 23440 10452 23446 10464
rect 23477 10455 23535 10461
rect 23477 10452 23489 10455
rect 23440 10424 23489 10452
rect 23440 10412 23446 10424
rect 23477 10421 23489 10424
rect 23523 10421 23535 10455
rect 23477 10415 23535 10421
rect 25317 10455 25375 10461
rect 25317 10421 25329 10455
rect 25363 10452 25375 10455
rect 25682 10452 25688 10464
rect 25363 10424 25688 10452
rect 25363 10421 25375 10424
rect 25317 10415 25375 10421
rect 25682 10412 25688 10424
rect 25740 10412 25746 10464
rect 26142 10452 26148 10464
rect 26103 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 26697 10455 26755 10461
rect 26697 10421 26709 10455
rect 26743 10452 26755 10455
rect 28718 10452 28724 10464
rect 26743 10424 28724 10452
rect 26743 10421 26755 10424
rect 26697 10415 26755 10421
rect 28718 10412 28724 10424
rect 28776 10412 28782 10464
rect 1104 10362 32016 10384
rect 1104 10310 11253 10362
rect 11305 10310 11317 10362
rect 11369 10310 11381 10362
rect 11433 10310 11445 10362
rect 11497 10310 11509 10362
rect 11561 10310 21557 10362
rect 21609 10310 21621 10362
rect 21673 10310 21685 10362
rect 21737 10310 21749 10362
rect 21801 10310 21813 10362
rect 21865 10310 32016 10362
rect 1104 10288 32016 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2096 10220 2421 10248
rect 2096 10208 2102 10220
rect 2409 10217 2421 10220
rect 2455 10248 2467 10251
rect 2682 10248 2688 10260
rect 2455 10220 2688 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5408 10220 5457 10248
rect 5408 10208 5414 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7745 10251 7803 10257
rect 7745 10248 7757 10251
rect 6880 10220 7757 10248
rect 6880 10208 6886 10220
rect 7745 10217 7757 10220
rect 7791 10217 7803 10251
rect 8478 10248 8484 10260
rect 8439 10220 8484 10248
rect 7745 10211 7803 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 10284 10220 10333 10248
rect 10284 10208 10290 10220
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 10321 10211 10379 10217
rect 2958 10140 2964 10192
rect 3016 10180 3022 10192
rect 3522 10183 3580 10189
rect 3522 10180 3534 10183
rect 3016 10152 3534 10180
rect 3016 10140 3022 10152
rect 3522 10149 3534 10152
rect 3568 10149 3580 10183
rect 3522 10143 3580 10149
rect 4632 10152 5488 10180
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 3200 10084 4537 10112
rect 3200 10072 3206 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 3786 10004 3792 10056
rect 3844 10044 3850 10056
rect 4632 10044 4660 10152
rect 5460 10124 5488 10152
rect 6454 10140 6460 10192
rect 6512 10180 6518 10192
rect 6610 10183 6668 10189
rect 6610 10180 6622 10183
rect 6512 10152 6622 10180
rect 6512 10140 6518 10152
rect 6610 10149 6622 10152
rect 6656 10149 6668 10183
rect 6610 10143 6668 10149
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 9186 10183 9244 10189
rect 9186 10180 9198 10183
rect 7708 10152 9198 10180
rect 7708 10140 7714 10152
rect 9186 10149 9198 10152
rect 9232 10149 9244 10183
rect 9186 10143 9244 10149
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 5350 10112 5356 10124
rect 4764 10084 5356 10112
rect 4764 10072 4770 10084
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 5500 10084 6377 10112
rect 5500 10072 5506 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 10336 10112 10364 10211
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 10468 10220 13001 10248
rect 10468 10208 10474 10220
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 12989 10211 13047 10217
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 14366 10248 14372 10260
rect 14323 10220 14372 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 18046 10248 18052 10260
rect 17552 10220 18052 10248
rect 17552 10208 17558 10220
rect 18046 10208 18052 10220
rect 18104 10248 18110 10260
rect 19426 10248 19432 10260
rect 18104 10220 19288 10248
rect 19387 10220 19432 10248
rect 18104 10208 18110 10220
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12345 10183 12403 10189
rect 12345 10180 12357 10183
rect 11940 10152 12357 10180
rect 11940 10140 11946 10152
rect 12345 10149 12357 10152
rect 12391 10180 12403 10183
rect 12618 10180 12624 10192
rect 12391 10152 12624 10180
rect 12391 10149 12403 10152
rect 12345 10143 12403 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 19150 10180 19156 10192
rect 18064 10152 19156 10180
rect 10781 10115 10839 10121
rect 10781 10112 10793 10115
rect 10336 10084 10793 10112
rect 6365 10075 6423 10081
rect 10781 10081 10793 10084
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 3844 10016 4660 10044
rect 5261 10047 5319 10053
rect 3844 10004 3850 10016
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 1949 9911 2007 9917
rect 1949 9877 1961 9911
rect 1995 9908 2007 9911
rect 2130 9908 2136 9920
rect 1995 9880 2136 9908
rect 1995 9877 2007 9880
rect 1949 9871 2007 9877
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 4433 9911 4491 9917
rect 4433 9877 4445 9911
rect 4479 9908 4491 9911
rect 4706 9908 4712 9920
rect 4479 9880 4712 9908
rect 4479 9877 4491 9880
rect 4433 9871 4491 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 5276 9908 5304 10007
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 7708 10016 8953 10044
rect 7708 10004 7714 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 11808 9976 11836 10075
rect 12710 10072 12716 10124
rect 12768 10112 12774 10124
rect 13078 10112 13084 10124
rect 12768 10084 13084 10112
rect 12768 10072 12774 10084
rect 13078 10072 13084 10084
rect 13136 10112 13142 10124
rect 13541 10115 13599 10121
rect 13541 10112 13553 10115
rect 13136 10084 13553 10112
rect 13136 10072 13142 10084
rect 13541 10081 13553 10084
rect 13587 10081 13599 10115
rect 13722 10112 13728 10124
rect 13683 10084 13728 10112
rect 13541 10075 13599 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 13872 10084 13917 10112
rect 13872 10072 13878 10084
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 14056 10084 14105 10112
rect 14056 10072 14062 10084
rect 14093 10081 14105 10084
rect 14139 10112 14151 10115
rect 14550 10112 14556 10124
rect 14139 10084 14556 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14826 10072 14832 10124
rect 14884 10112 14890 10124
rect 18064 10121 18092 10152
rect 19150 10140 19156 10152
rect 19208 10140 19214 10192
rect 19260 10180 19288 10220
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 20257 10251 20315 10257
rect 20257 10217 20269 10251
rect 20303 10248 20315 10251
rect 20346 10248 20352 10260
rect 20303 10220 20352 10248
rect 20303 10217 20315 10220
rect 20257 10211 20315 10217
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22278 10248 22284 10260
rect 21968 10220 22284 10248
rect 21968 10208 21974 10220
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 23198 10248 23204 10260
rect 23159 10220 23204 10248
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 30742 10248 30748 10260
rect 23308 10220 30748 10248
rect 19260 10152 20760 10180
rect 14993 10115 15051 10121
rect 14993 10112 15005 10115
rect 14884 10084 15005 10112
rect 14884 10072 14890 10084
rect 14993 10081 15005 10084
rect 15039 10081 15051 10115
rect 14993 10075 15051 10081
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 18316 10115 18374 10121
rect 18316 10081 18328 10115
rect 18362 10112 18374 10115
rect 18690 10112 18696 10124
rect 18362 10084 18696 10112
rect 18362 10081 18374 10084
rect 18316 10075 18374 10081
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 19886 10072 19892 10124
rect 19944 10112 19950 10124
rect 20732 10121 20760 10152
rect 20806 10140 20812 10192
rect 20864 10180 20870 10192
rect 23308 10180 23336 10220
rect 30742 10208 30748 10220
rect 30800 10208 30806 10260
rect 30926 10248 30932 10260
rect 30887 10220 30932 10248
rect 30926 10208 30932 10220
rect 30984 10208 30990 10260
rect 20864 10152 23336 10180
rect 20864 10140 20870 10152
rect 24578 10140 24584 10192
rect 24636 10180 24642 10192
rect 24857 10183 24915 10189
rect 24857 10180 24869 10183
rect 24636 10152 24869 10180
rect 24636 10140 24642 10152
rect 24857 10149 24869 10152
rect 24903 10149 24915 10183
rect 29270 10180 29276 10192
rect 24857 10143 24915 10149
rect 25424 10152 29276 10180
rect 20073 10115 20131 10121
rect 20073 10112 20085 10115
rect 19944 10084 20085 10112
rect 19944 10072 19950 10084
rect 20073 10081 20085 10084
rect 20119 10081 20131 10115
rect 20073 10075 20131 10081
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 21450 10072 21456 10124
rect 21508 10112 21514 10124
rect 21726 10112 21732 10124
rect 21508 10084 21732 10112
rect 21508 10072 21514 10084
rect 21726 10072 21732 10084
rect 21784 10112 21790 10124
rect 22005 10115 22063 10121
rect 22005 10112 22017 10115
rect 21784 10084 22017 10112
rect 21784 10072 21790 10084
rect 22005 10081 22017 10084
rect 22051 10081 22063 10115
rect 22278 10112 22284 10124
rect 22239 10084 22284 10112
rect 22005 10075 22063 10081
rect 22278 10072 22284 10084
rect 22336 10072 22342 10124
rect 22370 10072 22376 10124
rect 22428 10112 22434 10124
rect 22465 10115 22523 10121
rect 22465 10112 22477 10115
rect 22428 10084 22477 10112
rect 22428 10072 22434 10084
rect 22465 10081 22477 10084
rect 22511 10081 22523 10115
rect 23382 10112 23388 10124
rect 23343 10084 23388 10112
rect 22465 10075 22523 10081
rect 23382 10072 23388 10084
rect 23440 10072 23446 10124
rect 24026 10112 24032 10124
rect 23987 10084 24032 10112
rect 24026 10072 24032 10084
rect 24084 10072 24090 10124
rect 24121 10115 24179 10121
rect 24121 10081 24133 10115
rect 24167 10112 24179 10115
rect 24673 10115 24731 10121
rect 24673 10112 24685 10115
rect 24167 10084 24685 10112
rect 24167 10081 24179 10084
rect 24121 10075 24179 10081
rect 24673 10081 24685 10084
rect 24719 10081 24731 10115
rect 24673 10075 24731 10081
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 13909 10047 13967 10053
rect 13909 10044 13921 10047
rect 12575 10016 13921 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 13909 10013 13921 10016
rect 13955 10044 13967 10047
rect 14366 10044 14372 10056
rect 13955 10016 14372 10044
rect 13955 10013 13967 10016
rect 13909 10007 13967 10013
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14734 10044 14740 10056
rect 14647 10016 14740 10044
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 16022 10004 16028 10056
rect 16080 10044 16086 10056
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 16080 10016 17233 10044
rect 16080 10004 16086 10016
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 17586 10044 17592 10056
rect 17543 10016 17592 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10044 22247 10047
rect 23014 10044 23020 10056
rect 22235 10016 23020 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 14090 9976 14096 9988
rect 11808 9948 14096 9976
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 5626 9908 5632 9920
rect 5276 9880 5632 9908
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 5813 9911 5871 9917
rect 5813 9877 5825 9911
rect 5859 9908 5871 9911
rect 7834 9908 7840 9920
rect 5859 9880 7840 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 11146 9908 11152 9920
rect 10919 9880 11152 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 11698 9908 11704 9920
rect 11659 9880 11704 9908
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 12618 9868 12624 9920
rect 12676 9908 12682 9920
rect 12802 9908 12808 9920
rect 12676 9880 12808 9908
rect 12676 9868 12682 9880
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 14752 9908 14780 10004
rect 22094 9936 22100 9988
rect 22152 9976 22158 9988
rect 24044 9976 24072 10072
rect 24688 10044 24716 10075
rect 25314 10044 25320 10056
rect 24688 10016 25320 10044
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 25424 9976 25452 10152
rect 29270 10140 29276 10152
rect 29328 10140 29334 10192
rect 29816 10183 29874 10189
rect 29816 10149 29828 10183
rect 29862 10180 29874 10183
rect 30282 10180 30288 10192
rect 29862 10152 30288 10180
rect 29862 10149 29874 10152
rect 29816 10143 29874 10149
rect 30282 10140 30288 10152
rect 30340 10140 30346 10192
rect 25501 10115 25559 10121
rect 25501 10081 25513 10115
rect 25547 10081 25559 10115
rect 25501 10075 25559 10081
rect 25869 10115 25927 10121
rect 25869 10081 25881 10115
rect 25915 10112 25927 10115
rect 25958 10112 25964 10124
rect 25915 10084 25964 10112
rect 25915 10081 25927 10084
rect 25869 10075 25927 10081
rect 22152 9948 22197 9976
rect 24044 9948 25452 9976
rect 25516 9976 25544 10075
rect 25958 10072 25964 10084
rect 26016 10072 26022 10124
rect 27338 10072 27344 10124
rect 27396 10112 27402 10124
rect 28086 10115 28144 10121
rect 28086 10112 28098 10115
rect 27396 10084 28098 10112
rect 27396 10072 27402 10084
rect 28086 10081 28098 10084
rect 28132 10081 28144 10115
rect 28086 10075 28144 10081
rect 28353 10047 28411 10053
rect 28353 10013 28365 10047
rect 28399 10044 28411 10047
rect 28994 10044 29000 10056
rect 28399 10016 29000 10044
rect 28399 10013 28411 10016
rect 28353 10007 28411 10013
rect 28994 10004 29000 10016
rect 29052 10044 29058 10056
rect 29546 10044 29552 10056
rect 29052 10016 29552 10044
rect 29052 10004 29058 10016
rect 29546 10004 29552 10016
rect 29604 10004 29610 10056
rect 26602 9976 26608 9988
rect 25516 9948 26608 9976
rect 22152 9936 22158 9948
rect 15746 9908 15752 9920
rect 14752 9880 15752 9908
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 16114 9908 16120 9920
rect 16075 9880 16120 9908
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16850 9868 16856 9920
rect 16908 9908 16914 9920
rect 20809 9911 20867 9917
rect 20809 9908 20821 9911
rect 16908 9880 20821 9908
rect 16908 9868 16914 9880
rect 20809 9877 20821 9880
rect 20855 9877 20867 9911
rect 21818 9908 21824 9920
rect 21779 9880 21824 9908
rect 20809 9871 20867 9877
rect 21818 9868 21824 9880
rect 21876 9868 21882 9920
rect 25038 9908 25044 9920
rect 24999 9880 25044 9908
rect 25038 9868 25044 9880
rect 25096 9868 25102 9920
rect 25424 9908 25452 9948
rect 26602 9936 26608 9948
rect 26660 9976 26666 9988
rect 26973 9979 27031 9985
rect 26973 9976 26985 9979
rect 26660 9948 26985 9976
rect 26660 9936 26666 9948
rect 26973 9945 26985 9948
rect 27019 9945 27031 9979
rect 26973 9939 27031 9945
rect 25593 9911 25651 9917
rect 25593 9908 25605 9911
rect 25424 9880 25605 9908
rect 25593 9877 25605 9880
rect 25639 9877 25651 9911
rect 25593 9871 25651 9877
rect 26053 9911 26111 9917
rect 26053 9877 26065 9911
rect 26099 9908 26111 9911
rect 26418 9908 26424 9920
rect 26099 9880 26424 9908
rect 26099 9877 26111 9880
rect 26053 9871 26111 9877
rect 26418 9868 26424 9880
rect 26476 9868 26482 9920
rect 27614 9868 27620 9920
rect 27672 9908 27678 9920
rect 28813 9911 28871 9917
rect 28813 9908 28825 9911
rect 27672 9880 28825 9908
rect 27672 9868 27678 9880
rect 28813 9877 28825 9880
rect 28859 9877 28871 9911
rect 28813 9871 28871 9877
rect 1104 9818 32016 9840
rect 1104 9766 6102 9818
rect 6154 9766 6166 9818
rect 6218 9766 6230 9818
rect 6282 9766 6294 9818
rect 6346 9766 6358 9818
rect 6410 9766 16405 9818
rect 16457 9766 16469 9818
rect 16521 9766 16533 9818
rect 16585 9766 16597 9818
rect 16649 9766 16661 9818
rect 16713 9766 26709 9818
rect 26761 9766 26773 9818
rect 26825 9766 26837 9818
rect 26889 9766 26901 9818
rect 26953 9766 26965 9818
rect 27017 9766 32016 9818
rect 1104 9744 32016 9766
rect 3326 9664 3332 9716
rect 3384 9704 3390 9716
rect 3878 9704 3884 9716
rect 3384 9676 3884 9704
rect 3384 9664 3390 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 7006 9704 7012 9716
rect 4672 9676 7012 9704
rect 4672 9664 4678 9676
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 14826 9704 14832 9716
rect 14787 9676 14832 9704
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 22094 9664 22100 9716
rect 22152 9704 22158 9716
rect 22741 9707 22799 9713
rect 22741 9704 22753 9707
rect 22152 9676 22753 9704
rect 22152 9664 22158 9676
rect 22741 9673 22753 9676
rect 22787 9673 22799 9707
rect 23566 9704 23572 9716
rect 23479 9676 23572 9704
rect 22741 9667 22799 9673
rect 23566 9664 23572 9676
rect 23624 9704 23630 9716
rect 24486 9704 24492 9716
rect 23624 9676 24492 9704
rect 23624 9664 23630 9676
rect 24486 9664 24492 9676
rect 24544 9664 24550 9716
rect 27246 9664 27252 9716
rect 27304 9704 27310 9716
rect 30006 9704 30012 9716
rect 27304 9676 30012 9704
rect 27304 9664 27310 9676
rect 30006 9664 30012 9676
rect 30064 9664 30070 9716
rect 4522 9596 4528 9648
rect 4580 9596 4586 9648
rect 4893 9639 4951 9645
rect 4893 9605 4905 9639
rect 4939 9636 4951 9639
rect 4982 9636 4988 9648
rect 4939 9608 4988 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 5445 9639 5503 9645
rect 5445 9605 5457 9639
rect 5491 9636 5503 9639
rect 5994 9636 6000 9648
rect 5491 9608 6000 9636
rect 5491 9605 5503 9608
rect 5445 9599 5503 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 7374 9636 7380 9648
rect 7335 9608 7380 9636
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 10318 9596 10324 9648
rect 10376 9636 10382 9648
rect 10413 9639 10471 9645
rect 10413 9636 10425 9639
rect 10376 9608 10425 9636
rect 10376 9596 10382 9608
rect 10413 9605 10425 9608
rect 10459 9605 10471 9639
rect 10413 9599 10471 9605
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 13170 9636 13176 9648
rect 12492 9608 12537 9636
rect 12820 9608 13176 9636
rect 12492 9596 12498 9608
rect 2498 9460 2504 9512
rect 2556 9509 2562 9512
rect 2556 9500 2568 9509
rect 2777 9503 2835 9509
rect 2556 9472 2601 9500
rect 2556 9463 2568 9472
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 3786 9500 3792 9512
rect 2823 9472 3792 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 2556 9460 2562 9463
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 4246 9500 4252 9512
rect 4207 9472 4252 9500
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4430 9500 4436 9512
rect 4391 9472 4436 9500
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 4540 9509 4568 9596
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 8386 9528 8392 9580
rect 8444 9568 8450 9580
rect 12710 9568 12716 9580
rect 8444 9540 12716 9568
rect 8444 9528 8450 9540
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 4528 9503 4586 9509
rect 4528 9469 4540 9503
rect 4574 9469 4586 9503
rect 4528 9463 4586 9469
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 4672 9472 4717 9500
rect 4672 9460 4678 9472
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5684 9472 6101 9500
rect 5684 9460 5690 9472
rect 6089 9469 6101 9472
rect 6135 9500 6147 9503
rect 6840 9500 6868 9528
rect 6135 9472 6868 9500
rect 8297 9503 8355 9509
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 8297 9469 8309 9503
rect 8343 9500 8355 9503
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 8343 9472 9045 9500
rect 8343 9469 8355 9472
rect 8297 9463 8355 9469
rect 9033 9469 9045 9472
rect 9079 9500 9091 9503
rect 9122 9500 9128 9512
rect 9079 9472 9128 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9306 9500 9312 9512
rect 9267 9472 9312 9500
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 11609 9503 11667 9509
rect 11609 9469 11621 9503
rect 11655 9500 11667 9503
rect 12820 9500 12848 9608
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 15010 9596 15016 9648
rect 15068 9596 15074 9648
rect 15562 9596 15568 9648
rect 15620 9596 15626 9648
rect 16758 9636 16764 9648
rect 16719 9608 16764 9636
rect 16758 9596 16764 9608
rect 16816 9596 16822 9648
rect 17954 9636 17960 9648
rect 17915 9608 17960 9636
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 20165 9639 20223 9645
rect 20165 9636 20177 9639
rect 19392 9608 20177 9636
rect 19392 9596 19398 9608
rect 20165 9605 20177 9608
rect 20211 9605 20223 9639
rect 22186 9636 22192 9648
rect 22147 9608 22192 9636
rect 20165 9599 20223 9605
rect 22186 9596 22192 9608
rect 22244 9596 22250 9648
rect 30098 9636 30104 9648
rect 30059 9608 30104 9636
rect 30098 9596 30104 9608
rect 30156 9596 30162 9648
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 15028 9568 15056 9596
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 15028 9540 15301 9568
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15580 9568 15608 9596
rect 15289 9531 15347 9537
rect 15488 9540 15608 9568
rect 11655 9472 12848 9500
rect 11655 9469 11667 9472
rect 11609 9463 11667 9469
rect 12894 9460 12900 9512
rect 12952 9500 12958 9512
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 12952 9472 14105 9500
rect 12952 9460 12958 9472
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9469 15071 9503
rect 15197 9503 15255 9509
rect 15197 9490 15209 9503
rect 15243 9490 15255 9503
rect 15013 9463 15071 9469
rect 4264 9432 4292 9460
rect 4890 9432 4896 9444
rect 4264 9404 4896 9432
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 6546 9432 6552 9444
rect 6012 9404 6552 9432
rect 1397 9367 1455 9373
rect 1397 9333 1409 9367
rect 1443 9364 1455 9367
rect 2222 9364 2228 9376
rect 1443 9336 2228 9364
rect 1443 9333 1455 9336
rect 1397 9327 1455 9333
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 6012 9373 6040 9404
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 6825 9435 6883 9441
rect 6825 9401 6837 9435
rect 6871 9432 6883 9435
rect 7374 9432 7380 9444
rect 6871 9404 7380 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 11425 9435 11483 9441
rect 11425 9401 11437 9435
rect 11471 9432 11483 9435
rect 12805 9435 12863 9441
rect 11471 9404 11652 9432
rect 11471 9401 11483 9404
rect 11425 9395 11483 9401
rect 11624 9376 11652 9404
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 14369 9435 14427 9441
rect 14369 9432 14381 9435
rect 12851 9404 14381 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 14369 9401 14381 9404
rect 14415 9401 14427 9435
rect 14369 9395 14427 9401
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5684 9336 6009 9364
rect 5684 9324 5690 9336
rect 5997 9333 6009 9336
rect 6043 9333 6055 9367
rect 5997 9327 6055 9333
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6420 9336 6745 9364
rect 6420 9324 6426 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 11020 9336 11253 9364
rect 11020 9324 11026 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 11606 9324 11612 9376
rect 11664 9324 11670 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 13998 9364 14004 9376
rect 12943 9336 14004 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 15028 9364 15056 9463
rect 15194 9438 15200 9490
rect 15252 9438 15258 9490
rect 15304 9444 15332 9531
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9500 15439 9503
rect 15488 9500 15516 9540
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16172 9540 20116 9568
rect 16172 9528 16178 9540
rect 15427 9472 15516 9500
rect 15565 9503 15623 9509
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15654 9500 15660 9512
rect 15611 9472 15660 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 15654 9460 15660 9472
rect 15712 9500 15718 9512
rect 16022 9500 16028 9512
rect 15712 9472 16028 9500
rect 15712 9460 15718 9472
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 16224 9509 16252 9540
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 16301 9503 16359 9509
rect 16301 9469 16313 9503
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 16577 9503 16635 9509
rect 16577 9469 16589 9503
rect 16623 9500 16635 9503
rect 17494 9500 17500 9512
rect 16623 9472 17500 9500
rect 16623 9469 16635 9472
rect 16577 9463 16635 9469
rect 15286 9392 15292 9444
rect 15344 9432 15350 9444
rect 16316 9432 16344 9463
rect 15344 9404 16344 9432
rect 16408 9432 16436 9463
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 19621 9503 19679 9509
rect 18064 9472 19334 9500
rect 17126 9432 17132 9444
rect 16408 9404 17132 9432
rect 15344 9392 15350 9404
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 17313 9435 17371 9441
rect 17313 9401 17325 9435
rect 17359 9432 17371 9435
rect 18064 9432 18092 9472
rect 17359 9404 18092 9432
rect 18141 9435 18199 9441
rect 17359 9401 17371 9404
rect 17313 9395 17371 9401
rect 18141 9401 18153 9435
rect 18187 9401 18199 9435
rect 19306 9432 19334 9472
rect 19621 9469 19633 9503
rect 19667 9500 19679 9503
rect 19886 9500 19892 9512
rect 19667 9472 19892 9500
rect 19667 9469 19679 9472
rect 19621 9463 19679 9469
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 20088 9509 20116 9540
rect 21818 9528 21824 9580
rect 21876 9528 21882 9580
rect 22002 9568 22008 9580
rect 21928 9540 22008 9568
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 20809 9503 20867 9509
rect 20809 9500 20821 9503
rect 20496 9472 20821 9500
rect 20496 9460 20502 9472
rect 20809 9469 20821 9472
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 21076 9503 21134 9509
rect 21076 9469 21088 9503
rect 21122 9500 21134 9503
rect 21836 9500 21864 9528
rect 21122 9472 21864 9500
rect 21122 9469 21134 9472
rect 21076 9463 21134 9469
rect 21928 9432 21956 9540
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 24765 9571 24823 9577
rect 24765 9537 24777 9571
rect 24811 9568 24823 9571
rect 26697 9571 26755 9577
rect 24811 9540 25544 9568
rect 24811 9537 24823 9540
rect 24765 9531 24823 9537
rect 22554 9460 22560 9512
rect 22612 9500 22618 9512
rect 22833 9503 22891 9509
rect 22833 9500 22845 9503
rect 22612 9472 22845 9500
rect 22612 9460 22618 9472
rect 22833 9469 22845 9472
rect 22879 9500 22891 9503
rect 24026 9500 24032 9512
rect 22879 9472 24032 9500
rect 22879 9469 22891 9472
rect 22833 9463 22891 9469
rect 24026 9460 24032 9472
rect 24084 9460 24090 9512
rect 24578 9460 24584 9512
rect 24636 9500 24642 9512
rect 24673 9503 24731 9509
rect 24673 9500 24685 9503
rect 24636 9472 24685 9500
rect 24636 9460 24642 9472
rect 24673 9469 24685 9472
rect 24719 9469 24731 9503
rect 25314 9500 25320 9512
rect 25275 9472 25320 9500
rect 24673 9463 24731 9469
rect 25314 9460 25320 9472
rect 25372 9460 25378 9512
rect 25516 9509 25544 9540
rect 26697 9537 26709 9571
rect 26743 9568 26755 9571
rect 27430 9568 27436 9580
rect 26743 9540 27436 9568
rect 26743 9537 26755 9540
rect 26697 9531 26755 9537
rect 27430 9528 27436 9540
rect 27488 9528 27494 9580
rect 25501 9503 25559 9509
rect 25501 9469 25513 9503
rect 25547 9500 25559 9503
rect 25958 9500 25964 9512
rect 25547 9472 25964 9500
rect 25547 9469 25559 9472
rect 25501 9463 25559 9469
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 26421 9503 26479 9509
rect 26421 9469 26433 9503
rect 26467 9500 26479 9503
rect 26510 9500 26516 9512
rect 26467 9472 26516 9500
rect 26467 9469 26479 9472
rect 26421 9463 26479 9469
rect 26510 9460 26516 9472
rect 26568 9460 26574 9512
rect 26602 9460 26608 9512
rect 26660 9500 26666 9512
rect 26789 9503 26847 9509
rect 26660 9472 26705 9500
rect 26660 9460 26666 9472
rect 26789 9469 26801 9503
rect 26835 9469 26847 9503
rect 26789 9463 26847 9469
rect 26973 9503 27031 9509
rect 26973 9469 26985 9503
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 24854 9432 24860 9444
rect 19306 9404 21956 9432
rect 22103 9404 24860 9432
rect 18141 9395 18199 9401
rect 16114 9364 16120 9376
rect 15028 9336 16120 9364
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16942 9364 16948 9376
rect 16356 9336 16948 9364
rect 16356 9324 16362 9336
rect 16942 9324 16948 9336
rect 17000 9364 17006 9376
rect 17328 9364 17356 9395
rect 17000 9336 17356 9364
rect 17405 9367 17463 9373
rect 17000 9324 17006 9336
rect 17405 9333 17417 9367
rect 17451 9364 17463 9367
rect 17494 9364 17500 9376
rect 17451 9336 17500 9364
rect 17451 9333 17463 9336
rect 17405 9327 17463 9333
rect 17494 9324 17500 9336
rect 17552 9364 17558 9376
rect 18156 9364 18184 9395
rect 19426 9364 19432 9376
rect 17552 9336 18184 9364
rect 19387 9336 19432 9364
rect 17552 9324 17558 9336
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 22103 9364 22131 9404
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 25685 9435 25743 9441
rect 25685 9401 25697 9435
rect 25731 9401 25743 9435
rect 25685 9395 25743 9401
rect 20312 9336 22131 9364
rect 25700 9364 25728 9395
rect 26234 9392 26240 9444
rect 26292 9432 26298 9444
rect 26804 9432 26832 9463
rect 26878 9432 26884 9444
rect 26292 9404 26884 9432
rect 26292 9392 26298 9404
rect 26878 9392 26884 9404
rect 26936 9392 26942 9444
rect 26694 9364 26700 9376
rect 25700 9336 26700 9364
rect 20312 9324 20318 9336
rect 26694 9324 26700 9336
rect 26752 9324 26758 9376
rect 26988 9364 27016 9463
rect 27522 9460 27528 9512
rect 27580 9500 27586 9512
rect 28994 9500 29000 9512
rect 27580 9472 28856 9500
rect 28955 9472 29000 9500
rect 27580 9460 27586 9472
rect 27157 9435 27215 9441
rect 27157 9401 27169 9435
rect 27203 9432 27215 9435
rect 28730 9435 28788 9441
rect 28730 9432 28742 9435
rect 27203 9404 28742 9432
rect 27203 9401 27215 9404
rect 27157 9395 27215 9401
rect 28730 9401 28742 9404
rect 28776 9401 28788 9435
rect 28828 9432 28856 9472
rect 28994 9460 29000 9472
rect 29052 9460 29058 9512
rect 31113 9503 31171 9509
rect 31113 9469 31125 9503
rect 31159 9469 31171 9503
rect 31113 9463 31171 9469
rect 31128 9432 31156 9463
rect 28828 9404 31156 9432
rect 28730 9395 28788 9401
rect 27522 9364 27528 9376
rect 26988 9336 27528 9364
rect 27522 9324 27528 9336
rect 27580 9364 27586 9376
rect 27617 9367 27675 9373
rect 27617 9364 27629 9367
rect 27580 9336 27629 9364
rect 27580 9324 27586 9336
rect 27617 9333 27629 9336
rect 27663 9333 27675 9367
rect 27617 9327 27675 9333
rect 28810 9324 28816 9376
rect 28868 9364 28874 9376
rect 29549 9367 29607 9373
rect 29549 9364 29561 9367
rect 28868 9336 29561 9364
rect 28868 9324 28874 9336
rect 29549 9333 29561 9336
rect 29595 9333 29607 9367
rect 29549 9327 29607 9333
rect 31297 9367 31355 9373
rect 31297 9333 31309 9367
rect 31343 9364 31355 9367
rect 31343 9336 32076 9364
rect 31343 9333 31355 9336
rect 31297 9327 31355 9333
rect 1104 9274 32016 9296
rect 0 9228 800 9242
rect 0 9200 1072 9228
rect 1104 9222 11253 9274
rect 11305 9222 11317 9274
rect 11369 9222 11381 9274
rect 11433 9222 11445 9274
rect 11497 9222 11509 9274
rect 11561 9222 21557 9274
rect 21609 9222 21621 9274
rect 21673 9222 21685 9274
rect 21737 9222 21749 9274
rect 21801 9222 21813 9274
rect 21865 9222 32016 9274
rect 1104 9200 32016 9222
rect 32048 9228 32076 9336
rect 32320 9228 33120 9242
rect 32048 9200 33120 9228
rect 0 9186 800 9200
rect 1044 9092 1072 9200
rect 32320 9186 33120 9200
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1728 9132 1961 9160
rect 1728 9120 1734 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 1949 9123 2007 9129
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 2501 9163 2559 9169
rect 2501 9160 2513 9163
rect 2464 9132 2513 9160
rect 2464 9120 2470 9132
rect 2501 9129 2513 9132
rect 2547 9129 2559 9163
rect 2501 9123 2559 9129
rect 3789 9163 3847 9169
rect 3789 9129 3801 9163
rect 3835 9160 3847 9163
rect 4798 9160 4804 9172
rect 3835 9132 4804 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 5408 9132 5549 9160
rect 5408 9120 5414 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 5537 9123 5595 9129
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 16298 9160 16304 9172
rect 11756 9132 16304 9160
rect 11756 9120 11762 9132
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17586 9160 17592 9172
rect 17368 9132 17592 9160
rect 17368 9120 17374 9132
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22646 9160 22652 9172
rect 22152 9132 22652 9160
rect 22152 9120 22158 9132
rect 22646 9120 22652 9132
rect 22704 9120 22710 9172
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 24213 9163 24271 9169
rect 24213 9160 24225 9163
rect 23532 9132 24225 9160
rect 23532 9120 23538 9132
rect 24213 9129 24225 9132
rect 24259 9129 24271 9163
rect 27614 9160 27620 9172
rect 24213 9123 24271 9129
rect 24872 9132 27620 9160
rect 7190 9092 7196 9104
rect 1044 9064 1900 9092
rect 1872 9033 1900 9064
rect 4448 9064 5672 9092
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2038 9024 2044 9036
rect 1903 8996 2044 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 2774 9024 2780 9036
rect 2280 8996 2780 9024
rect 2280 8984 2286 8996
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 4448 9033 4476 9064
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4433 8987 4491 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4801 9027 4859 9033
rect 4801 8993 4813 9027
rect 4847 9024 4859 9027
rect 4890 9024 4896 9036
rect 4847 8996 4896 9024
rect 4847 8993 4859 8996
rect 4801 8987 4859 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 8993 5043 9027
rect 4985 8987 5043 8993
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8925 4767 8959
rect 5000 8956 5028 8987
rect 5074 8984 5080 9036
rect 5132 9022 5138 9036
rect 5644 9033 5672 9064
rect 6564 9064 7196 9092
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 5184 9022 5457 9024
rect 5132 8996 5457 9022
rect 5132 8994 5212 8996
rect 5132 8984 5138 8994
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 5810 9024 5816 9036
rect 5675 8996 5816 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 6362 9024 6368 9036
rect 6323 8996 6368 9024
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6564 9033 6592 9064
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 9122 9052 9128 9104
rect 9180 9092 9186 9104
rect 10873 9095 10931 9101
rect 9180 9064 9674 9092
rect 9180 9052 9186 9064
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 8993 6607 9027
rect 6549 8987 6607 8993
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6880 8996 6929 9024
rect 6880 8984 6886 8996
rect 6917 8993 6929 8996
rect 6963 8993 6975 9027
rect 7650 9024 7656 9036
rect 7611 8996 7656 9024
rect 6917 8987 6975 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 7920 9027 7978 9033
rect 7920 8993 7932 9027
rect 7966 9024 7978 9027
rect 8938 9024 8944 9036
rect 7966 8996 8944 9024
rect 7966 8993 7978 8996
rect 7920 8987 7978 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 5534 8956 5540 8968
rect 5000 8928 5540 8956
rect 4709 8919 4767 8925
rect 4522 8888 4528 8900
rect 3160 8860 4528 8888
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 3160 8829 3188 8860
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 4724 8888 4752 8919
rect 5534 8916 5540 8928
rect 5592 8956 5598 8968
rect 6380 8956 6408 8984
rect 5592 8928 6408 8956
rect 5592 8916 5598 8928
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6512 8928 6653 8956
rect 6512 8916 6518 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 6472 8888 6500 8916
rect 6748 8888 6776 8919
rect 4724 8860 6500 8888
rect 6656 8860 6776 8888
rect 9033 8891 9091 8897
rect 3145 8823 3203 8829
rect 3145 8820 3157 8823
rect 2280 8792 3157 8820
rect 2280 8780 2286 8792
rect 3145 8789 3157 8792
rect 3191 8789 3203 8823
rect 4246 8820 4252 8832
rect 4207 8792 4252 8820
rect 3145 8783 3203 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 6656 8820 6684 8860
rect 9033 8857 9045 8891
rect 9079 8888 9091 8891
rect 9122 8888 9128 8900
rect 9079 8860 9128 8888
rect 9079 8857 9091 8860
rect 9033 8851 9091 8857
rect 9122 8848 9128 8860
rect 9180 8888 9186 8900
rect 9508 8888 9536 8987
rect 9646 8956 9674 9064
rect 10873 9061 10885 9095
rect 10919 9092 10931 9095
rect 11790 9092 11796 9104
rect 10919 9064 11796 9092
rect 10919 9061 10931 9064
rect 10873 9055 10931 9061
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 11885 9095 11943 9101
rect 11885 9061 11897 9095
rect 11931 9092 11943 9095
rect 13446 9092 13452 9104
rect 11931 9064 13452 9092
rect 11931 9061 11943 9064
rect 11885 9055 11943 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 16206 9092 16212 9104
rect 14200 9064 16212 9092
rect 14200 9036 14228 9064
rect 16206 9052 16212 9064
rect 16264 9092 16270 9104
rect 18877 9095 18935 9101
rect 18877 9092 18889 9095
rect 16264 9064 18889 9092
rect 16264 9052 16270 9064
rect 18877 9061 18889 9064
rect 18923 9092 18935 9095
rect 21174 9092 21180 9104
rect 18923 9064 21180 9092
rect 18923 9061 18935 9064
rect 18877 9055 18935 9061
rect 21174 9052 21180 9064
rect 21232 9052 21238 9104
rect 23842 9092 23848 9104
rect 22296 9064 23704 9092
rect 23803 9064 23848 9092
rect 10134 9024 10140 9036
rect 10095 8996 10140 9024
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 9024 11023 9027
rect 11606 9024 11612 9036
rect 11011 8996 11612 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 11606 8984 11612 8996
rect 11664 9024 11670 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11664 8996 11713 9024
rect 11664 8984 11670 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 12342 9024 12348 9036
rect 12303 8996 12348 9024
rect 11701 8987 11759 8993
rect 11238 8956 11244 8968
rect 9646 8928 11244 8956
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 9180 8860 9536 8888
rect 9585 8891 9643 8897
rect 9180 8848 9186 8860
rect 9585 8857 9597 8891
rect 9631 8888 9643 8891
rect 11606 8888 11612 8900
rect 9631 8860 11612 8888
rect 9631 8857 9643 8860
rect 9585 8851 9643 8857
rect 11606 8848 11612 8860
rect 11664 8848 11670 8900
rect 11716 8888 11744 8987
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12618 9024 12624 9036
rect 12579 8996 12624 9024
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 12805 9027 12863 9033
rect 12805 8993 12817 9027
rect 12851 9024 12863 9027
rect 13630 9024 13636 9036
rect 12851 8996 13636 9024
rect 12851 8993 12863 8996
rect 12805 8987 12863 8993
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12492 8928 12541 8956
rect 12492 8916 12498 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12728 8956 12756 8987
rect 13630 8984 13636 8996
rect 13688 9024 13694 9036
rect 13725 9027 13783 9033
rect 13725 9024 13737 9027
rect 13688 8996 13737 9024
rect 13688 8984 13694 8996
rect 13725 8993 13737 8996
rect 13771 9024 13783 9027
rect 13998 9024 14004 9036
rect 13771 8996 14004 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 13998 8984 14004 8996
rect 14056 8984 14062 9036
rect 14182 9024 14188 9036
rect 14143 8996 14188 9024
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 9024 16727 9027
rect 17218 9024 17224 9036
rect 16715 8996 17224 9024
rect 16715 8993 16727 8996
rect 16669 8987 16727 8993
rect 13078 8956 13084 8968
rect 12728 8928 13084 8956
rect 12529 8919 12587 8925
rect 13078 8916 13084 8928
rect 13136 8956 13142 8968
rect 16684 8956 16712 8987
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 17678 9024 17684 9036
rect 17639 8996 17684 9024
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 18138 9024 18144 9036
rect 17788 8996 18144 9024
rect 17788 8965 17816 8996
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 20530 8984 20536 9036
rect 20588 9024 20594 9036
rect 21985 9027 22043 9033
rect 21985 9024 21997 9027
rect 20588 8996 21997 9024
rect 20588 8984 20594 8996
rect 21985 8993 21997 8996
rect 22031 8993 22043 9027
rect 22296 9026 22324 9064
rect 22204 9022 22324 9026
rect 21985 8987 22043 8993
rect 22112 8998 22324 9022
rect 22112 8994 22232 8998
rect 17773 8959 17831 8965
rect 17773 8956 17785 8959
rect 13136 8928 16712 8956
rect 17236 8928 17785 8956
rect 13136 8916 13142 8928
rect 14274 8888 14280 8900
rect 11716 8860 14280 8888
rect 14274 8848 14280 8860
rect 14332 8848 14338 8900
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 16206 8888 16212 8900
rect 15528 8860 16212 8888
rect 15528 8848 15534 8860
rect 16206 8848 16212 8860
rect 16264 8888 16270 8900
rect 17236 8888 17264 8928
rect 17773 8925 17785 8928
rect 17819 8925 17831 8959
rect 17773 8919 17831 8925
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 20254 8956 20260 8968
rect 17920 8928 20260 8956
rect 17920 8916 17926 8928
rect 20254 8916 20260 8928
rect 20312 8956 20318 8968
rect 22112 8956 22140 8994
rect 22554 8984 22560 9036
rect 22612 9024 22618 9036
rect 22649 9027 22707 9033
rect 22649 9024 22661 9027
rect 22612 8996 22661 9024
rect 22612 8984 22618 8996
rect 22649 8993 22661 8996
rect 22695 8993 22707 9027
rect 22649 8987 22707 8993
rect 22830 8984 22836 9036
rect 22888 9024 22894 9036
rect 23201 9027 23259 9033
rect 22888 8996 23152 9024
rect 22888 8984 22894 8996
rect 20312 8928 22140 8956
rect 22189 8959 22247 8965
rect 20312 8916 20318 8928
rect 22189 8925 22201 8959
rect 22235 8925 22247 8959
rect 22189 8919 22247 8925
rect 16264 8860 17264 8888
rect 16264 8848 16270 8860
rect 17310 8848 17316 8900
rect 17368 8888 17374 8900
rect 18322 8888 18328 8900
rect 17368 8860 18328 8888
rect 17368 8848 17374 8860
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 18506 8848 18512 8900
rect 18564 8888 18570 8900
rect 20070 8888 20076 8900
rect 18564 8860 20076 8888
rect 18564 8848 18570 8860
rect 20070 8848 20076 8860
rect 20128 8888 20134 8900
rect 20128 8860 21229 8888
rect 20128 8848 20134 8860
rect 7098 8820 7104 8832
rect 4764 8792 6684 8820
rect 7059 8792 7104 8820
rect 4764 8780 4770 8792
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 10226 8820 10232 8832
rect 10187 8792 10232 8820
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 10744 8792 11529 8820
rect 10744 8780 10750 8792
rect 11517 8789 11529 8792
rect 11563 8789 11575 8823
rect 11517 8783 11575 8789
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12308 8792 13001 8820
rect 12308 8780 12314 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 13630 8820 13636 8832
rect 13591 8792 13636 8820
rect 12989 8783 13047 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 15657 8823 15715 8829
rect 15657 8789 15669 8823
rect 15703 8820 15715 8823
rect 15746 8820 15752 8832
rect 15703 8792 15752 8820
rect 15703 8789 15715 8792
rect 15657 8783 15715 8789
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16761 8823 16819 8829
rect 16761 8789 16773 8823
rect 16807 8820 16819 8823
rect 16850 8820 16856 8832
rect 16807 8792 16856 8820
rect 16807 8789 16819 8792
rect 16761 8783 16819 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17862 8820 17868 8832
rect 17823 8792 17868 8820
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 18049 8823 18107 8829
rect 18049 8820 18061 8823
rect 18012 8792 18061 8820
rect 18012 8780 18018 8792
rect 18049 8789 18061 8792
rect 18095 8789 18107 8823
rect 18049 8783 18107 8789
rect 19150 8780 19156 8832
rect 19208 8820 19214 8832
rect 20165 8823 20223 8829
rect 20165 8820 20177 8823
rect 19208 8792 20177 8820
rect 19208 8780 19214 8792
rect 20165 8789 20177 8792
rect 20211 8820 20223 8823
rect 20438 8820 20444 8832
rect 20211 8792 20444 8820
rect 20211 8789 20223 8792
rect 20165 8783 20223 8789
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 21201 8820 21229 8860
rect 21266 8848 21272 8900
rect 21324 8888 21330 8900
rect 22204 8888 22232 8919
rect 22278 8916 22284 8968
rect 22336 8956 22342 8968
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 22336 8928 22937 8956
rect 22336 8916 22342 8928
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8925 23075 8959
rect 23124 8956 23152 8996
rect 23201 8993 23213 9027
rect 23247 9024 23259 9027
rect 23566 9024 23572 9036
rect 23247 8996 23572 9024
rect 23247 8993 23259 8996
rect 23201 8987 23259 8993
rect 23566 8984 23572 8996
rect 23624 8984 23630 9036
rect 23676 9024 23704 9064
rect 23842 9052 23848 9064
rect 23900 9052 23906 9104
rect 24061 9095 24119 9101
rect 24061 9061 24073 9095
rect 24107 9092 24119 9095
rect 24762 9092 24768 9104
rect 24107 9064 24768 9092
rect 24107 9061 24119 9064
rect 24061 9055 24119 9061
rect 24762 9052 24768 9064
rect 24820 9052 24826 9104
rect 24872 9024 24900 9132
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 28534 9120 28540 9172
rect 28592 9160 28598 9172
rect 28592 9132 28764 9160
rect 28592 9120 28598 9132
rect 25682 9052 25688 9104
rect 25740 9092 25746 9104
rect 28629 9095 28687 9101
rect 28629 9092 28641 9095
rect 25740 9064 26188 9092
rect 25740 9052 25746 9064
rect 26160 9036 26188 9064
rect 26252 9064 28641 9092
rect 25866 9024 25872 9036
rect 23676 8996 24900 9024
rect 25827 8996 25872 9024
rect 25866 8984 25872 8996
rect 25924 8984 25930 9036
rect 26142 9024 26148 9036
rect 26055 8996 26148 9024
rect 26142 8984 26148 8996
rect 26200 8984 26206 9036
rect 26252 9033 26280 9064
rect 28629 9061 28641 9064
rect 28675 9061 28687 9095
rect 28736 9092 28764 9132
rect 29086 9120 29092 9172
rect 29144 9160 29150 9172
rect 29181 9163 29239 9169
rect 29181 9160 29193 9163
rect 29144 9132 29193 9160
rect 29144 9120 29150 9132
rect 29181 9129 29193 9132
rect 29227 9129 29239 9163
rect 29181 9123 29239 9129
rect 30285 9095 30343 9101
rect 30285 9092 30297 9095
rect 28736 9064 30297 9092
rect 28629 9055 28687 9061
rect 30285 9061 30297 9064
rect 30331 9061 30343 9095
rect 30285 9055 30343 9061
rect 26237 9027 26295 9033
rect 26237 8993 26249 9027
rect 26283 8993 26295 9027
rect 26418 9024 26424 9036
rect 26379 8996 26424 9024
rect 26237 8987 26295 8993
rect 26418 8984 26424 8996
rect 26476 8984 26482 9036
rect 26510 8984 26516 9036
rect 26568 9024 26574 9036
rect 27341 9027 27399 9033
rect 27341 9024 27353 9027
rect 26568 8996 27353 9024
rect 26568 8984 26574 8996
rect 27341 8993 27353 8996
rect 27387 8993 27399 9027
rect 27522 9024 27528 9036
rect 27483 8996 27528 9024
rect 27341 8987 27399 8993
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 27890 9024 27896 9036
rect 27851 8996 27896 9024
rect 27890 8984 27896 8996
rect 27948 9024 27954 9036
rect 28537 9027 28595 9033
rect 28537 9024 28549 9027
rect 27948 8996 28549 9024
rect 27948 8984 27954 8996
rect 28537 8993 28549 8996
rect 28583 8993 28595 9027
rect 28537 8987 28595 8993
rect 29362 8984 29368 9036
rect 29420 9024 29426 9036
rect 30374 9024 30380 9036
rect 29420 8996 30380 9024
rect 29420 8984 29426 8996
rect 30374 8984 30380 8996
rect 30432 8984 30438 9036
rect 23382 8956 23388 8968
rect 23124 8928 23388 8956
rect 23017 8919 23075 8925
rect 21324 8860 22324 8888
rect 21324 8848 21330 8860
rect 21634 8820 21640 8832
rect 21201 8792 21640 8820
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 21818 8820 21824 8832
rect 21779 8792 21824 8820
rect 21818 8780 21824 8792
rect 21876 8780 21882 8832
rect 22296 8820 22324 8860
rect 22462 8848 22468 8900
rect 22520 8888 22526 8900
rect 23032 8888 23060 8919
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 25038 8916 25044 8968
rect 25096 8956 25102 8968
rect 26050 8956 26056 8968
rect 25096 8928 26056 8956
rect 25096 8916 25102 8928
rect 26050 8916 26056 8928
rect 26108 8916 26114 8968
rect 27430 8916 27436 8968
rect 27488 8956 27494 8968
rect 27617 8959 27675 8965
rect 27617 8956 27629 8959
rect 27488 8928 27629 8956
rect 27488 8916 27494 8928
rect 27617 8925 27629 8928
rect 27663 8925 27675 8959
rect 27617 8919 27675 8925
rect 27709 8959 27767 8965
rect 27709 8925 27721 8959
rect 27755 8925 27767 8959
rect 27709 8919 27767 8925
rect 22520 8860 23060 8888
rect 22520 8848 22526 8860
rect 23566 8848 23572 8900
rect 23624 8888 23630 8900
rect 23624 8860 25820 8888
rect 23624 8848 23630 8860
rect 22370 8820 22376 8832
rect 22283 8792 22376 8820
rect 22370 8780 22376 8792
rect 22428 8820 22434 8832
rect 23198 8820 23204 8832
rect 22428 8792 23204 8820
rect 22428 8780 22434 8792
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 23385 8823 23443 8829
rect 23385 8789 23397 8823
rect 23431 8820 23443 8823
rect 23474 8820 23480 8832
rect 23431 8792 23480 8820
rect 23431 8789 23443 8792
rect 23385 8783 23443 8789
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 23934 8780 23940 8832
rect 23992 8820 23998 8832
rect 24029 8823 24087 8829
rect 24029 8820 24041 8823
rect 23992 8792 24041 8820
rect 23992 8780 23998 8792
rect 24029 8789 24041 8792
rect 24075 8820 24087 8823
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 24075 8792 24685 8820
rect 24075 8789 24087 8792
rect 24029 8783 24087 8789
rect 24673 8789 24685 8792
rect 24719 8820 24731 8823
rect 25130 8820 25136 8832
rect 24719 8792 25136 8820
rect 24719 8789 24731 8792
rect 24673 8783 24731 8789
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 25682 8820 25688 8832
rect 25643 8792 25688 8820
rect 25682 8780 25688 8792
rect 25740 8780 25746 8832
rect 25792 8820 25820 8860
rect 26418 8848 26424 8900
rect 26476 8888 26482 8900
rect 26694 8888 26700 8900
rect 26476 8860 26700 8888
rect 26476 8848 26482 8860
rect 26694 8848 26700 8860
rect 26752 8848 26758 8900
rect 27062 8848 27068 8900
rect 27120 8888 27126 8900
rect 27724 8888 27752 8919
rect 27120 8860 27752 8888
rect 28077 8891 28135 8897
rect 27120 8848 27126 8860
rect 28077 8857 28089 8891
rect 28123 8888 28135 8891
rect 29362 8888 29368 8900
rect 28123 8860 29368 8888
rect 28123 8857 28135 8860
rect 28077 8851 28135 8857
rect 29362 8848 29368 8860
rect 29420 8848 29426 8900
rect 29086 8820 29092 8832
rect 25792 8792 29092 8820
rect 29086 8780 29092 8792
rect 29144 8820 29150 8832
rect 29733 8823 29791 8829
rect 29733 8820 29745 8823
rect 29144 8792 29745 8820
rect 29144 8780 29150 8792
rect 29733 8789 29745 8792
rect 29779 8789 29791 8823
rect 30834 8820 30840 8832
rect 30795 8792 30840 8820
rect 29733 8783 29791 8789
rect 30834 8780 30840 8792
rect 30892 8780 30898 8832
rect 1104 8730 32016 8752
rect 1104 8678 6102 8730
rect 6154 8678 6166 8730
rect 6218 8678 6230 8730
rect 6282 8678 6294 8730
rect 6346 8678 6358 8730
rect 6410 8678 16405 8730
rect 16457 8678 16469 8730
rect 16521 8678 16533 8730
rect 16585 8678 16597 8730
rect 16649 8678 16661 8730
rect 16713 8678 26709 8730
rect 26761 8678 26773 8730
rect 26825 8678 26837 8730
rect 26889 8678 26901 8730
rect 26953 8678 26965 8730
rect 27017 8678 32016 8730
rect 1104 8656 32016 8678
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5810 8616 5816 8628
rect 5399 8588 5816 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 8386 8616 8392 8628
rect 8347 8588 8392 8616
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10192 8588 10609 8616
rect 10192 8576 10198 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 11793 8619 11851 8625
rect 10597 8579 10655 8585
rect 10888 8588 11652 8616
rect 2130 8508 2136 8560
rect 2188 8548 2194 8560
rect 2317 8551 2375 8557
rect 2317 8548 2329 8551
rect 2188 8520 2329 8548
rect 2188 8508 2194 8520
rect 2317 8517 2329 8520
rect 2363 8548 2375 8551
rect 2363 8520 4016 8548
rect 2363 8517 2375 8520
rect 2317 8511 2375 8517
rect 2498 8440 2504 8492
rect 2556 8480 2562 8492
rect 2556 8452 2601 8480
rect 2556 8440 2562 8452
rect 2682 8440 2688 8492
rect 2740 8480 2746 8492
rect 3988 8480 4016 8520
rect 5074 8508 5080 8560
rect 5132 8548 5138 8560
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 5132 8520 6469 8548
rect 5132 8508 5138 8520
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 6822 8548 6828 8560
rect 6503 8520 6828 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 10888 8548 10916 8588
rect 10284 8520 10916 8548
rect 10284 8508 10290 8520
rect 2740 8452 3188 8480
rect 3988 8452 4108 8480
rect 2740 8440 2746 8452
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8381 1823 8415
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 1765 8375 1823 8381
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 1673 8347 1731 8353
rect 1673 8344 1685 8347
rect 1636 8316 1685 8344
rect 1636 8304 1642 8316
rect 1673 8313 1685 8316
rect 1719 8313 1731 8347
rect 1780 8344 1808 8375
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2700 8412 2728 8440
rect 2332 8384 2728 8412
rect 2332 8344 2360 8384
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 3160 8421 3188 8452
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2832 8384 2973 8412
rect 2832 8372 2838 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 3786 8372 3792 8424
rect 3844 8412 3850 8424
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3844 8384 3985 8412
rect 3844 8372 3850 8384
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 1780 8316 2360 8344
rect 2501 8347 2559 8353
rect 1673 8307 1731 8313
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 3234 8344 3240 8356
rect 2547 8316 3240 8344
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 4080 8344 4108 8452
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11333 8483 11391 8489
rect 11333 8480 11345 8483
rect 11020 8452 11345 8480
rect 11020 8440 11026 8452
rect 11333 8449 11345 8452
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 4246 8421 4252 8424
rect 4240 8412 4252 8421
rect 4207 8384 4252 8412
rect 4240 8375 4252 8384
rect 4246 8372 4252 8375
rect 4304 8372 4310 8424
rect 5902 8412 5908 8424
rect 4356 8384 5908 8412
rect 4356 8344 4384 8384
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7570 8415 7628 8421
rect 7570 8412 7582 8415
rect 7156 8384 7582 8412
rect 7156 8372 7162 8384
rect 7570 8381 7582 8384
rect 7616 8381 7628 8415
rect 7570 8375 7628 8381
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 7800 8384 7849 8412
rect 7800 8372 7806 8384
rect 7837 8381 7849 8384
rect 7883 8381 7895 8415
rect 7837 8375 7895 8381
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8412 9275 8415
rect 10870 8412 10876 8424
rect 9263 8384 10876 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11054 8412 11060 8424
rect 11015 8384 11060 8412
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 11624 8421 11652 8588
rect 11793 8585 11805 8619
rect 11839 8616 11851 8619
rect 12618 8616 12624 8628
rect 11839 8588 12624 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12894 8616 12900 8628
rect 12855 8588 12900 8616
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 14090 8616 14096 8628
rect 14051 8588 14096 8616
rect 14090 8576 14096 8588
rect 14148 8616 14154 8628
rect 14826 8616 14832 8628
rect 14148 8588 14832 8616
rect 14148 8576 14154 8588
rect 14826 8576 14832 8588
rect 14884 8616 14890 8628
rect 15562 8616 15568 8628
rect 14884 8588 15568 8616
rect 14884 8576 14890 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 19518 8616 19524 8628
rect 18840 8588 19524 8616
rect 18840 8576 18846 8588
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 20990 8576 20996 8628
rect 21048 8616 21054 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 21048 8588 21373 8616
rect 21048 8576 21054 8588
rect 13078 8548 13084 8560
rect 12636 8520 13084 8548
rect 12066 8440 12072 8492
rect 12124 8480 12130 8492
rect 12636 8489 12664 8520
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 16942 8508 16948 8560
rect 17000 8548 17006 8560
rect 17126 8548 17132 8560
rect 17000 8520 17132 8548
rect 17000 8508 17006 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17770 8508 17776 8560
rect 17828 8508 17834 8560
rect 18141 8551 18199 8557
rect 18141 8517 18153 8551
rect 18187 8548 18199 8551
rect 18230 8548 18236 8560
rect 18187 8520 18236 8548
rect 18187 8517 18199 8520
rect 18141 8511 18199 8517
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 18417 8551 18475 8557
rect 18417 8517 18429 8551
rect 18463 8548 18475 8551
rect 19334 8548 19340 8560
rect 18463 8520 19340 8548
rect 18463 8517 18475 8520
rect 18417 8511 18475 8517
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12124 8452 12541 8480
rect 12124 8440 12130 8452
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8449 12679 8483
rect 13630 8480 13636 8492
rect 12621 8443 12679 8449
rect 12728 8452 13636 8480
rect 11241 8415 11299 8421
rect 11241 8412 11253 8415
rect 11204 8384 11253 8412
rect 11204 8372 11210 8384
rect 11241 8381 11253 8384
rect 11287 8381 11299 8415
rect 11241 8375 11299 8381
rect 11425 8415 11483 8421
rect 11425 8381 11437 8415
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8381 11667 8415
rect 12250 8412 12256 8424
rect 12211 8384 12256 8412
rect 11609 8375 11667 8381
rect 4080 8316 4384 8344
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 9484 8347 9542 8353
rect 5408 8316 6132 8344
rect 5408 8304 5414 8316
rect 1394 8236 1400 8288
rect 1452 8276 1458 8288
rect 2222 8276 2228 8288
rect 1452 8248 2228 8276
rect 1452 8236 1458 8248
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 3050 8276 3056 8288
rect 3011 8248 3056 8276
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 5905 8279 5963 8285
rect 5905 8245 5917 8279
rect 5951 8276 5963 8279
rect 5994 8276 6000 8288
rect 5951 8248 6000 8276
rect 5951 8245 5963 8248
rect 5905 8239 5963 8245
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 6104 8276 6132 8316
rect 9484 8313 9496 8347
rect 9530 8344 9542 8347
rect 9582 8344 9588 8356
rect 9530 8316 9588 8344
rect 9530 8313 9542 8316
rect 9484 8307 9542 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11440 8344 11468 8375
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12728 8421 12756 8452
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 17788 8480 17816 8508
rect 15405 8452 17816 8480
rect 18049 8483 18107 8489
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 10744 8316 11468 8344
rect 12452 8344 12480 8375
rect 13170 8372 13176 8424
rect 13228 8412 13234 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 13228 8384 13369 8412
rect 13228 8372 13234 8384
rect 13357 8381 13369 8384
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 15405 8412 15433 8452
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18322 8480 18328 8492
rect 18095 8452 18328 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19208 8452 19993 8480
rect 19208 8440 19214 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 21201 8480 21229 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 23566 8616 23572 8628
rect 21692 8588 23572 8616
rect 21692 8576 21698 8588
rect 23566 8576 23572 8588
rect 23624 8576 23630 8628
rect 24762 8616 24768 8628
rect 24723 8588 24768 8616
rect 24762 8576 24768 8588
rect 24820 8576 24826 8628
rect 27338 8616 27344 8628
rect 27299 8588 27344 8616
rect 27338 8576 27344 8588
rect 27396 8576 27402 8628
rect 28074 8576 28080 8628
rect 28132 8616 28138 8628
rect 28445 8619 28503 8625
rect 28445 8616 28457 8619
rect 28132 8588 28457 8616
rect 28132 8576 28138 8588
rect 28445 8585 28457 8588
rect 28491 8585 28503 8619
rect 28445 8579 28503 8585
rect 29454 8576 29460 8628
rect 29512 8616 29518 8628
rect 29549 8619 29607 8625
rect 29549 8616 29561 8619
rect 29512 8588 29561 8616
rect 29512 8576 29518 8588
rect 29549 8585 29561 8588
rect 29595 8585 29607 8619
rect 29549 8579 29607 8585
rect 21450 8508 21456 8560
rect 21508 8548 21514 8560
rect 21910 8548 21916 8560
rect 21508 8520 21916 8548
rect 21508 8508 21514 8520
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 23753 8551 23811 8557
rect 23753 8548 23765 8551
rect 23440 8520 23765 8548
rect 23440 8508 23446 8520
rect 23753 8517 23765 8520
rect 23799 8548 23811 8551
rect 24946 8548 24952 8560
rect 23799 8520 24952 8548
rect 23799 8517 23811 8520
rect 23753 8511 23811 8517
rect 24946 8508 24952 8520
rect 25004 8508 25010 8560
rect 25866 8508 25872 8560
rect 25924 8548 25930 8560
rect 27893 8551 27951 8557
rect 27893 8548 27905 8551
rect 25924 8520 27905 8548
rect 25924 8508 25930 8520
rect 27893 8517 27905 8520
rect 27939 8517 27951 8551
rect 27893 8511 27951 8517
rect 28166 8508 28172 8560
rect 28224 8548 28230 8560
rect 30653 8551 30711 8557
rect 30653 8548 30665 8551
rect 28224 8520 30665 8548
rect 28224 8508 28230 8520
rect 30653 8517 30665 8520
rect 30699 8517 30711 8551
rect 30653 8511 30711 8517
rect 25409 8483 25467 8489
rect 21201 8452 21972 8480
rect 19981 8443 20039 8449
rect 13596 8384 15433 8412
rect 15473 8415 15531 8421
rect 13596 8372 13602 8384
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15746 8412 15752 8424
rect 15519 8384 15752 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 16264 8384 16313 8412
rect 16264 8372 16270 8384
rect 16301 8381 16313 8384
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 16393 8415 16451 8421
rect 16393 8381 16405 8415
rect 16439 8412 16451 8415
rect 17770 8412 17776 8424
rect 16439 8384 17632 8412
rect 17731 8384 17776 8412
rect 16439 8381 16451 8384
rect 16393 8375 16451 8381
rect 14366 8344 14372 8356
rect 12452 8316 14372 8344
rect 10744 8304 10750 8316
rect 14366 8304 14372 8316
rect 14424 8304 14430 8356
rect 14918 8304 14924 8356
rect 14976 8344 14982 8356
rect 15206 8347 15264 8353
rect 15206 8344 15218 8347
rect 14976 8316 15218 8344
rect 14976 8304 14982 8316
rect 15206 8313 15218 8316
rect 15252 8313 15264 8347
rect 15206 8307 15264 8313
rect 17034 8304 17040 8356
rect 17092 8344 17098 8356
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 17092 8316 17141 8344
rect 17092 8304 17098 8316
rect 17129 8313 17141 8316
rect 17175 8313 17187 8347
rect 17310 8344 17316 8356
rect 17271 8316 17316 8344
rect 17129 8307 17187 8313
rect 17310 8304 17316 8316
rect 17368 8304 17374 8356
rect 17604 8344 17632 8384
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 17954 8412 17960 8424
rect 17915 8384 17960 8412
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18233 8415 18291 8421
rect 18233 8381 18245 8415
rect 18279 8381 18291 8415
rect 18233 8375 18291 8381
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8412 19395 8415
rect 21818 8412 21824 8424
rect 19383 8384 21824 8412
rect 19383 8381 19395 8384
rect 19337 8375 19395 8381
rect 18046 8344 18052 8356
rect 17604 8316 18052 8344
rect 18046 8304 18052 8316
rect 18104 8344 18110 8356
rect 18248 8344 18276 8375
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 21944 8412 21972 8452
rect 25409 8449 25421 8483
rect 25455 8480 25467 8483
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 25455 8452 26065 8480
rect 25455 8449 25467 8452
rect 25409 8443 25467 8449
rect 26053 8449 26065 8452
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 26694 8440 26700 8492
rect 26752 8480 26758 8492
rect 26752 8452 27200 8480
rect 26752 8440 26758 8452
rect 22370 8412 22376 8424
rect 21944 8384 22232 8412
rect 22331 8384 22376 8412
rect 20226 8347 20284 8353
rect 20226 8344 20238 8347
rect 18104 8316 18276 8344
rect 19536 8316 20238 8344
rect 18104 8304 18110 8316
rect 11698 8276 11704 8288
rect 6104 8248 11704 8276
rect 11698 8236 11704 8248
rect 11756 8236 11762 8288
rect 16942 8276 16948 8288
rect 16903 8248 16948 8276
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 18138 8276 18144 8288
rect 18012 8248 18144 8276
rect 18012 8236 18018 8248
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 19242 8276 19248 8288
rect 18564 8248 19248 8276
rect 18564 8236 18570 8248
rect 19242 8236 19248 8248
rect 19300 8236 19306 8288
rect 19536 8285 19564 8316
rect 20226 8313 20238 8316
rect 20272 8313 20284 8347
rect 20226 8307 20284 8313
rect 21358 8304 21364 8356
rect 21416 8344 21422 8356
rect 22094 8344 22100 8356
rect 21416 8316 22100 8344
rect 21416 8304 21422 8316
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 22204 8344 22232 8384
rect 22370 8372 22376 8384
rect 22428 8372 22434 8424
rect 23934 8412 23940 8424
rect 22583 8384 23940 8412
rect 22583 8344 22611 8384
rect 23934 8372 23940 8384
rect 23992 8372 23998 8424
rect 25958 8412 25964 8424
rect 25919 8384 25964 8412
rect 25958 8372 25964 8384
rect 26016 8372 26022 8424
rect 26145 8415 26203 8421
rect 26145 8381 26157 8415
rect 26191 8412 26203 8415
rect 26418 8412 26424 8424
rect 26191 8384 26424 8412
rect 26191 8381 26203 8384
rect 26145 8375 26203 8381
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 26510 8372 26516 8424
rect 26568 8412 26574 8424
rect 26605 8415 26663 8421
rect 26605 8412 26617 8415
rect 26568 8384 26617 8412
rect 26568 8372 26574 8384
rect 26605 8381 26617 8384
rect 26651 8381 26663 8415
rect 26605 8375 26663 8381
rect 26789 8415 26847 8421
rect 26789 8381 26801 8415
rect 26835 8381 26847 8415
rect 26789 8375 26847 8381
rect 26881 8415 26939 8421
rect 26881 8381 26893 8415
rect 26927 8381 26939 8415
rect 26881 8375 26939 8381
rect 26973 8415 27031 8421
rect 26973 8381 26985 8415
rect 27019 8412 27031 8415
rect 27062 8412 27068 8424
rect 27019 8384 27068 8412
rect 27019 8381 27031 8384
rect 26973 8375 27031 8381
rect 22646 8353 22652 8356
rect 22204 8316 22611 8344
rect 22640 8307 22652 8353
rect 22704 8344 22710 8356
rect 22704 8316 22740 8344
rect 22646 8304 22652 8307
rect 22704 8304 22710 8316
rect 24762 8304 24768 8356
rect 24820 8344 24826 8356
rect 25133 8347 25191 8353
rect 25133 8344 25145 8347
rect 24820 8316 25145 8344
rect 24820 8304 24826 8316
rect 25133 8313 25145 8316
rect 25179 8313 25191 8347
rect 25133 8307 25191 8313
rect 25225 8347 25283 8353
rect 25225 8313 25237 8347
rect 25271 8344 25283 8347
rect 26326 8344 26332 8356
rect 25271 8316 26332 8344
rect 25271 8313 25283 8316
rect 25225 8307 25283 8313
rect 26326 8304 26332 8316
rect 26384 8344 26390 8356
rect 26804 8344 26832 8375
rect 26384 8316 26832 8344
rect 26896 8344 26924 8375
rect 27062 8372 27068 8384
rect 27120 8372 27126 8424
rect 27172 8421 27200 8452
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 30926 8480 30932 8492
rect 28960 8452 30932 8480
rect 28960 8440 28966 8452
rect 30926 8440 30932 8452
rect 30984 8480 30990 8492
rect 31205 8483 31263 8489
rect 31205 8480 31217 8483
rect 30984 8452 31217 8480
rect 30984 8440 30990 8452
rect 31205 8449 31217 8452
rect 31251 8449 31263 8483
rect 31205 8443 31263 8449
rect 27157 8415 27215 8421
rect 27157 8381 27169 8415
rect 27203 8381 27215 8415
rect 27157 8375 27215 8381
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 27801 8415 27859 8421
rect 27801 8412 27813 8415
rect 27580 8384 27813 8412
rect 27580 8372 27586 8384
rect 27801 8381 27813 8384
rect 27847 8381 27859 8415
rect 27801 8375 27859 8381
rect 27430 8344 27436 8356
rect 26896 8316 27436 8344
rect 26384 8304 26390 8316
rect 27430 8304 27436 8316
rect 27488 8304 27494 8356
rect 30193 8347 30251 8353
rect 30193 8313 30205 8347
rect 30239 8344 30251 8347
rect 30374 8344 30380 8356
rect 30239 8316 30380 8344
rect 30239 8313 30251 8316
rect 30193 8307 30251 8313
rect 19521 8279 19579 8285
rect 19521 8245 19533 8279
rect 19567 8245 19579 8279
rect 19521 8239 19579 8245
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 21082 8276 21088 8288
rect 20772 8248 21088 8276
rect 20772 8236 20778 8248
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 21266 8236 21272 8288
rect 21324 8276 21330 8288
rect 30208 8276 30236 8307
rect 30374 8304 30380 8316
rect 30432 8304 30438 8356
rect 21324 8248 30236 8276
rect 21324 8236 21330 8248
rect 1104 8186 32016 8208
rect 1104 8134 11253 8186
rect 11305 8134 11317 8186
rect 11369 8134 11381 8186
rect 11433 8134 11445 8186
rect 11497 8134 11509 8186
rect 11561 8134 21557 8186
rect 21609 8134 21621 8186
rect 21673 8134 21685 8186
rect 21737 8134 21749 8186
rect 21801 8134 21813 8186
rect 21865 8134 32016 8186
rect 1104 8112 32016 8134
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 8297 8075 8355 8081
rect 2464 8044 2774 8072
rect 2464 8032 2470 8044
rect 1670 7964 1676 8016
rect 1728 8004 1734 8016
rect 2746 8004 2774 8044
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 9582 8072 9588 8084
rect 8343 8044 9444 8072
rect 9543 8044 9588 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 6730 8004 6736 8016
rect 1728 7976 2084 8004
rect 2746 7976 6736 8004
rect 1728 7964 1734 7976
rect 2056 7945 2084 7976
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 9122 8004 9128 8016
rect 9048 7976 9128 8004
rect 2021 7939 2084 7945
rect 2021 7905 2033 7939
rect 2067 7905 2084 7939
rect 2021 7899 2084 7905
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7905 2191 7939
rect 2133 7899 2191 7905
rect 2222 7899 2228 7951
rect 2280 7939 2286 7951
rect 2409 7939 2467 7945
rect 2280 7911 2325 7939
rect 2280 7899 2286 7911
rect 2409 7905 2421 7939
rect 2455 7936 2467 7939
rect 2682 7936 2688 7948
rect 2455 7908 2688 7936
rect 2455 7905 2467 7908
rect 2409 7899 2467 7905
rect 2056 7800 2084 7899
rect 2148 7868 2176 7899
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 3234 7936 3240 7948
rect 3195 7908 3240 7936
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3881 7939 3939 7945
rect 3881 7936 3893 7939
rect 3344 7908 3893 7936
rect 2958 7868 2964 7880
rect 2148 7840 2964 7868
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3142 7828 3148 7880
rect 3200 7868 3206 7880
rect 3344 7868 3372 7908
rect 3881 7905 3893 7908
rect 3927 7905 3939 7939
rect 3881 7899 3939 7905
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 4856 7908 5457 7936
rect 4856 7896 4862 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 5810 7936 5816 7948
rect 5675 7908 5816 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6880 7908 6929 7936
rect 6880 7896 6886 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 8386 7936 8392 7948
rect 8347 7908 8392 7936
rect 7469 7899 7527 7905
rect 3510 7868 3516 7880
rect 3200 7840 3372 7868
rect 3471 7840 3516 7868
rect 3200 7828 3206 7840
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4706 7868 4712 7880
rect 4295 7840 4712 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5534 7868 5540 7880
rect 5040 7840 5540 7868
rect 5040 7828 5046 7840
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 7484 7868 7512 7899
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 8846 7936 8852 7948
rect 8807 7908 8852 7936
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 9048 7945 9076 7976
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 9306 7964 9312 8016
rect 9364 7964 9370 8016
rect 9416 8004 9444 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10336 8044 11008 8072
rect 10336 8004 10364 8044
rect 10980 8004 11008 8044
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 11112 8044 11529 8072
rect 11112 8032 11118 8044
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 11756 8044 22600 8072
rect 11756 8032 11762 8044
rect 9416 7976 10364 8004
rect 10428 7976 10732 8004
rect 10980 7976 12112 8004
rect 9033 7939 9091 7945
rect 9033 7905 9045 7939
rect 9079 7905 9091 7939
rect 9324 7936 9352 7964
rect 9033 7899 9091 7905
rect 9140 7908 9352 7936
rect 9401 7939 9459 7945
rect 9140 7877 9168 7908
rect 9401 7905 9413 7939
rect 9447 7936 9459 7939
rect 10042 7936 10048 7948
rect 9447 7908 10048 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 10428 7945 10456 7976
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7905 10471 7939
rect 10413 7899 10471 7905
rect 10522 7939 10580 7945
rect 10522 7905 10534 7939
rect 10568 7936 10580 7939
rect 10704 7936 10732 7976
rect 10568 7908 10640 7936
rect 10704 7908 11468 7936
rect 10568 7905 10580 7908
rect 10522 7899 10580 7905
rect 5960 7840 7512 7868
rect 9125 7871 9183 7877
rect 5960 7828 5966 7840
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9306 7868 9312 7880
rect 9263 7840 9312 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 2682 7800 2688 7812
rect 2056 7772 2688 7800
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 3697 7803 3755 7809
rect 3697 7769 3709 7803
rect 3743 7800 3755 7803
rect 5350 7800 5356 7812
rect 3743 7772 5356 7800
rect 3743 7769 3755 7772
rect 3697 7763 3755 7769
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 6546 7800 6552 7812
rect 5460 7772 6552 7800
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 1765 7735 1823 7741
rect 1765 7732 1777 7735
rect 1728 7704 1777 7732
rect 1728 7692 1734 7704
rect 1765 7701 1777 7704
rect 1811 7701 1823 7735
rect 1765 7695 1823 7701
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 2774 7732 2780 7744
rect 2004 7704 2780 7732
rect 2004 7692 2010 7704
rect 2774 7692 2780 7704
rect 2832 7692 2838 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 4028 7704 4997 7732
rect 4028 7692 4034 7704
rect 4985 7701 4997 7704
rect 5031 7732 5043 7735
rect 5460 7732 5488 7772
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 6825 7803 6883 7809
rect 6825 7800 6837 7803
rect 6696 7772 6837 7800
rect 6696 7760 6702 7772
rect 6825 7769 6837 7772
rect 6871 7769 6883 7803
rect 6825 7763 6883 7769
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 10152 7800 10180 7899
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10612 7868 10640 7908
rect 10376 7840 10640 7868
rect 11440 7868 11468 7908
rect 11606 7896 11612 7948
rect 11664 7936 11670 7948
rect 12084 7945 12112 7976
rect 12250 7964 12256 8016
rect 12308 8004 12314 8016
rect 12713 8007 12771 8013
rect 12713 8004 12725 8007
rect 12308 7976 12725 8004
rect 12308 7964 12314 7976
rect 12713 7973 12725 7976
rect 12759 7973 12771 8007
rect 12713 7967 12771 7973
rect 12897 8007 12955 8013
rect 12897 7973 12909 8007
rect 12943 8004 12955 8007
rect 13446 8004 13452 8016
rect 12943 7976 13452 8004
rect 12943 7973 12955 7976
rect 12897 7967 12955 7973
rect 13446 7964 13452 7976
rect 13504 7964 13510 8016
rect 13541 8007 13599 8013
rect 13541 7973 13553 8007
rect 13587 8004 13599 8007
rect 13630 8004 13636 8016
rect 13587 7976 13636 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 17586 8004 17592 8016
rect 16546 7976 17592 8004
rect 11701 7939 11759 7945
rect 11701 7936 11713 7939
rect 11664 7908 11713 7936
rect 11664 7896 11670 7908
rect 11701 7905 11713 7908
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 11808 7868 11836 7899
rect 12342 7896 12348 7948
rect 12400 7936 12406 7948
rect 12526 7936 12532 7948
rect 12400 7908 12532 7936
rect 12400 7896 12406 7908
rect 12526 7896 12532 7908
rect 12584 7936 12590 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 12584 7908 13369 7936
rect 12584 7896 12590 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 13722 7936 13728 7948
rect 13683 7908 13728 7936
rect 13357 7899 13415 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 15390 7939 15448 7945
rect 15390 7936 15402 7939
rect 15068 7908 15402 7936
rect 15068 7896 15074 7908
rect 15390 7905 15402 7908
rect 15436 7905 15448 7939
rect 15390 7899 15448 7905
rect 13170 7868 13176 7880
rect 11440 7840 13176 7868
rect 10376 7828 10382 7840
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7868 15715 7871
rect 15746 7868 15752 7880
rect 15703 7840 15752 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 8352 7772 10180 7800
rect 8352 7760 8358 7772
rect 13906 7760 13912 7812
rect 13964 7800 13970 7812
rect 14277 7803 14335 7809
rect 14277 7800 14289 7803
rect 13964 7772 14289 7800
rect 13964 7760 13970 7772
rect 14277 7769 14289 7772
rect 14323 7769 14335 7803
rect 14277 7763 14335 7769
rect 5031 7704 5488 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5629 7735 5687 7741
rect 5629 7732 5641 7735
rect 5592 7704 5641 7732
rect 5592 7692 5598 7704
rect 5629 7701 5641 7704
rect 5675 7732 5687 7735
rect 6914 7732 6920 7744
rect 5675 7704 6920 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 10226 7732 10232 7744
rect 10187 7704 10232 7732
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 10689 7735 10747 7741
rect 10689 7732 10701 7735
rect 10652 7704 10701 7732
rect 10652 7692 10658 7704
rect 10689 7701 10701 7704
rect 10735 7701 10747 7735
rect 10689 7695 10747 7701
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11977 7735 12035 7741
rect 11977 7732 11989 7735
rect 10836 7704 11989 7732
rect 10836 7692 10842 7704
rect 11977 7701 11989 7704
rect 12023 7732 12035 7735
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12023 7704 12541 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12529 7701 12541 7704
rect 12575 7732 12587 7735
rect 12710 7732 12716 7744
rect 12575 7704 12716 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 12710 7692 12716 7704
rect 12768 7732 12774 7744
rect 13814 7732 13820 7744
rect 12768 7704 13820 7732
rect 12768 7692 12774 7704
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 16546 7732 16574 7976
rect 17586 7964 17592 7976
rect 17644 7964 17650 8016
rect 18138 8004 18144 8016
rect 17972 7976 18144 8004
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7936 16727 7939
rect 16758 7936 16764 7948
rect 16715 7908 16764 7936
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 16853 7939 16911 7945
rect 16853 7905 16865 7939
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 16862 7868 16890 7899
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17221 7939 17279 7945
rect 17000 7908 17045 7936
rect 17000 7896 17006 7908
rect 17221 7905 17233 7939
rect 17267 7936 17279 7939
rect 17267 7908 17816 7936
rect 17267 7905 17279 7908
rect 17221 7899 17279 7905
rect 16684 7840 16890 7868
rect 17037 7871 17095 7877
rect 16684 7812 16712 7840
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 16666 7760 16672 7812
rect 16724 7760 16730 7812
rect 17052 7800 17080 7831
rect 17218 7800 17224 7812
rect 17052 7772 17224 7800
rect 17218 7760 17224 7772
rect 17276 7760 17282 7812
rect 17788 7800 17816 7908
rect 17972 7868 18000 7976
rect 18138 7964 18144 7976
rect 18196 7964 18202 8016
rect 18325 8007 18383 8013
rect 18325 7973 18337 8007
rect 18371 7973 18383 8007
rect 18325 7967 18383 7973
rect 19420 8007 19478 8013
rect 19420 7973 19432 8007
rect 19466 8004 19478 8007
rect 19518 8004 19524 8016
rect 19466 7976 19524 8004
rect 19466 7973 19478 7976
rect 19420 7967 19478 7973
rect 18233 7939 18291 7945
rect 18233 7905 18245 7939
rect 18279 7934 18291 7939
rect 18340 7936 18368 7967
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 21085 8007 21143 8013
rect 21085 7973 21097 8007
rect 21131 8004 21143 8007
rect 21266 8004 21272 8016
rect 21131 7976 21272 8004
rect 21131 7973 21143 7976
rect 21085 7967 21143 7973
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 22572 8004 22600 8044
rect 22646 8032 22652 8084
rect 22704 8072 22710 8084
rect 22741 8075 22799 8081
rect 22741 8072 22753 8075
rect 22704 8044 22753 8072
rect 22704 8032 22710 8044
rect 22741 8041 22753 8044
rect 22787 8041 22799 8075
rect 22741 8035 22799 8041
rect 24486 8032 24492 8084
rect 24544 8072 24550 8084
rect 24581 8075 24639 8081
rect 24581 8072 24593 8075
rect 24544 8044 24593 8072
rect 24544 8032 24550 8044
rect 24581 8041 24593 8044
rect 24627 8041 24639 8075
rect 24581 8035 24639 8041
rect 25777 8075 25835 8081
rect 25777 8041 25789 8075
rect 25823 8072 25835 8075
rect 25958 8072 25964 8084
rect 25823 8044 25964 8072
rect 25823 8041 25835 8044
rect 25777 8035 25835 8041
rect 25958 8032 25964 8044
rect 26016 8032 26022 8084
rect 27890 8072 27896 8084
rect 27264 8044 27896 8072
rect 23474 8013 23480 8016
rect 23468 8004 23480 8013
rect 22572 7976 22784 8004
rect 23435 7976 23480 8004
rect 19702 7936 19708 7948
rect 18340 7934 19380 7936
rect 19518 7934 19708 7936
rect 18279 7905 18312 7934
rect 18340 7908 19708 7934
rect 19352 7906 19546 7908
rect 18233 7899 18312 7905
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17972 7840 18061 7868
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18284 7868 18312 7899
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 22005 7939 22063 7945
rect 22005 7905 22017 7939
rect 22051 7905 22063 7939
rect 22005 7899 22063 7905
rect 18874 7868 18880 7880
rect 18284 7840 18880 7868
rect 18049 7831 18107 7837
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19150 7868 19156 7880
rect 19111 7840 19156 7868
rect 19150 7828 19156 7840
rect 19208 7828 19214 7880
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 22020 7868 22048 7899
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22189 7939 22247 7945
rect 22189 7936 22201 7939
rect 22152 7908 22201 7936
rect 22152 7896 22158 7908
rect 22189 7905 22201 7908
rect 22235 7905 22247 7939
rect 22462 7936 22468 7948
rect 22189 7899 22247 7905
rect 22388 7908 22468 7936
rect 22278 7868 22284 7880
rect 20404 7840 22140 7868
rect 22239 7840 22284 7868
rect 20404 7828 20410 7840
rect 18506 7800 18512 7812
rect 17788 7772 18512 7800
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 20530 7800 20536 7812
rect 20491 7772 20536 7800
rect 20530 7760 20536 7772
rect 20588 7760 20594 7812
rect 21266 7760 21272 7812
rect 21324 7800 21330 7812
rect 22002 7800 22008 7812
rect 21324 7772 22008 7800
rect 21324 7760 21330 7772
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 22112 7800 22140 7840
rect 22278 7828 22284 7840
rect 22336 7828 22342 7880
rect 22388 7877 22416 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 22568 7939 22626 7945
rect 22568 7905 22580 7939
rect 22614 7905 22626 7939
rect 22756 7936 22784 7976
rect 23468 7967 23480 7976
rect 23474 7964 23480 7967
rect 23532 7964 23538 8016
rect 25498 7964 25504 8016
rect 25556 8004 25562 8016
rect 25556 7976 26280 8004
rect 25556 7964 25562 7976
rect 22756 7908 24256 7936
rect 22568 7899 22626 7905
rect 22373 7871 22431 7877
rect 22373 7837 22385 7871
rect 22419 7837 22431 7871
rect 22572 7868 22600 7899
rect 22830 7868 22836 7880
rect 22572 7840 22836 7868
rect 22373 7831 22431 7837
rect 22830 7828 22836 7840
rect 22888 7828 22894 7880
rect 23201 7871 23259 7877
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 22646 7800 22652 7812
rect 22112 7772 22652 7800
rect 22646 7760 22652 7772
rect 22704 7760 22710 7812
rect 16172 7704 16574 7732
rect 17405 7735 17463 7741
rect 16172 7692 16178 7704
rect 17405 7701 17417 7735
rect 17451 7732 17463 7735
rect 18414 7732 18420 7744
rect 17451 7704 18420 7732
rect 17451 7701 17463 7704
rect 17405 7695 17463 7701
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 18693 7735 18751 7741
rect 18693 7701 18705 7735
rect 18739 7732 18751 7735
rect 19794 7732 19800 7744
rect 18739 7704 19800 7732
rect 18739 7701 18751 7704
rect 18693 7695 18751 7701
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 22020 7732 22048 7760
rect 22922 7732 22928 7744
rect 22020 7704 22928 7732
rect 22922 7692 22928 7704
rect 22980 7692 22986 7744
rect 23216 7732 23244 7831
rect 24228 7800 24256 7908
rect 24670 7896 24676 7948
rect 24728 7936 24734 7948
rect 25409 7939 25467 7945
rect 25409 7936 25421 7939
rect 24728 7908 25421 7936
rect 24728 7896 24734 7908
rect 25409 7905 25421 7908
rect 25455 7905 25467 7939
rect 25590 7936 25596 7948
rect 25551 7908 25596 7936
rect 25409 7899 25467 7905
rect 25424 7868 25452 7899
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 26252 7945 26280 7976
rect 26237 7939 26295 7945
rect 26237 7905 26249 7939
rect 26283 7905 26295 7939
rect 26237 7899 26295 7905
rect 26510 7896 26516 7948
rect 26568 7936 26574 7948
rect 27264 7945 27292 8044
rect 27890 8032 27896 8044
rect 27948 8072 27954 8084
rect 28261 8075 28319 8081
rect 28261 8072 28273 8075
rect 27948 8044 28273 8072
rect 27948 8032 27954 8044
rect 28261 8041 28273 8044
rect 28307 8041 28319 8075
rect 28261 8035 28319 8041
rect 28350 8032 28356 8084
rect 28408 8072 28414 8084
rect 30653 8075 30711 8081
rect 30653 8072 30665 8075
rect 28408 8044 30665 8072
rect 28408 8032 28414 8044
rect 30653 8041 30665 8044
rect 30699 8041 30711 8075
rect 30653 8035 30711 8041
rect 30742 8032 30748 8084
rect 30800 8072 30806 8084
rect 31205 8075 31263 8081
rect 31205 8072 31217 8075
rect 30800 8044 31217 8072
rect 30800 8032 30806 8044
rect 31205 8041 31217 8044
rect 31251 8041 31263 8075
rect 31205 8035 31263 8041
rect 27430 8004 27436 8016
rect 27356 7976 27436 8004
rect 27356 7945 27384 7976
rect 27430 7964 27436 7976
rect 27488 7964 27494 8016
rect 29362 7964 29368 8016
rect 29420 8013 29426 8016
rect 29420 8004 29432 8013
rect 29420 7976 29465 8004
rect 29420 7967 29432 7976
rect 29420 7964 29426 7967
rect 27065 7939 27123 7945
rect 27065 7936 27077 7939
rect 26568 7908 27077 7936
rect 26568 7896 26574 7908
rect 27065 7905 27077 7908
rect 27111 7905 27123 7939
rect 27065 7899 27123 7905
rect 27249 7939 27307 7945
rect 27249 7905 27261 7939
rect 27295 7905 27307 7939
rect 27249 7899 27307 7905
rect 27341 7939 27399 7945
rect 27341 7905 27353 7939
rect 27387 7905 27399 7939
rect 27614 7936 27620 7948
rect 27575 7908 27620 7936
rect 27341 7899 27399 7905
rect 27614 7896 27620 7908
rect 27672 7896 27678 7948
rect 30101 7939 30159 7945
rect 30101 7936 30113 7939
rect 27724 7908 30113 7936
rect 26329 7871 26387 7877
rect 26329 7868 26341 7871
rect 25424 7840 26341 7868
rect 26329 7837 26341 7840
rect 26375 7837 26387 7871
rect 26329 7831 26387 7837
rect 27154 7828 27160 7880
rect 27212 7868 27218 7880
rect 27433 7871 27491 7877
rect 27433 7868 27445 7871
rect 27212 7840 27445 7868
rect 27212 7828 27218 7840
rect 27433 7837 27445 7840
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 27724 7800 27752 7908
rect 30101 7905 30113 7908
rect 30147 7905 30159 7939
rect 30101 7899 30159 7905
rect 29641 7871 29699 7877
rect 29641 7837 29653 7871
rect 29687 7837 29699 7871
rect 29641 7831 29699 7837
rect 24228 7772 27752 7800
rect 23934 7732 23940 7744
rect 23216 7704 23940 7732
rect 23934 7692 23940 7704
rect 23992 7692 23998 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 25038 7732 25044 7744
rect 24176 7704 25044 7732
rect 24176 7692 24182 7704
rect 25038 7692 25044 7704
rect 25096 7732 25102 7744
rect 26326 7732 26332 7744
rect 25096 7704 26332 7732
rect 25096 7692 25102 7704
rect 26326 7692 26332 7704
rect 26384 7692 26390 7744
rect 27798 7732 27804 7744
rect 27759 7704 27804 7732
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 28994 7692 29000 7744
rect 29052 7732 29058 7744
rect 29656 7732 29684 7831
rect 29052 7704 29684 7732
rect 29052 7692 29058 7704
rect 1104 7642 32016 7664
rect 1104 7590 6102 7642
rect 6154 7590 6166 7642
rect 6218 7590 6230 7642
rect 6282 7590 6294 7642
rect 6346 7590 6358 7642
rect 6410 7590 16405 7642
rect 16457 7590 16469 7642
rect 16521 7590 16533 7642
rect 16585 7590 16597 7642
rect 16649 7590 16661 7642
rect 16713 7590 26709 7642
rect 26761 7590 26773 7642
rect 26825 7590 26837 7642
rect 26889 7590 26901 7642
rect 26953 7590 26965 7642
rect 27017 7590 32016 7642
rect 1104 7568 32016 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 3510 7528 3516 7540
rect 1811 7500 3516 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 3970 7528 3976 7540
rect 3931 7500 3976 7528
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4706 7528 4712 7540
rect 4667 7500 4712 7528
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 5500 7500 6224 7528
rect 5500 7488 5506 7500
rect 3142 7460 3148 7472
rect 3103 7432 3148 7460
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 3789 7463 3847 7469
rect 3789 7460 3801 7463
rect 3252 7432 3801 7460
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2314 7392 2320 7404
rect 1903 7364 2320 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2608 7392 2774 7400
rect 3050 7392 3056 7404
rect 2547 7372 3056 7392
rect 2547 7364 2636 7372
rect 2746 7364 3056 7372
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3252 7401 3280 7432
rect 3789 7429 3801 7432
rect 3835 7429 3847 7463
rect 5994 7460 6000 7472
rect 3789 7423 3847 7429
rect 3896 7432 6000 7460
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3896 7392 3924 7432
rect 5994 7420 6000 7432
rect 6052 7460 6058 7472
rect 6089 7463 6147 7469
rect 6089 7460 6101 7463
rect 6052 7432 6101 7460
rect 6052 7420 6058 7432
rect 6089 7429 6101 7432
rect 6135 7429 6147 7463
rect 6196 7460 6224 7500
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6604 7500 6837 7528
rect 6604 7488 6610 7500
rect 6825 7497 6837 7500
rect 6871 7528 6883 7531
rect 7282 7528 7288 7540
rect 6871 7500 7288 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 8938 7528 8944 7540
rect 8899 7500 8944 7528
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10778 7528 10784 7540
rect 10284 7500 10784 7528
rect 10284 7488 10290 7500
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 13078 7528 13084 7540
rect 12299 7500 13084 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 14277 7531 14335 7537
rect 14277 7528 14289 7531
rect 13780 7500 14289 7528
rect 13780 7488 13786 7500
rect 14277 7497 14289 7500
rect 14323 7497 14335 7531
rect 14277 7491 14335 7497
rect 6638 7460 6644 7472
rect 6196 7432 6644 7460
rect 6089 7423 6147 7429
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 9582 7460 9588 7472
rect 8904 7432 9588 7460
rect 8904 7420 8910 7432
rect 9582 7420 9588 7432
rect 9640 7460 9646 7472
rect 9640 7432 9720 7460
rect 9640 7420 9646 7432
rect 5350 7392 5356 7404
rect 3237 7355 3295 7361
rect 3436 7364 3924 7392
rect 5311 7364 5356 7392
rect 1394 7284 1400 7336
rect 1452 7324 1458 7336
rect 1949 7327 2007 7333
rect 1949 7324 1961 7327
rect 1452 7296 1961 7324
rect 1452 7284 1458 7296
rect 1949 7293 1961 7296
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 1964 7256 1992 7287
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2464 7296 2605 7324
rect 2464 7284 2470 7296
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 2869 7327 2927 7333
rect 2869 7324 2881 7327
rect 2740 7296 2881 7324
rect 2740 7284 2746 7296
rect 2869 7293 2881 7296
rect 2915 7324 2927 7327
rect 3436 7324 3464 7364
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5460 7364 5672 7392
rect 2915 7296 3464 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 3568 7296 4629 7324
rect 3568 7284 3574 7296
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 5132 7296 5273 7324
rect 5132 7284 5138 7296
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 5261 7287 5319 7293
rect 2774 7256 2780 7268
rect 1964 7228 2780 7256
rect 2774 7216 2780 7228
rect 2832 7256 2838 7268
rect 3970 7265 3976 7268
rect 3957 7259 3976 7265
rect 2832 7228 3280 7256
rect 2832 7216 2838 7228
rect 0 7188 800 7202
rect 1670 7188 1676 7200
rect 0 7160 1676 7188
rect 0 7146 800 7160
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 3252 7188 3280 7228
rect 3957 7225 3969 7259
rect 3957 7219 3976 7225
rect 3970 7216 3976 7219
rect 4028 7216 4034 7268
rect 4157 7259 4215 7265
rect 4157 7225 4169 7259
rect 4203 7225 4215 7259
rect 4157 7219 4215 7225
rect 4172 7188 4200 7219
rect 4246 7216 4252 7268
rect 4304 7256 4310 7268
rect 5460 7256 5488 7364
rect 5644 7333 5672 7364
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8444 7364 9536 7392
rect 8444 7352 8450 7364
rect 9508 7336 9536 7364
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 4304 7228 5488 7256
rect 5552 7256 5580 7287
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 6086 7324 6092 7336
rect 5776 7296 6092 7324
rect 5776 7284 5782 7296
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 6914 7324 6920 7336
rect 6856 7293 6920 7324
rect 6638 7256 6644 7268
rect 5552 7228 5764 7256
rect 6599 7228 6644 7256
rect 4304 7216 4310 7228
rect 5736 7200 5764 7228
rect 6638 7216 6644 7228
rect 6696 7216 6702 7268
rect 6856 7262 6883 7293
rect 6871 7259 6883 7262
rect 6917 7284 6920 7293
rect 6972 7284 6978 7336
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7929 7327 7987 7333
rect 7929 7324 7941 7327
rect 7064 7296 7941 7324
rect 7064 7284 7070 7296
rect 7929 7293 7941 7296
rect 7975 7293 7987 7327
rect 9122 7324 9128 7336
rect 9083 7296 9128 7324
rect 7929 7287 7987 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9306 7324 9312 7336
rect 9267 7296 9312 7324
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 6917 7259 6929 7284
rect 6871 7253 6929 7259
rect 9214 7216 9220 7268
rect 9272 7256 9278 7268
rect 9416 7256 9444 7287
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9692 7333 9720 7432
rect 13998 7420 14004 7472
rect 14056 7460 14062 7472
rect 14292 7460 14320 7491
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 14424 7500 14473 7528
rect 14424 7488 14430 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 14918 7528 14924 7540
rect 14879 7500 14924 7528
rect 14461 7491 14519 7497
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 15160 7500 16129 7528
rect 15160 7488 15166 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16758 7528 16764 7540
rect 16719 7500 16764 7528
rect 16117 7491 16175 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17221 7531 17279 7537
rect 17221 7528 17233 7531
rect 17184 7500 17233 7528
rect 17184 7488 17190 7500
rect 17221 7497 17233 7500
rect 17267 7497 17279 7531
rect 18230 7528 18236 7540
rect 17221 7491 17279 7497
rect 18064 7500 18236 7528
rect 16850 7460 16856 7472
rect 14056 7432 14228 7460
rect 14292 7432 16856 7460
rect 14056 7420 14062 7432
rect 10686 7352 10692 7404
rect 10744 7392 10750 7404
rect 14200 7401 14228 7432
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 17770 7420 17776 7472
rect 17828 7460 17834 7472
rect 18064 7469 18092 7500
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7528 19671 7531
rect 19886 7528 19892 7540
rect 19659 7500 19892 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 22741 7531 22799 7537
rect 22741 7528 22753 7531
rect 22152 7500 22753 7528
rect 22152 7488 22158 7500
rect 22741 7497 22753 7500
rect 22787 7528 22799 7531
rect 23106 7528 23112 7540
rect 22787 7500 23112 7528
rect 22787 7497 22799 7500
rect 22741 7491 22799 7497
rect 23106 7488 23112 7500
rect 23164 7488 23170 7540
rect 24762 7528 24768 7540
rect 24723 7500 24768 7528
rect 24762 7488 24768 7500
rect 24820 7488 24826 7540
rect 25332 7500 29040 7528
rect 18049 7463 18107 7469
rect 17828 7432 17873 7460
rect 17828 7420 17834 7432
rect 18049 7429 18061 7463
rect 18095 7429 18107 7463
rect 18414 7460 18420 7472
rect 18049 7423 18107 7429
rect 18284 7432 18420 7460
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 10744 7364 10977 7392
rect 10744 7352 10750 7364
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 14185 7395 14243 7401
rect 11379 7364 14136 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 9677 7327 9735 7333
rect 9548 7296 9641 7324
rect 9548 7284 9554 7296
rect 9677 7293 9689 7327
rect 9723 7293 9735 7327
rect 10594 7324 10600 7336
rect 10555 7296 10600 7324
rect 9677 7287 9735 7293
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 10778 7324 10784 7336
rect 10739 7296 10784 7324
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11054 7324 11060 7336
rect 10919 7296 11060 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11149 7327 11207 7333
rect 11149 7293 11161 7327
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 9272 7228 9444 7256
rect 9272 7216 9278 7228
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 11164 7256 11192 7287
rect 11790 7284 11796 7336
rect 11848 7324 11854 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11848 7296 11989 7324
rect 11848 7284 11854 7296
rect 11977 7293 11989 7296
rect 12023 7324 12035 7327
rect 12250 7324 12256 7336
rect 12023 7296 12256 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 12345 7327 12403 7333
rect 12345 7293 12357 7327
rect 12391 7324 12403 7327
rect 12526 7324 12532 7336
rect 12391 7296 12532 7324
rect 12391 7293 12403 7296
rect 12345 7287 12403 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13078 7324 13084 7336
rect 12851 7296 13084 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 14108 7333 14136 7364
rect 14185 7361 14197 7395
rect 14231 7361 14243 7395
rect 15286 7392 15292 7404
rect 15247 7364 15292 7392
rect 14185 7355 14243 7361
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 16298 7392 16304 7404
rect 16259 7364 16304 7392
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 16448 7364 16620 7392
rect 16448 7352 16454 7364
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14884 7296 15117 7324
rect 14884 7284 14890 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15378 7324 15384 7336
rect 15339 7296 15384 7324
rect 15105 7287 15163 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 15473 7327 15531 7333
rect 15473 7293 15485 7327
rect 15519 7293 15531 7327
rect 15654 7324 15660 7336
rect 15615 7296 15660 7324
rect 15473 7287 15531 7293
rect 10008 7228 11192 7256
rect 12268 7256 12296 7284
rect 12989 7259 13047 7265
rect 12989 7256 13001 7259
rect 12268 7228 13001 7256
rect 10008 7216 10014 7228
rect 12989 7225 13001 7228
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 15488 7256 15516 7287
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 16592 7333 16620 7364
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17126 7392 17132 7404
rect 17000 7364 17132 7392
rect 17000 7352 17006 7364
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 18064 7392 18092 7423
rect 17236 7364 18092 7392
rect 18141 7395 18199 7401
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7324 16175 7327
rect 16209 7327 16267 7333
rect 16209 7324 16221 7327
rect 16163 7296 16221 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 16209 7293 16221 7296
rect 16255 7293 16267 7327
rect 16209 7287 16267 7293
rect 16485 7327 16543 7333
rect 16485 7293 16497 7327
rect 16531 7293 16543 7327
rect 16485 7287 16543 7293
rect 16577 7327 16635 7333
rect 16577 7293 16589 7327
rect 16623 7293 16635 7327
rect 16577 7287 16635 7293
rect 13964 7228 15516 7256
rect 16500 7256 16528 7287
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 17236 7324 17264 7364
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18284 7392 18312 7432
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 22554 7420 22560 7472
rect 22612 7460 22618 7472
rect 23293 7463 23351 7469
rect 23293 7460 23305 7463
rect 22612 7432 23305 7460
rect 22612 7420 22618 7432
rect 23293 7429 23305 7432
rect 23339 7460 23351 7463
rect 25332 7460 25360 7500
rect 25498 7460 25504 7472
rect 23339 7432 25360 7460
rect 25459 7432 25504 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 25498 7420 25504 7432
rect 25556 7420 25562 7472
rect 29012 7460 29040 7500
rect 29270 7488 29276 7540
rect 29328 7528 29334 7540
rect 29549 7531 29607 7537
rect 29549 7528 29561 7531
rect 29328 7500 29561 7528
rect 29328 7488 29334 7500
rect 29549 7497 29561 7500
rect 29595 7497 29607 7531
rect 29549 7491 29607 7497
rect 30006 7488 30012 7540
rect 30064 7528 30070 7540
rect 30101 7531 30159 7537
rect 30101 7528 30113 7531
rect 30064 7500 30113 7528
rect 30064 7488 30070 7500
rect 30101 7497 30113 7500
rect 30147 7497 30159 7531
rect 30101 7491 30159 7497
rect 30834 7460 30840 7472
rect 29012 7432 30840 7460
rect 30834 7420 30840 7432
rect 30892 7420 30898 7472
rect 18690 7392 18696 7404
rect 18187 7364 18312 7392
rect 18340 7364 18696 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 16816 7296 17264 7324
rect 16816 7284 16822 7296
rect 17402 7284 17408 7336
rect 17460 7324 17466 7336
rect 17954 7324 17960 7336
rect 17460 7302 17632 7324
rect 17460 7296 17816 7302
rect 17915 7296 17960 7324
rect 17460 7284 17466 7296
rect 17604 7274 17816 7296
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7324 18291 7327
rect 18340 7324 18368 7364
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 20346 7392 20352 7404
rect 20307 7364 20352 7392
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 24486 7352 24492 7404
rect 24544 7392 24550 7404
rect 26326 7392 26332 7404
rect 24544 7364 25636 7392
rect 26287 7364 26332 7392
rect 24544 7352 24550 7364
rect 18279 7296 18368 7324
rect 18418 7327 18476 7333
rect 18279 7293 18291 7296
rect 18233 7287 18291 7293
rect 18418 7293 18430 7327
rect 18464 7324 18476 7327
rect 18506 7324 18512 7336
rect 18464 7296 18512 7324
rect 18464 7293 18476 7296
rect 18418 7287 18476 7293
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 19245 7327 19303 7333
rect 19245 7293 19257 7327
rect 19291 7293 19303 7327
rect 19426 7324 19432 7336
rect 19387 7296 19432 7324
rect 19245 7287 19303 7293
rect 16942 7256 16948 7268
rect 16500 7228 16948 7256
rect 13964 7216 13970 7228
rect 15120 7200 15148 7228
rect 16942 7216 16948 7228
rect 17000 7216 17006 7268
rect 17788 7256 17816 7274
rect 19260 7256 19288 7287
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 20073 7327 20131 7333
rect 20073 7324 20085 7327
rect 19518 7296 20085 7324
rect 17788 7228 19288 7256
rect 3252 7160 4200 7188
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5166 7188 5172 7200
rect 4948 7160 5172 7188
rect 4948 7148 4954 7160
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5261 7191 5319 7197
rect 5261 7157 5273 7191
rect 5307 7188 5319 7191
rect 5353 7191 5411 7197
rect 5353 7188 5365 7191
rect 5307 7160 5365 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 5353 7157 5365 7160
rect 5399 7157 5411 7191
rect 5353 7151 5411 7157
rect 5718 7148 5724 7200
rect 5776 7148 5782 7200
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7098 7188 7104 7200
rect 7055 7160 7104 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 8018 7188 8024 7200
rect 7979 7160 8024 7188
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11756 7160 11805 7188
rect 11756 7148 11762 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 13170 7188 13176 7200
rect 13083 7160 13176 7188
rect 11793 7151 11851 7157
rect 13170 7148 13176 7160
rect 13228 7188 13234 7200
rect 13630 7188 13636 7200
rect 13228 7160 13636 7188
rect 13228 7148 13234 7160
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 15102 7148 15108 7200
rect 15160 7148 15166 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 17402 7188 17408 7200
rect 16172 7160 17408 7188
rect 16172 7148 16178 7160
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17494 7148 17500 7200
rect 17552 7188 17558 7200
rect 19518 7188 19546 7296
rect 20073 7293 20085 7296
rect 20119 7293 20131 7327
rect 20073 7287 20131 7293
rect 20438 7284 20444 7336
rect 20496 7324 20502 7336
rect 21361 7327 21419 7333
rect 21361 7324 21373 7327
rect 20496 7296 21373 7324
rect 20496 7284 20502 7296
rect 21361 7293 21373 7296
rect 21407 7324 21419 7327
rect 22370 7324 22376 7336
rect 21407 7296 22376 7324
rect 21407 7293 21419 7296
rect 21361 7287 21419 7293
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 24765 7327 24823 7333
rect 24765 7293 24777 7327
rect 24811 7293 24823 7327
rect 24765 7287 24823 7293
rect 20162 7216 20168 7268
rect 20220 7256 20226 7268
rect 20806 7256 20812 7268
rect 20220 7228 20812 7256
rect 20220 7216 20226 7228
rect 20806 7216 20812 7228
rect 20864 7216 20870 7268
rect 21628 7259 21686 7265
rect 21628 7225 21640 7259
rect 21674 7256 21686 7259
rect 22002 7256 22008 7268
rect 21674 7228 22008 7256
rect 21674 7225 21686 7228
rect 21628 7219 21686 7225
rect 22002 7216 22008 7228
rect 22060 7216 22066 7268
rect 24780 7256 24808 7287
rect 24854 7284 24860 7336
rect 24912 7324 24918 7336
rect 25608 7333 25636 7364
rect 26326 7352 26332 7364
rect 26384 7352 26390 7404
rect 26510 7352 26516 7404
rect 26568 7392 26574 7404
rect 26605 7395 26663 7401
rect 26605 7392 26617 7395
rect 26568 7364 26617 7392
rect 26568 7352 26574 7364
rect 26605 7361 26617 7364
rect 26651 7361 26663 7395
rect 26605 7355 26663 7361
rect 25409 7327 25467 7333
rect 25409 7324 25421 7327
rect 24912 7296 25421 7324
rect 24912 7284 24918 7296
rect 25409 7293 25421 7296
rect 25455 7293 25467 7327
rect 25409 7287 25467 7293
rect 25593 7327 25651 7333
rect 25593 7293 25605 7327
rect 25639 7293 25651 7327
rect 25593 7287 25651 7293
rect 25682 7284 25688 7336
rect 25740 7324 25746 7336
rect 25869 7327 25927 7333
rect 25740 7296 25785 7324
rect 25740 7284 25746 7296
rect 25869 7293 25881 7327
rect 25915 7324 25927 7327
rect 25958 7324 25964 7336
rect 25915 7296 25964 7324
rect 25915 7293 25927 7296
rect 25869 7287 25927 7293
rect 25958 7284 25964 7296
rect 26016 7284 26022 7336
rect 26344 7324 26372 7352
rect 27062 7324 27068 7336
rect 26344 7296 27068 7324
rect 27062 7284 27068 7296
rect 27120 7284 27126 7336
rect 27798 7284 27804 7336
rect 27856 7324 27862 7336
rect 28730 7327 28788 7333
rect 28730 7324 28742 7327
rect 27856 7296 28742 7324
rect 27856 7284 27862 7296
rect 28730 7293 28742 7296
rect 28776 7293 28788 7327
rect 28994 7324 29000 7336
rect 28955 7296 29000 7324
rect 28730 7287 28788 7293
rect 28994 7284 29000 7296
rect 29052 7284 29058 7336
rect 31110 7324 31116 7336
rect 31071 7296 31116 7324
rect 31110 7284 31116 7296
rect 31168 7284 31174 7336
rect 25774 7256 25780 7268
rect 24780 7228 25780 7256
rect 25774 7216 25780 7228
rect 25832 7216 25838 7268
rect 23750 7188 23756 7200
rect 17552 7160 19546 7188
rect 23711 7160 23756 7188
rect 17552 7148 17558 7160
rect 23750 7148 23756 7160
rect 23808 7148 23814 7200
rect 25130 7148 25136 7200
rect 25188 7188 25194 7200
rect 25225 7191 25283 7197
rect 25225 7188 25237 7191
rect 25188 7160 25237 7188
rect 25188 7148 25194 7160
rect 25225 7157 25237 7160
rect 25271 7157 25283 7191
rect 27614 7188 27620 7200
rect 27575 7160 27620 7188
rect 25225 7151 25283 7157
rect 27614 7148 27620 7160
rect 27672 7148 27678 7200
rect 31297 7191 31355 7197
rect 31297 7157 31309 7191
rect 31343 7188 31355 7191
rect 32320 7188 33120 7202
rect 31343 7160 33120 7188
rect 31343 7157 31355 7160
rect 31297 7151 31355 7157
rect 32320 7146 33120 7160
rect 1104 7098 32016 7120
rect 1104 7046 11253 7098
rect 11305 7046 11317 7098
rect 11369 7046 11381 7098
rect 11433 7046 11445 7098
rect 11497 7046 11509 7098
rect 11561 7046 21557 7098
rect 21609 7046 21621 7098
rect 21673 7046 21685 7098
rect 21737 7046 21749 7098
rect 21801 7046 21813 7098
rect 21865 7046 32016 7098
rect 1104 7024 32016 7046
rect 1946 6984 1952 6996
rect 1780 6956 1952 6984
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1673 6851 1731 6857
rect 1673 6848 1685 6851
rect 1636 6820 1685 6848
rect 1636 6808 1642 6820
rect 1673 6817 1685 6820
rect 1719 6817 1731 6851
rect 1780 6848 1808 6956
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 3510 6984 3516 6996
rect 3471 6956 3516 6984
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 5350 6984 5356 6996
rect 5215 6956 5356 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 5718 6984 5724 6996
rect 5460 6956 5724 6984
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 3145 6919 3203 6925
rect 3145 6916 3157 6919
rect 2464 6888 3157 6916
rect 2464 6876 2470 6888
rect 3145 6885 3157 6888
rect 3191 6916 3203 6919
rect 3970 6916 3976 6928
rect 3191 6888 3976 6916
rect 3191 6885 3203 6888
rect 3145 6879 3203 6885
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 5460 6916 5488 6956
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 8018 6984 8024 6996
rect 5868 6956 8024 6984
rect 5868 6944 5874 6956
rect 8018 6944 8024 6956
rect 8076 6944 8082 6996
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 15654 6944 15660 6996
rect 15712 6944 15718 6996
rect 17218 6984 17224 6996
rect 17179 6956 17224 6984
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 20073 6987 20131 6993
rect 20073 6984 20085 6987
rect 18196 6956 20085 6984
rect 18196 6944 18202 6956
rect 20073 6953 20085 6956
rect 20119 6953 20131 6987
rect 22002 6984 22008 6996
rect 21963 6956 22008 6984
rect 20073 6947 20131 6953
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 22922 6944 22928 6996
rect 22980 6984 22986 6996
rect 28350 6984 28356 6996
rect 22980 6956 28356 6984
rect 22980 6944 22986 6956
rect 28350 6944 28356 6956
rect 28408 6944 28414 6996
rect 31110 6944 31116 6996
rect 31168 6984 31174 6996
rect 31297 6987 31355 6993
rect 31297 6984 31309 6987
rect 31168 6956 31309 6984
rect 31168 6944 31174 6956
rect 31297 6953 31309 6956
rect 31343 6953 31355 6987
rect 31297 6947 31355 6953
rect 4120 6888 5488 6916
rect 5552 6888 5764 6916
rect 4120 6876 4126 6888
rect 1836 6851 1894 6857
rect 1836 6848 1848 6851
rect 1780 6820 1848 6848
rect 1673 6811 1731 6817
rect 1836 6817 1848 6820
rect 1882 6848 1894 6851
rect 1882 6817 1900 6848
rect 1836 6811 1900 6817
rect 1872 6712 1900 6811
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 2087 6851 2145 6857
rect 2004 6820 2049 6848
rect 2004 6808 2010 6820
rect 2087 6817 2099 6851
rect 2133 6848 2145 6851
rect 2682 6848 2688 6860
rect 2133 6820 2688 6848
rect 2133 6817 2145 6820
rect 2087 6811 2145 6817
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3016 6820 3188 6848
rect 3016 6808 3022 6820
rect 3160 6792 3188 6820
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 3602 6848 3608 6860
rect 3384 6820 3608 6848
rect 3384 6808 3390 6820
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4212 6820 4445 6848
rect 4212 6808 4218 6820
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 5258 6848 5264 6860
rect 4571 6820 5264 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2498 6780 2504 6792
rect 2363 6752 2504 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 2869 6743 2927 6749
rect 2884 6712 2912 6743
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 4540 6780 4568 6811
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5442 6848 5448 6860
rect 5403 6820 5448 6848
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 5552 6857 5580 6888
rect 5736 6860 5764 6888
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 3200 6752 4568 6780
rect 4709 6783 4767 6789
rect 3200 6740 3206 6752
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5166 6780 5172 6792
rect 4755 6752 5172 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 2958 6712 2964 6724
rect 1872 6684 2544 6712
rect 2884 6684 2964 6712
rect 2516 6656 2544 6684
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 5644 6712 5672 6811
rect 5718 6808 5724 6860
rect 5776 6808 5782 6860
rect 5828 6857 5856 6944
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 10744 6888 11008 6916
rect 10744 6876 10750 6888
rect 5825 6851 5883 6857
rect 5825 6817 5837 6851
rect 5871 6817 5883 6851
rect 5825 6811 5883 6817
rect 7285 6851 7343 6857
rect 7285 6817 7297 6851
rect 7331 6848 7343 6851
rect 8386 6848 8392 6860
rect 7331 6820 8392 6848
rect 7331 6817 7343 6820
rect 7285 6811 7343 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10606 6851 10664 6857
rect 10606 6848 10618 6851
rect 9916 6820 10618 6848
rect 9916 6808 9922 6820
rect 10606 6817 10618 6820
rect 10652 6817 10664 6851
rect 10870 6848 10876 6860
rect 10831 6820 10876 6848
rect 10606 6811 10664 6817
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10980 6848 11008 6888
rect 11532 6888 12020 6916
rect 11532 6848 11560 6888
rect 11698 6848 11704 6860
rect 10980 6820 11560 6848
rect 11659 6820 11704 6848
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 11885 6851 11943 6857
rect 11885 6848 11897 6851
rect 11848 6820 11897 6848
rect 11848 6808 11854 6820
rect 11885 6817 11897 6820
rect 11931 6817 11943 6851
rect 11992 6848 12020 6888
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 14734 6916 14740 6928
rect 12768 6888 14740 6916
rect 12768 6876 12774 6888
rect 14734 6876 14740 6888
rect 14792 6876 14798 6928
rect 15672 6916 15700 6944
rect 15672 6888 15792 6916
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 11992 6820 12081 6848
rect 11885 6811 11943 6817
rect 12069 6817 12081 6820
rect 12115 6817 12127 6851
rect 12250 6848 12256 6860
rect 12211 6820 12256 6848
rect 12069 6811 12127 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13998 6848 14004 6860
rect 14056 6857 14062 6860
rect 12492 6820 12537 6848
rect 13968 6820 14004 6848
rect 12492 6808 12498 6820
rect 13998 6808 14004 6820
rect 14056 6811 14068 6857
rect 15010 6848 15016 6860
rect 14971 6820 15016 6848
rect 14056 6808 14062 6811
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 15197 6851 15255 6857
rect 15197 6848 15209 6851
rect 15160 6820 15209 6848
rect 15160 6808 15166 6820
rect 15197 6817 15209 6820
rect 15243 6817 15255 6851
rect 15378 6848 15384 6860
rect 15339 6820 15384 6848
rect 15197 6811 15255 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 15654 6848 15660 6860
rect 15611 6820 15660 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 15764 6857 15792 6888
rect 15930 6876 15936 6928
rect 15988 6916 15994 6928
rect 23750 6916 23756 6928
rect 15988 6888 23756 6916
rect 15988 6876 15994 6888
rect 23750 6876 23756 6888
rect 23808 6876 23814 6928
rect 24854 6876 24860 6928
rect 24912 6916 24918 6928
rect 24912 6888 26280 6916
rect 24912 6876 24918 6888
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 15838 6848 15844 6860
rect 15795 6820 15844 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16850 6848 16856 6860
rect 16811 6820 16856 6848
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17034 6848 17040 6860
rect 16995 6820 17040 6848
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 18049 6851 18107 6857
rect 18049 6817 18061 6851
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11112 6752 11989 6780
rect 11112 6740 11118 6752
rect 11977 6749 11989 6752
rect 12023 6749 12035 6783
rect 14274 6780 14280 6792
rect 14235 6752 14280 6780
rect 11977 6743 12035 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 15470 6780 15476 6792
rect 15431 6752 15476 6780
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 17862 6780 17868 6792
rect 16172 6752 17868 6780
rect 16172 6740 16178 6752
rect 17862 6740 17868 6752
rect 17920 6780 17926 6792
rect 18064 6780 18092 6811
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 18233 6851 18291 6857
rect 18233 6848 18245 6851
rect 18196 6820 18245 6848
rect 18196 6808 18202 6820
rect 18233 6817 18245 6820
rect 18279 6817 18291 6851
rect 19334 6848 19340 6860
rect 19295 6820 19340 6848
rect 18233 6811 18291 6817
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 19521 6851 19579 6857
rect 19521 6817 19533 6851
rect 19567 6848 19579 6851
rect 19702 6848 19708 6860
rect 19567 6820 19708 6848
rect 19567 6817 19579 6820
rect 19521 6811 19579 6817
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 19981 6851 20039 6857
rect 19981 6817 19993 6851
rect 20027 6817 20039 6851
rect 19981 6811 20039 6817
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 20625 6851 20683 6857
rect 20625 6817 20637 6851
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 17920 6752 18092 6780
rect 18417 6783 18475 6789
rect 17920 6740 17926 6752
rect 18417 6749 18429 6783
rect 18463 6780 18475 6783
rect 18506 6780 18512 6792
rect 18463 6752 18512 6780
rect 18463 6749 18475 6752
rect 18417 6743 18475 6749
rect 18506 6740 18512 6752
rect 18564 6780 18570 6792
rect 19996 6780 20024 6811
rect 18564 6752 20024 6780
rect 18564 6740 18570 6752
rect 4488 6684 5672 6712
rect 4488 6672 4494 6684
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 6086 6712 6092 6724
rect 5868 6684 6092 6712
rect 5868 6672 5874 6684
rect 6086 6672 6092 6684
rect 6144 6712 6150 6724
rect 6365 6715 6423 6721
rect 6365 6712 6377 6715
rect 6144 6684 6377 6712
rect 6144 6672 6150 6684
rect 6365 6681 6377 6684
rect 6411 6681 6423 6715
rect 6365 6675 6423 6681
rect 7742 6672 7748 6724
rect 7800 6712 7806 6724
rect 8573 6715 8631 6721
rect 8573 6712 8585 6715
rect 7800 6684 8585 6712
rect 7800 6672 7806 6684
rect 8573 6681 8585 6684
rect 8619 6681 8631 6715
rect 8573 6675 8631 6681
rect 16298 6672 16304 6724
rect 16356 6712 16362 6724
rect 17586 6712 17592 6724
rect 16356 6684 17592 6712
rect 16356 6672 16362 6684
rect 17586 6672 17592 6684
rect 17644 6712 17650 6724
rect 20180 6712 20208 6811
rect 20640 6712 20668 6811
rect 22094 6808 22100 6860
rect 22152 6848 22158 6860
rect 22189 6851 22247 6857
rect 22189 6848 22201 6851
rect 22152 6820 22201 6848
rect 22152 6808 22158 6820
rect 22189 6817 22201 6820
rect 22235 6817 22247 6851
rect 22189 6811 22247 6817
rect 22278 6808 22284 6860
rect 22336 6848 22342 6860
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 22336 6820 22477 6848
rect 22336 6808 22342 6820
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6817 22615 6851
rect 22557 6811 22615 6817
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6749 22431 6783
rect 22572 6780 22600 6811
rect 22646 6808 22652 6860
rect 22704 6848 22710 6860
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22704 6820 22753 6848
rect 22704 6808 22710 6820
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 22741 6811 22799 6817
rect 23474 6808 23480 6860
rect 23532 6848 23538 6860
rect 23661 6851 23719 6857
rect 23661 6848 23673 6851
rect 23532 6820 23673 6848
rect 23532 6808 23538 6820
rect 23661 6817 23673 6820
rect 23707 6817 23719 6851
rect 23661 6811 23719 6817
rect 24673 6851 24731 6857
rect 24673 6817 24685 6851
rect 24719 6848 24731 6851
rect 24946 6848 24952 6860
rect 24719 6820 24952 6848
rect 24719 6817 24731 6820
rect 24673 6811 24731 6817
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 25130 6848 25136 6860
rect 25091 6820 25136 6848
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 25317 6851 25375 6857
rect 25317 6848 25329 6851
rect 25240 6820 25329 6848
rect 23842 6780 23848 6792
rect 22572 6752 23848 6780
rect 22373 6743 22431 6749
rect 17644 6684 20208 6712
rect 20272 6684 20668 6712
rect 17644 6672 17650 6684
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 5994 6644 6000 6656
rect 4663 6616 6000 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 10134 6644 10140 6656
rect 9732 6616 10140 6644
rect 9732 6604 9738 6616
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 12526 6604 12532 6656
rect 12584 6644 12590 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12584 6616 12909 6644
rect 12584 6604 12590 6616
rect 12897 6613 12909 6616
rect 12943 6644 12955 6647
rect 13538 6644 13544 6656
rect 12943 6616 13544 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 20272 6644 20300 6684
rect 21082 6672 21088 6724
rect 21140 6712 21146 6724
rect 22388 6712 22416 6743
rect 23842 6740 23848 6752
rect 23900 6740 23906 6792
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24854 6780 24860 6792
rect 24627 6752 24860 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24854 6740 24860 6752
rect 24912 6740 24918 6792
rect 22462 6712 22468 6724
rect 21140 6684 22094 6712
rect 22375 6684 22468 6712
rect 21140 6672 21146 6684
rect 20714 6644 20720 6656
rect 15620 6616 20300 6644
rect 20675 6616 20720 6644
rect 15620 6604 15626 6616
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 22066 6644 22094 6684
rect 22462 6672 22468 6684
rect 22520 6712 22526 6724
rect 22922 6712 22928 6724
rect 22520 6684 22928 6712
rect 22520 6672 22526 6684
rect 22922 6672 22928 6684
rect 22980 6672 22986 6724
rect 24305 6715 24363 6721
rect 24305 6681 24317 6715
rect 24351 6712 24363 6715
rect 25240 6712 25268 6820
rect 25317 6817 25329 6820
rect 25363 6817 25375 6851
rect 25590 6848 25596 6860
rect 25551 6820 25596 6848
rect 25317 6811 25375 6817
rect 25590 6808 25596 6820
rect 25648 6808 25654 6860
rect 25774 6848 25780 6860
rect 25735 6820 25780 6848
rect 25774 6808 25780 6820
rect 25832 6808 25838 6860
rect 26252 6857 26280 6888
rect 26237 6851 26295 6857
rect 26237 6817 26249 6851
rect 26283 6817 26295 6851
rect 26237 6811 26295 6817
rect 26510 6808 26516 6860
rect 26568 6848 26574 6860
rect 27157 6851 27215 6857
rect 27157 6848 27169 6851
rect 26568 6820 27169 6848
rect 26568 6808 26574 6820
rect 27157 6817 27169 6820
rect 27203 6817 27215 6851
rect 27157 6811 27215 6817
rect 27341 6851 27399 6857
rect 27341 6817 27353 6851
rect 27387 6848 27399 6851
rect 27614 6848 27620 6860
rect 27387 6820 27620 6848
rect 27387 6817 27399 6820
rect 27341 6811 27399 6817
rect 27614 6808 27620 6820
rect 27672 6808 27678 6860
rect 27709 6851 27767 6857
rect 27709 6817 27721 6851
rect 27755 6848 27767 6851
rect 28442 6848 28448 6860
rect 27755 6820 28448 6848
rect 27755 6817 27767 6820
rect 27709 6811 27767 6817
rect 28442 6808 28448 6820
rect 28500 6808 28506 6860
rect 28997 6851 29055 6857
rect 28997 6817 29009 6851
rect 29043 6848 29055 6851
rect 29086 6848 29092 6860
rect 29043 6820 29092 6848
rect 29043 6817 29055 6820
rect 28997 6811 29055 6817
rect 29086 6808 29092 6820
rect 29144 6808 29150 6860
rect 29270 6808 29276 6860
rect 29328 6848 29334 6860
rect 30561 6851 30619 6857
rect 30561 6848 30573 6851
rect 29328 6820 30573 6848
rect 29328 6808 29334 6820
rect 30561 6817 30573 6820
rect 30607 6817 30619 6851
rect 30561 6811 30619 6817
rect 31113 6851 31171 6857
rect 31113 6817 31125 6851
rect 31159 6848 31171 6851
rect 31294 6848 31300 6860
rect 31159 6820 31300 6848
rect 31159 6817 31171 6820
rect 31113 6811 31171 6817
rect 31294 6808 31300 6820
rect 31352 6808 31358 6860
rect 25498 6780 25504 6792
rect 25459 6752 25504 6780
rect 25498 6740 25504 6752
rect 25556 6740 25562 6792
rect 25608 6780 25636 6808
rect 26329 6783 26387 6789
rect 26329 6780 26341 6783
rect 25608 6752 26341 6780
rect 26329 6749 26341 6752
rect 26375 6749 26387 6783
rect 27430 6780 27436 6792
rect 27391 6752 27436 6780
rect 26329 6743 26387 6749
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 27522 6740 27528 6792
rect 27580 6780 27586 6792
rect 27580 6752 27625 6780
rect 27580 6740 27586 6752
rect 28718 6740 28724 6792
rect 28776 6780 28782 6792
rect 30742 6780 30748 6792
rect 28776 6752 30748 6780
rect 28776 6740 28782 6752
rect 30742 6740 30748 6752
rect 30800 6740 30806 6792
rect 25406 6712 25412 6724
rect 24351 6684 25268 6712
rect 25367 6684 25412 6712
rect 24351 6681 24363 6684
rect 24305 6675 24363 6681
rect 25406 6672 25412 6684
rect 25464 6672 25470 6724
rect 30009 6715 30067 6721
rect 30009 6712 30021 6715
rect 28368 6684 30021 6712
rect 28368 6656 28396 6684
rect 30009 6681 30021 6684
rect 30055 6681 30067 6715
rect 30009 6675 30067 6681
rect 23658 6644 23664 6656
rect 22066 6616 23664 6644
rect 23658 6604 23664 6616
rect 23716 6604 23722 6656
rect 23753 6647 23811 6653
rect 23753 6613 23765 6647
rect 23799 6644 23811 6647
rect 24394 6644 24400 6656
rect 23799 6616 24400 6644
rect 23799 6613 23811 6616
rect 23753 6607 23811 6613
rect 24394 6604 24400 6616
rect 24452 6604 24458 6656
rect 24670 6644 24676 6656
rect 24631 6616 24676 6644
rect 24670 6604 24676 6616
rect 24728 6604 24734 6656
rect 27890 6644 27896 6656
rect 27851 6616 27896 6644
rect 27890 6604 27896 6616
rect 27948 6604 27954 6656
rect 28350 6644 28356 6656
rect 28311 6616 28356 6644
rect 28350 6604 28356 6616
rect 28408 6604 28414 6656
rect 28626 6604 28632 6656
rect 28684 6644 28690 6656
rect 29457 6647 29515 6653
rect 29457 6644 29469 6647
rect 28684 6616 29469 6644
rect 28684 6604 28690 6616
rect 29457 6613 29469 6616
rect 29503 6613 29515 6647
rect 29457 6607 29515 6613
rect 1104 6554 32016 6576
rect 1104 6502 6102 6554
rect 6154 6502 6166 6554
rect 6218 6502 6230 6554
rect 6282 6502 6294 6554
rect 6346 6502 6358 6554
rect 6410 6502 16405 6554
rect 16457 6502 16469 6554
rect 16521 6502 16533 6554
rect 16585 6502 16597 6554
rect 16649 6502 16661 6554
rect 16713 6502 26709 6554
rect 26761 6502 26773 6554
rect 26825 6502 26837 6554
rect 26889 6502 26901 6554
rect 26953 6502 26965 6554
rect 27017 6502 32016 6554
rect 1104 6480 32016 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 2740 6412 2973 6440
rect 2740 6400 2746 6412
rect 2961 6409 2973 6412
rect 3007 6440 3019 6443
rect 3050 6440 3056 6452
rect 3007 6412 3056 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4798 6440 4804 6452
rect 4019 6412 4804 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 5132 6412 5856 6440
rect 5132 6400 5138 6412
rect 1946 6332 1952 6384
rect 2004 6372 2010 6384
rect 2041 6375 2099 6381
rect 2041 6372 2053 6375
rect 2004 6344 2053 6372
rect 2004 6332 2010 6344
rect 2041 6341 2053 6344
rect 2087 6372 2099 6375
rect 4062 6372 4068 6384
rect 2087 6344 4068 6372
rect 2087 6341 2099 6344
rect 2041 6335 2099 6341
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5718 6304 5724 6316
rect 5399 6276 5724 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5828 6304 5856 6412
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 10410 6440 10416 6452
rect 9272 6412 10416 6440
rect 9272 6400 9278 6412
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 11425 6443 11483 6449
rect 11425 6409 11437 6443
rect 11471 6440 11483 6443
rect 11606 6440 11612 6452
rect 11471 6412 11612 6440
rect 11471 6409 11483 6412
rect 11425 6403 11483 6409
rect 11606 6400 11612 6412
rect 11664 6440 11670 6452
rect 11882 6440 11888 6452
rect 11664 6412 11888 6440
rect 11664 6400 11670 6412
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 12308 6412 13277 6440
rect 12308 6400 12314 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 13265 6403 13323 6409
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 14093 6443 14151 6449
rect 14093 6440 14105 6443
rect 14056 6412 14105 6440
rect 14056 6400 14062 6412
rect 14093 6409 14105 6412
rect 14139 6409 14151 6443
rect 14093 6403 14151 6409
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 15933 6443 15991 6449
rect 14608 6412 14688 6440
rect 14608 6400 14614 6412
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 7101 6375 7159 6381
rect 5960 6344 6005 6372
rect 5960 6332 5966 6344
rect 7101 6341 7113 6375
rect 7147 6372 7159 6375
rect 8389 6375 8447 6381
rect 7147 6344 8340 6372
rect 7147 6341 7159 6344
rect 7101 6335 7159 6341
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 5828 6276 6929 6304
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7616 6276 7665 6304
rect 7616 6264 7622 6276
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 8312 6304 8340 6344
rect 8389 6341 8401 6375
rect 8435 6372 8447 6375
rect 10226 6372 10232 6384
rect 8435 6344 10232 6372
rect 8435 6341 8447 6344
rect 8389 6335 8447 6341
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10336 6344 10732 6372
rect 8662 6304 8668 6316
rect 8312 6276 8668 6304
rect 7653 6267 7711 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 10336 6304 10364 6344
rect 9140 6276 10364 6304
rect 10505 6307 10563 6313
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4430 6236 4436 6248
rect 4111 6208 4436 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4430 6196 4436 6208
rect 4488 6236 4494 6248
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4488 6208 4537 6236
rect 4488 6196 4494 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 5074 6236 5080 6248
rect 4755 6208 5080 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 5534 6236 5540 6248
rect 5495 6208 5540 6236
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6052 6208 6653 6236
rect 6052 6196 6058 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7248 6208 7297 6236
rect 7248 6196 7254 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 9140 6245 9168 6276
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10594 6304 10600 6316
rect 10551 6276 10600 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8904 6208 8953 6236
rect 8904 6196 8910 6208
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 9125 6239 9183 6245
rect 9125 6238 9137 6239
rect 8941 6199 8999 6205
rect 9068 6210 9137 6238
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 1857 6171 1915 6177
rect 1857 6168 1869 6171
rect 1728 6140 1869 6168
rect 1728 6128 1734 6140
rect 1857 6137 1869 6140
rect 1903 6137 1915 6171
rect 1857 6131 1915 6137
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 2958 6168 2964 6180
rect 2915 6140 2964 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 5626 6168 5632 6180
rect 4540 6140 5632 6168
rect 4540 6112 4568 6140
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 9068 6168 9096 6210
rect 9125 6205 9137 6210
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9211 6239 9269 6245
rect 9211 6226 9223 6239
rect 9257 6226 9269 6239
rect 9309 6239 9367 6245
rect 9211 6199 9220 6226
rect 9214 6174 9220 6199
rect 9272 6174 9278 6226
rect 9309 6205 9321 6239
rect 9355 6205 9367 6239
rect 9309 6199 9367 6205
rect 8812 6140 9096 6168
rect 9324 6168 9352 6199
rect 9490 6196 9496 6248
rect 9548 6245 9554 6248
rect 9548 6239 9562 6245
rect 9550 6236 9562 6239
rect 9677 6239 9735 6245
rect 9550 6208 9593 6236
rect 9550 6205 9562 6208
rect 9548 6199 9562 6205
rect 9677 6205 9689 6239
rect 9723 6234 9735 6239
rect 9858 6234 9864 6248
rect 9723 6206 9864 6234
rect 9723 6205 9735 6206
rect 9677 6199 9735 6205
rect 9548 6196 9554 6199
rect 9858 6196 9864 6206
rect 9916 6196 9922 6248
rect 10134 6236 10140 6248
rect 10095 6208 10140 6236
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 9398 6168 9404 6180
rect 9324 6140 9404 6168
rect 8812 6128 8818 6140
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 10042 6128 10048 6180
rect 10100 6168 10106 6180
rect 10336 6168 10364 6199
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 10704 6245 10732 6344
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 12400 6276 14565 6304
rect 12400 6264 12406 6276
rect 14553 6273 14565 6276
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 10689 6239 10747 6245
rect 10468 6208 10513 6236
rect 10468 6196 10474 6208
rect 10689 6205 10701 6239
rect 10735 6205 10747 6239
rect 10689 6199 10747 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 12710 6236 12716 6248
rect 12671 6208 12716 6236
rect 12437 6199 12495 6205
rect 10100 6140 10364 6168
rect 12452 6168 12480 6199
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 12860 6208 13185 6236
rect 12860 6196 12866 6208
rect 13173 6205 13185 6208
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 13596 6208 14289 6236
rect 13596 6196 13602 6208
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14660 6245 14688 6412
rect 15933 6409 15945 6443
rect 15979 6440 15991 6443
rect 16114 6440 16120 6452
rect 15979 6412 16120 6440
rect 15979 6409 15991 6412
rect 15933 6403 15991 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 16577 6443 16635 6449
rect 16577 6409 16589 6443
rect 16623 6440 16635 6443
rect 16850 6440 16856 6452
rect 16623 6412 16856 6440
rect 16623 6409 16635 6412
rect 16577 6403 16635 6409
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17034 6400 17040 6452
rect 17092 6440 17098 6452
rect 17497 6443 17555 6449
rect 17092 6412 17448 6440
rect 17092 6400 17098 6412
rect 17310 6372 17316 6384
rect 16960 6344 17316 6372
rect 16960 6304 16988 6344
rect 17310 6332 17316 6344
rect 17368 6332 17374 6384
rect 16684 6276 16988 6304
rect 16684 6245 16712 6276
rect 14461 6239 14519 6245
rect 14461 6236 14473 6239
rect 14424 6208 14473 6236
rect 14424 6196 14430 6208
rect 14461 6205 14473 6208
rect 14507 6205 14519 6239
rect 14461 6199 14519 6205
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16669 6239 16727 6245
rect 16669 6205 16681 6239
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 12618 6168 12624 6180
rect 12452 6140 12624 6168
rect 10100 6128 10106 6140
rect 12618 6128 12624 6140
rect 12676 6168 12682 6180
rect 13446 6168 13452 6180
rect 12676 6140 13452 6168
rect 12676 6128 12682 6140
rect 13446 6128 13452 6140
rect 13504 6168 13510 6180
rect 14844 6168 14872 6199
rect 13504 6140 14872 6168
rect 16040 6168 16068 6199
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 17129 6239 17187 6245
rect 17129 6236 17141 6239
rect 16908 6208 17141 6236
rect 16908 6196 16914 6208
rect 17129 6205 17141 6208
rect 17175 6205 17187 6239
rect 17420 6236 17448 6412
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17586 6440 17592 6452
rect 17543 6412 17592 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 18693 6443 18751 6449
rect 18693 6409 18705 6443
rect 18739 6440 18751 6443
rect 21266 6440 21272 6452
rect 18739 6412 21272 6440
rect 18739 6409 18751 6412
rect 18693 6403 18751 6409
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 21910 6400 21916 6452
rect 21968 6440 21974 6452
rect 23106 6440 23112 6452
rect 21968 6412 23112 6440
rect 21968 6400 21974 6412
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 27062 6440 27068 6452
rect 27023 6412 27068 6440
rect 27062 6400 27068 6412
rect 27120 6400 27126 6452
rect 28350 6440 28356 6452
rect 27264 6412 28356 6440
rect 20254 6332 20260 6384
rect 20312 6372 20318 6384
rect 20717 6375 20775 6381
rect 20717 6372 20729 6375
rect 20312 6344 20729 6372
rect 20312 6332 20318 6344
rect 20717 6341 20729 6344
rect 20763 6341 20775 6375
rect 20717 6335 20775 6341
rect 23658 6332 23664 6384
rect 23716 6372 23722 6384
rect 27264 6372 27292 6412
rect 28350 6400 28356 6412
rect 28408 6440 28414 6452
rect 28718 6440 28724 6452
rect 28408 6412 28724 6440
rect 28408 6400 28414 6412
rect 28718 6400 28724 6412
rect 28776 6400 28782 6452
rect 29270 6400 29276 6452
rect 29328 6440 29334 6452
rect 29549 6443 29607 6449
rect 29549 6440 29561 6443
rect 29328 6412 29561 6440
rect 29328 6400 29334 6412
rect 29549 6409 29561 6412
rect 29595 6409 29607 6443
rect 30098 6440 30104 6452
rect 30059 6412 30104 6440
rect 29549 6403 29607 6409
rect 30098 6400 30104 6412
rect 30156 6400 30162 6452
rect 30929 6443 30987 6449
rect 30929 6409 30941 6443
rect 30975 6440 30987 6443
rect 31018 6440 31024 6452
rect 30975 6412 31024 6440
rect 30975 6409 30987 6412
rect 30929 6403 30987 6409
rect 31018 6400 31024 6412
rect 31076 6440 31082 6452
rect 31570 6440 31576 6452
rect 31076 6412 31576 6440
rect 31076 6400 31082 6412
rect 31570 6400 31576 6412
rect 31628 6400 31634 6452
rect 23716 6344 27292 6372
rect 23716 6332 23722 6344
rect 27338 6332 27344 6384
rect 27396 6372 27402 6384
rect 27522 6372 27528 6384
rect 27396 6344 27528 6372
rect 27396 6332 27402 6344
rect 27522 6332 27528 6344
rect 27580 6332 27586 6384
rect 19886 6304 19892 6316
rect 19847 6276 19892 6304
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 20898 6264 20904 6316
rect 20956 6304 20962 6316
rect 21910 6304 21916 6316
rect 20956 6276 21916 6304
rect 20956 6264 20962 6276
rect 21910 6264 21916 6276
rect 21968 6304 21974 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 21968 6276 22109 6304
rect 21968 6264 21974 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22278 6264 22284 6316
rect 22336 6304 22342 6316
rect 22830 6304 22836 6316
rect 22336 6276 22836 6304
rect 22336 6264 22342 6276
rect 22830 6264 22836 6276
rect 22888 6264 22894 6316
rect 23750 6304 23756 6316
rect 23711 6276 23756 6304
rect 23750 6264 23756 6276
rect 23808 6304 23814 6316
rect 24397 6307 24455 6313
rect 24397 6304 24409 6307
rect 23808 6276 24409 6304
rect 23808 6264 23814 6276
rect 24397 6273 24409 6276
rect 24443 6273 24455 6307
rect 24397 6267 24455 6273
rect 26418 6264 26424 6316
rect 26476 6304 26482 6316
rect 26513 6307 26571 6313
rect 26513 6304 26525 6307
rect 26476 6276 26525 6304
rect 26476 6264 26482 6276
rect 26513 6273 26525 6276
rect 26559 6304 26571 6307
rect 27154 6304 27160 6316
rect 26559 6276 27160 6304
rect 26559 6273 26571 6276
rect 26513 6267 26571 6273
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 17420 6208 17969 6236
rect 17129 6199 17187 6205
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 19242 6196 19248 6248
rect 19300 6236 19306 6248
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 19300 6208 19533 6236
rect 19300 6196 19306 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 19705 6239 19763 6245
rect 19705 6205 19717 6239
rect 19751 6205 19763 6239
rect 19705 6199 19763 6205
rect 16758 6168 16764 6180
rect 16040 6140 16764 6168
rect 13504 6128 13510 6140
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 17313 6171 17371 6177
rect 17313 6137 17325 6171
rect 17359 6168 17371 6171
rect 17770 6168 17776 6180
rect 17359 6140 17776 6168
rect 17359 6137 17371 6140
rect 17313 6131 17371 6137
rect 17770 6128 17776 6140
rect 17828 6168 17834 6180
rect 18049 6171 18107 6177
rect 18049 6168 18061 6171
rect 17828 6140 18061 6168
rect 17828 6128 17834 6140
rect 18049 6137 18061 6140
rect 18095 6137 18107 6171
rect 18049 6131 18107 6137
rect 19058 6128 19064 6180
rect 19116 6168 19122 6180
rect 19720 6168 19748 6199
rect 19794 6196 19800 6248
rect 19852 6236 19858 6248
rect 20073 6239 20131 6245
rect 19852 6208 19897 6236
rect 19852 6196 19858 6208
rect 20073 6205 20085 6239
rect 20119 6236 20131 6239
rect 21082 6236 21088 6248
rect 20119 6208 21088 6236
rect 20119 6205 20131 6208
rect 20073 6199 20131 6205
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 21821 6239 21879 6245
rect 21821 6205 21833 6239
rect 21867 6236 21879 6239
rect 22002 6236 22008 6248
rect 21867 6208 22008 6236
rect 21867 6205 21879 6208
rect 21821 6199 21879 6205
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 22554 6236 22560 6248
rect 22515 6208 22560 6236
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 22741 6239 22799 6245
rect 22741 6205 22753 6239
rect 22787 6205 22799 6239
rect 22922 6236 22928 6248
rect 22883 6208 22928 6236
rect 22741 6199 22799 6205
rect 20898 6168 20904 6180
rect 19116 6140 19748 6168
rect 19812 6140 20904 6168
rect 19116 6128 19122 6140
rect 4522 6060 4528 6112
rect 4580 6060 4586 6112
rect 4617 6103 4675 6109
rect 4617 6069 4629 6103
rect 4663 6100 4675 6103
rect 5442 6100 5448 6112
rect 4663 6072 5448 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 8076 6072 10885 6100
rect 8076 6060 8082 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 15286 6100 15292 6112
rect 15247 6072 15292 6100
rect 10873 6063 10931 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 19812 6100 19840 6140
rect 20898 6128 20904 6140
rect 20956 6168 20962 6180
rect 22462 6168 22468 6180
rect 20956 6140 22468 6168
rect 20956 6128 20962 6140
rect 22462 6128 22468 6140
rect 22520 6128 22526 6180
rect 22756 6168 22784 6199
rect 22922 6196 22928 6208
rect 22980 6196 22986 6248
rect 23109 6239 23167 6245
rect 23109 6205 23121 6239
rect 23155 6236 23167 6239
rect 23842 6236 23848 6248
rect 23155 6208 23848 6236
rect 23155 6205 23167 6208
rect 23109 6199 23167 6205
rect 23842 6196 23848 6208
rect 23900 6196 23906 6248
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 24673 6239 24731 6245
rect 24673 6236 24685 6239
rect 24636 6208 24685 6236
rect 24636 6196 24642 6208
rect 24673 6205 24685 6208
rect 24719 6205 24731 6239
rect 24673 6199 24731 6205
rect 26237 6239 26295 6245
rect 26237 6205 26249 6239
rect 26283 6205 26295 6239
rect 26237 6199 26295 6205
rect 23474 6168 23480 6180
rect 22756 6140 23480 6168
rect 23474 6128 23480 6140
rect 23532 6128 23538 6180
rect 24762 6128 24768 6180
rect 24820 6168 24826 6180
rect 26142 6168 26148 6180
rect 24820 6140 26148 6168
rect 24820 6128 24826 6140
rect 26142 6128 26148 6140
rect 26200 6128 26206 6180
rect 26252 6168 26280 6199
rect 26326 6196 26332 6248
rect 26384 6236 26390 6248
rect 26602 6236 26608 6248
rect 26384 6208 26429 6236
rect 26563 6208 26608 6236
rect 26384 6196 26390 6208
rect 26602 6196 26608 6208
rect 26660 6196 26666 6248
rect 27522 6196 27528 6248
rect 27580 6236 27586 6248
rect 27890 6245 27896 6248
rect 27617 6239 27675 6245
rect 27617 6236 27629 6239
rect 27580 6208 27629 6236
rect 27580 6196 27586 6208
rect 27617 6205 27629 6208
rect 27663 6205 27675 6239
rect 27884 6236 27896 6245
rect 27851 6208 27896 6236
rect 27617 6199 27675 6205
rect 27884 6199 27896 6208
rect 27890 6196 27896 6199
rect 27948 6196 27954 6248
rect 28350 6168 28356 6180
rect 26252 6140 28356 6168
rect 28350 6128 28356 6140
rect 28408 6128 28414 6180
rect 16724 6072 19840 6100
rect 16724 6060 16730 6072
rect 20162 6060 20168 6112
rect 20220 6100 20226 6112
rect 20257 6103 20315 6109
rect 20257 6100 20269 6103
rect 20220 6072 20269 6100
rect 20220 6060 20226 6072
rect 20257 6069 20269 6072
rect 20303 6069 20315 6103
rect 23290 6100 23296 6112
rect 23251 6072 23296 6100
rect 20257 6063 20315 6069
rect 23290 6060 23296 6072
rect 23348 6060 23354 6112
rect 26053 6103 26111 6109
rect 26053 6069 26065 6103
rect 26099 6100 26111 6103
rect 26418 6100 26424 6112
rect 26099 6072 26424 6100
rect 26099 6069 26111 6072
rect 26053 6063 26111 6069
rect 26418 6060 26424 6072
rect 26476 6060 26482 6112
rect 28442 6060 28448 6112
rect 28500 6100 28506 6112
rect 28997 6103 29055 6109
rect 28997 6100 29009 6103
rect 28500 6072 29009 6100
rect 28500 6060 28506 6072
rect 28997 6069 29009 6072
rect 29043 6069 29055 6103
rect 28997 6063 29055 6069
rect 1104 6010 32016 6032
rect 1104 5958 11253 6010
rect 11305 5958 11317 6010
rect 11369 5958 11381 6010
rect 11433 5958 11445 6010
rect 11497 5958 11509 6010
rect 11561 5958 21557 6010
rect 21609 5958 21621 6010
rect 21673 5958 21685 6010
rect 21737 5958 21749 6010
rect 21801 5958 21813 6010
rect 21865 5958 32016 6010
rect 1104 5936 32016 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 2406 5896 2412 5908
rect 1627 5868 2412 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2832 5868 2881 5896
rect 2832 5856 2838 5868
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 3234 5856 3240 5908
rect 3292 5896 3298 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3292 5868 3433 5896
rect 3292 5856 3298 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 5166 5896 5172 5908
rect 5127 5868 5172 5896
rect 3421 5859 3479 5865
rect 2222 5828 2228 5840
rect 1504 5800 2228 5828
rect 1504 5769 1532 5800
rect 2222 5788 2228 5800
rect 2280 5788 2286 5840
rect 3436 5828 3464 5859
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 7190 5896 7196 5908
rect 5500 5868 6408 5896
rect 7151 5868 7196 5896
rect 5500 5856 5506 5868
rect 3436 5800 4476 5828
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5729 1547 5763
rect 1489 5723 1547 5729
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1636 5732 1685 5760
rect 1636 5720 1642 5732
rect 1673 5729 1685 5732
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 2498 5760 2504 5772
rect 2363 5732 2504 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 2958 5760 2964 5772
rect 2919 5732 2964 5760
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 4448 5769 4476 5800
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 4856 5800 5693 5828
rect 4856 5788 4862 5800
rect 5665 5772 5693 5800
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5729 4215 5763
rect 4157 5723 4215 5729
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 2130 5584 2136 5636
rect 2188 5624 2194 5636
rect 3142 5624 3148 5636
rect 2188 5596 3148 5624
rect 2188 5584 2194 5596
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 4172 5624 4200 5723
rect 4522 5720 4528 5772
rect 4580 5760 4586 5772
rect 4709 5763 4767 5769
rect 4580 5732 4625 5760
rect 4580 5720 4586 5732
rect 4709 5729 4721 5763
rect 4755 5760 4767 5763
rect 4982 5760 4988 5772
rect 4755 5732 4988 5760
rect 4755 5729 4767 5732
rect 4709 5723 4767 5729
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 5445 5763 5503 5769
rect 5445 5760 5457 5763
rect 5408 5732 5457 5760
rect 5408 5720 5414 5732
rect 5445 5729 5457 5732
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 5550 5763 5608 5769
rect 5550 5729 5562 5763
rect 5596 5729 5608 5763
rect 5550 5723 5608 5729
rect 5650 5766 5708 5772
rect 6380 5769 6408 5868
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8812 5868 9137 5896
rect 8812 5856 8818 5868
rect 9125 5865 9137 5868
rect 9171 5896 9183 5899
rect 9214 5896 9220 5908
rect 9171 5868 9220 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 10965 5899 11023 5905
rect 9784 5868 10548 5896
rect 6730 5828 6736 5840
rect 6656 5800 6736 5828
rect 6656 5769 6684 5800
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 8018 5837 8024 5840
rect 8012 5828 8024 5837
rect 7979 5800 8024 5828
rect 8012 5791 8024 5800
rect 8018 5788 8024 5791
rect 8076 5788 8082 5840
rect 8662 5788 8668 5840
rect 8720 5828 8726 5840
rect 9784 5828 9812 5868
rect 8720 5800 9812 5828
rect 8720 5788 8726 5800
rect 9858 5788 9864 5840
rect 9916 5828 9922 5840
rect 10520 5828 10548 5868
rect 10965 5865 10977 5899
rect 11011 5896 11023 5899
rect 12066 5896 12072 5908
rect 11011 5868 12072 5896
rect 11011 5865 11023 5868
rect 10965 5859 11023 5865
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 16666 5896 16672 5908
rect 12176 5868 16672 5896
rect 12176 5828 12204 5868
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 16761 5899 16819 5905
rect 16761 5865 16773 5899
rect 16807 5896 16819 5899
rect 16850 5896 16856 5908
rect 16807 5868 16856 5896
rect 16807 5865 16819 5868
rect 16761 5859 16819 5865
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17862 5896 17868 5908
rect 17460 5868 17868 5896
rect 17460 5856 17466 5868
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 19058 5896 19064 5908
rect 19019 5868 19064 5896
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 21910 5856 21916 5908
rect 21968 5896 21974 5908
rect 22097 5899 22155 5905
rect 22097 5896 22109 5899
rect 21968 5868 22109 5896
rect 21968 5856 21974 5868
rect 22097 5865 22109 5868
rect 22143 5865 22155 5899
rect 22097 5859 22155 5865
rect 22649 5899 22707 5905
rect 22649 5865 22661 5899
rect 22695 5896 22707 5899
rect 23842 5896 23848 5908
rect 22695 5868 23848 5896
rect 22695 5865 22707 5868
rect 22649 5859 22707 5865
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 24486 5896 24492 5908
rect 24447 5868 24492 5896
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 25406 5856 25412 5908
rect 25464 5896 25470 5908
rect 25685 5899 25743 5905
rect 25685 5896 25697 5899
rect 25464 5868 25697 5896
rect 25464 5856 25470 5868
rect 25685 5865 25697 5868
rect 25731 5865 25743 5899
rect 26510 5896 26516 5908
rect 25685 5859 25743 5865
rect 25792 5868 26516 5896
rect 15286 5828 15292 5840
rect 9916 5800 10456 5828
rect 10520 5800 12204 5828
rect 13832 5800 15292 5828
rect 9916 5788 9922 5800
rect 5650 5732 5662 5766
rect 5696 5732 5708 5766
rect 5650 5726 5708 5732
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5729 6699 5763
rect 7098 5760 7104 5772
rect 7059 5732 7104 5760
rect 6641 5723 6699 5729
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4614 5692 4620 5704
rect 4387 5664 4620 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5561 5692 5589 5723
rect 5368 5664 5589 5692
rect 5368 5636 5396 5664
rect 4172 5596 5212 5624
rect 5184 5568 5212 5596
rect 5350 5584 5356 5636
rect 5408 5584 5414 5636
rect 5828 5624 5856 5723
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7742 5760 7748 5772
rect 7703 5732 7748 5760
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 9585 5763 9643 5769
rect 9585 5729 9597 5763
rect 9631 5729 9643 5763
rect 9585 5723 9643 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 9950 5760 9956 5772
rect 9723 5732 9956 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6733 5695 6791 5701
rect 6733 5692 6745 5695
rect 6052 5664 6745 5692
rect 6052 5652 6058 5664
rect 6733 5661 6745 5664
rect 6779 5692 6791 5695
rect 6914 5692 6920 5704
rect 6779 5664 6920 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 9600 5692 9628 5723
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10428 5769 10456 5800
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5729 10287 5763
rect 10229 5723 10287 5729
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 10686 5760 10692 5772
rect 10643 5732 10692 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 10042 5692 10048 5704
rect 9180 5664 10048 5692
rect 9180 5652 9186 5664
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 7006 5624 7012 5636
rect 5828 5596 7012 5624
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 4062 5556 4068 5568
rect 4019 5528 4068 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 5828 5556 5856 5596
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 10244 5624 10272 5723
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11146 5760 11152 5772
rect 10827 5732 11152 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 11238 5720 11244 5772
rect 11296 5760 11302 5772
rect 11609 5763 11667 5769
rect 11609 5760 11621 5763
rect 11296 5732 11621 5760
rect 11296 5720 11302 5732
rect 11609 5729 11621 5732
rect 11655 5760 11667 5763
rect 13832 5760 13860 5800
rect 15286 5788 15292 5800
rect 15344 5788 15350 5840
rect 16945 5831 17003 5837
rect 16945 5797 16957 5831
rect 16991 5828 17003 5831
rect 16991 5800 17816 5828
rect 16991 5797 17003 5800
rect 16945 5791 17003 5797
rect 17788 5772 17816 5800
rect 13998 5760 14004 5772
rect 14056 5769 14062 5772
rect 11655 5732 13860 5760
rect 13968 5732 14004 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 13998 5720 14004 5732
rect 14056 5723 14068 5769
rect 15197 5763 15255 5769
rect 15197 5729 15209 5763
rect 15243 5729 15255 5763
rect 15470 5760 15476 5772
rect 15431 5732 15476 5760
rect 15197 5723 15255 5729
rect 14056 5720 14062 5723
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5692 10563 5695
rect 11054 5692 11060 5704
rect 10551 5664 11060 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 12342 5692 12348 5704
rect 11931 5664 12348 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 14274 5692 14280 5704
rect 14235 5664 14280 5692
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 15212 5624 15240 5723
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 15562 5720 15568 5772
rect 15620 5760 15626 5772
rect 15749 5763 15807 5769
rect 15620 5732 15665 5760
rect 15620 5720 15626 5732
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 15838 5760 15844 5772
rect 15795 5732 15844 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5760 17187 5763
rect 17310 5760 17316 5772
rect 17175 5732 17316 5760
rect 17175 5729 17187 5732
rect 17129 5723 17187 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17770 5760 17776 5772
rect 17731 5732 17776 5760
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 18141 5763 18199 5769
rect 18141 5729 18153 5763
rect 18187 5760 18199 5763
rect 19076 5760 19104 5856
rect 23290 5788 23296 5840
rect 23348 5828 23354 5840
rect 23762 5831 23820 5837
rect 23762 5828 23774 5831
rect 23348 5800 23774 5828
rect 23348 5788 23354 5800
rect 23762 5797 23774 5800
rect 23808 5797 23820 5831
rect 23762 5791 23820 5797
rect 24394 5788 24400 5840
rect 24452 5828 24458 5840
rect 24452 5800 25084 5828
rect 24452 5788 24458 5800
rect 18187 5732 19104 5760
rect 18187 5729 18199 5732
rect 18141 5723 18199 5729
rect 19610 5720 19616 5772
rect 19668 5760 19674 5772
rect 20174 5763 20232 5769
rect 20174 5760 20186 5763
rect 19668 5732 20186 5760
rect 19668 5720 19674 5732
rect 20174 5729 20186 5732
rect 20220 5729 20232 5763
rect 21082 5760 21088 5772
rect 21043 5732 21088 5760
rect 20174 5723 20232 5729
rect 21082 5720 21088 5732
rect 21140 5720 21146 5772
rect 23934 5720 23940 5772
rect 23992 5760 23998 5772
rect 24029 5763 24087 5769
rect 24029 5760 24041 5763
rect 23992 5732 24041 5760
rect 23992 5720 23998 5732
rect 24029 5729 24041 5732
rect 24075 5729 24087 5763
rect 24670 5760 24676 5772
rect 24631 5732 24676 5760
rect 24029 5723 24087 5729
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 24762 5720 24768 5772
rect 24820 5760 24826 5772
rect 25056 5769 25084 5800
rect 24949 5763 25007 5769
rect 24949 5760 24961 5763
rect 24820 5732 24961 5760
rect 24820 5720 24826 5732
rect 24949 5729 24961 5732
rect 24995 5729 25007 5763
rect 24949 5723 25007 5729
rect 25041 5763 25099 5769
rect 25041 5729 25053 5763
rect 25087 5729 25099 5763
rect 25222 5760 25228 5772
rect 25183 5732 25228 5760
rect 25041 5723 25099 5729
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 25792 5760 25820 5868
rect 26510 5856 26516 5868
rect 26568 5856 26574 5908
rect 26602 5856 26608 5908
rect 26660 5896 26666 5908
rect 27709 5899 27767 5905
rect 27709 5896 27721 5899
rect 26660 5868 27721 5896
rect 26660 5856 26666 5868
rect 27709 5865 27721 5868
rect 27755 5865 27767 5899
rect 28350 5896 28356 5908
rect 28311 5868 28356 5896
rect 27709 5859 27767 5865
rect 28350 5856 28356 5868
rect 28408 5856 28414 5908
rect 28997 5899 29055 5905
rect 28997 5865 29009 5899
rect 29043 5896 29055 5899
rect 29270 5896 29276 5908
rect 29043 5868 29276 5896
rect 29043 5865 29055 5868
rect 28997 5859 29055 5865
rect 29270 5856 29276 5868
rect 29328 5856 29334 5908
rect 30558 5896 30564 5908
rect 30519 5868 30564 5896
rect 30558 5856 30564 5868
rect 30616 5856 30622 5908
rect 31110 5896 31116 5908
rect 31071 5868 31116 5896
rect 31110 5856 31116 5868
rect 31168 5856 31174 5908
rect 25869 5763 25927 5769
rect 25869 5760 25881 5763
rect 25792 5732 25881 5760
rect 25869 5729 25881 5732
rect 25915 5729 25927 5763
rect 26050 5760 26056 5772
rect 25869 5723 25927 5729
rect 25973 5732 26056 5760
rect 15378 5692 15384 5704
rect 15339 5664 15384 5692
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15654 5624 15660 5636
rect 10244 5596 13400 5624
rect 15212 5596 15660 5624
rect 5224 5528 5856 5556
rect 5224 5516 5230 5528
rect 10226 5516 10232 5568
rect 10284 5556 10290 5568
rect 10962 5556 10968 5568
rect 10284 5528 10968 5556
rect 10284 5516 10290 5528
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12860 5528 12909 5556
rect 12860 5516 12866 5528
rect 12897 5525 12909 5528
rect 12943 5525 12955 5559
rect 13372 5556 13400 5596
rect 15654 5584 15660 5596
rect 15712 5584 15718 5636
rect 14550 5556 14556 5568
rect 13372 5528 14556 5556
rect 12897 5519 12955 5525
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 15010 5556 15016 5568
rect 14971 5528 15016 5556
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 17328 5556 17356 5720
rect 17402 5652 17408 5704
rect 17460 5692 17466 5704
rect 18598 5692 18604 5704
rect 17460 5664 18604 5692
rect 17460 5652 17466 5664
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 20438 5692 20444 5704
rect 20399 5664 20444 5692
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 21450 5652 21456 5704
rect 21508 5692 21514 5704
rect 22278 5692 22284 5704
rect 21508 5664 22284 5692
rect 21508 5652 21514 5664
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5692 24915 5695
rect 25973 5692 26001 5732
rect 26050 5720 26056 5732
rect 26108 5720 26114 5772
rect 26249 5761 26307 5767
rect 26249 5727 26261 5761
rect 26295 5727 26307 5761
rect 26249 5721 26307 5727
rect 26151 5692 26157 5704
rect 24903 5664 26001 5692
rect 26112 5664 26157 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 26151 5652 26157 5664
rect 26209 5652 26215 5704
rect 26264 5692 26292 5721
rect 26418 5720 26424 5772
rect 26476 5760 26482 5772
rect 26476 5732 26521 5760
rect 26476 5720 26482 5732
rect 26602 5720 26608 5772
rect 26660 5760 26666 5772
rect 27157 5763 27215 5769
rect 27157 5760 27169 5763
rect 26660 5732 27169 5760
rect 26660 5720 26666 5732
rect 27157 5729 27169 5732
rect 27203 5729 27215 5763
rect 27614 5760 27620 5772
rect 27575 5732 27620 5760
rect 27157 5723 27215 5729
rect 27614 5720 27620 5732
rect 27672 5720 27678 5772
rect 28442 5760 28448 5772
rect 28355 5732 28448 5760
rect 28442 5720 28448 5732
rect 28500 5720 28506 5772
rect 27065 5695 27123 5701
rect 27065 5692 27077 5695
rect 26264 5664 27077 5692
rect 27065 5661 27077 5664
rect 27111 5661 27123 5695
rect 27065 5655 27123 5661
rect 27246 5652 27252 5704
rect 27304 5692 27310 5704
rect 28460 5692 28488 5720
rect 27304 5664 28488 5692
rect 27304 5652 27310 5664
rect 17589 5627 17647 5633
rect 17589 5593 17601 5627
rect 17635 5624 17647 5627
rect 17954 5624 17960 5636
rect 17635 5596 17960 5624
rect 17635 5593 17647 5596
rect 17589 5587 17647 5593
rect 17954 5584 17960 5596
rect 18012 5584 18018 5636
rect 29457 5627 29515 5633
rect 29457 5624 29469 5627
rect 20824 5596 22094 5624
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 17328 5528 17785 5556
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 17773 5519 17831 5525
rect 18046 5516 18052 5568
rect 18104 5556 18110 5568
rect 20824 5556 20852 5596
rect 20990 5556 20996 5568
rect 18104 5528 20852 5556
rect 20951 5528 20996 5556
rect 18104 5516 18110 5528
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 22066 5556 22094 5596
rect 25056 5596 29469 5624
rect 25056 5556 25084 5596
rect 29457 5593 29469 5596
rect 29503 5624 29515 5627
rect 30009 5627 30067 5633
rect 30009 5624 30021 5627
rect 29503 5596 30021 5624
rect 29503 5593 29515 5596
rect 29457 5587 29515 5593
rect 30009 5593 30021 5596
rect 30055 5593 30067 5627
rect 30009 5587 30067 5593
rect 22066 5528 25084 5556
rect 25222 5516 25228 5568
rect 25280 5556 25286 5568
rect 30098 5556 30104 5568
rect 25280 5528 30104 5556
rect 25280 5516 25286 5528
rect 30098 5516 30104 5528
rect 30156 5516 30162 5568
rect 1104 5466 32016 5488
rect 1104 5414 6102 5466
rect 6154 5414 6166 5466
rect 6218 5414 6230 5466
rect 6282 5414 6294 5466
rect 6346 5414 6358 5466
rect 6410 5414 16405 5466
rect 16457 5414 16469 5466
rect 16521 5414 16533 5466
rect 16585 5414 16597 5466
rect 16649 5414 16661 5466
rect 16713 5414 26709 5466
rect 26761 5414 26773 5466
rect 26825 5414 26837 5466
rect 26889 5414 26901 5466
rect 26953 5414 26965 5466
rect 27017 5414 32016 5466
rect 1104 5392 32016 5414
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 3016 5324 3065 5352
rect 3016 5312 3022 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 5166 5352 5172 5364
rect 5127 5324 5172 5352
rect 3053 5315 3111 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 11974 5352 11980 5364
rect 9640 5324 11980 5352
rect 9640 5312 9646 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 17221 5355 17279 5361
rect 17221 5321 17233 5355
rect 17267 5352 17279 5355
rect 17678 5352 17684 5364
rect 17267 5324 17684 5352
rect 17267 5321 17279 5324
rect 17221 5315 17279 5321
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 18230 5312 18236 5364
rect 18288 5312 18294 5364
rect 18690 5352 18696 5364
rect 18651 5324 18696 5352
rect 18690 5312 18696 5324
rect 18748 5312 18754 5364
rect 19245 5355 19303 5361
rect 19245 5321 19257 5355
rect 19291 5352 19303 5355
rect 19291 5324 22600 5352
rect 19291 5321 19303 5324
rect 19245 5315 19303 5321
rect 9125 5287 9183 5293
rect 9125 5253 9137 5287
rect 9171 5284 9183 5287
rect 10778 5284 10784 5296
rect 9171 5256 10784 5284
rect 9171 5253 9183 5256
rect 9125 5247 9183 5253
rect 10778 5244 10784 5256
rect 10836 5244 10842 5296
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 11238 5284 11244 5296
rect 11112 5256 11244 5284
rect 11112 5244 11118 5256
rect 11238 5244 11244 5256
rect 11296 5244 11302 5296
rect 12710 5284 12716 5296
rect 12268 5256 12716 5284
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 7742 5216 7748 5228
rect 7515 5188 7748 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9646 5188 10241 5216
rect 0 5148 800 5162
rect 1670 5148 1676 5160
rect 0 5120 888 5148
rect 1631 5120 1676 5148
rect 0 5106 800 5120
rect 860 5012 888 5120
rect 1670 5108 1676 5120
rect 1728 5148 1734 5160
rect 3786 5148 3792 5160
rect 1728 5120 3792 5148
rect 1728 5108 1734 5120
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4062 5157 4068 5160
rect 4056 5148 4068 5157
rect 4023 5120 4068 5148
rect 4056 5111 4068 5120
rect 4062 5108 4068 5111
rect 4120 5108 4126 5160
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 6822 5148 6828 5160
rect 5776 5120 6828 5148
rect 5776 5108 5782 5120
rect 1762 5040 1768 5092
rect 1820 5080 1826 5092
rect 1918 5083 1976 5089
rect 1918 5080 1930 5083
rect 1820 5052 1930 5080
rect 1820 5040 1826 5052
rect 1918 5049 1930 5052
rect 1964 5049 1976 5083
rect 1918 5043 1976 5049
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 5626 5080 5632 5092
rect 4212 5052 5632 5080
rect 4212 5040 4218 5052
rect 5626 5040 5632 5052
rect 5684 5080 5690 5092
rect 5994 5080 6000 5092
rect 5684 5052 6000 5080
rect 5684 5040 5690 5052
rect 5994 5040 6000 5052
rect 6052 5040 6058 5092
rect 768 4984 888 5012
rect 768 4740 796 4984
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2682 5012 2688 5024
rect 2372 4984 2688 5012
rect 2372 4972 2378 4984
rect 2682 4972 2688 4984
rect 2740 5012 2746 5024
rect 5350 5012 5356 5024
rect 2740 4984 5356 5012
rect 2740 4972 2746 4984
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 6104 5021 6132 5120
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 6880 5120 7941 5148
rect 6880 5108 6886 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 9214 5148 9220 5160
rect 9175 5120 9220 5148
rect 7929 5111 7987 5117
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9646 5148 9674 5188
rect 10229 5185 10241 5188
rect 10275 5216 10287 5219
rect 10594 5216 10600 5228
rect 10275 5188 10600 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 10594 5176 10600 5188
rect 10652 5176 10658 5228
rect 10962 5216 10968 5228
rect 10875 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5216 11026 5228
rect 12268 5216 12296 5256
rect 12710 5244 12716 5256
rect 12768 5244 12774 5296
rect 14366 5284 14372 5296
rect 13004 5256 14372 5284
rect 11020 5188 12296 5216
rect 11020 5176 11026 5188
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 13004 5225 13032 5256
rect 14366 5244 14372 5256
rect 14424 5244 14430 5296
rect 17126 5284 17132 5296
rect 16776 5256 17132 5284
rect 16776 5225 16804 5256
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12400 5188 12909 5216
rect 12400 5176 12406 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5216 16911 5219
rect 17218 5216 17224 5228
rect 16899 5188 17224 5216
rect 16899 5185 16911 5188
rect 16853 5179 16911 5185
rect 9456 5120 9674 5148
rect 10505 5151 10563 5157
rect 9456 5108 9462 5120
rect 10505 5117 10517 5151
rect 10551 5117 10563 5151
rect 10505 5111 10563 5117
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7202 5083 7260 5089
rect 7202 5080 7214 5083
rect 7156 5052 7214 5080
rect 7156 5040 7162 5052
rect 7202 5049 7214 5052
rect 7248 5049 7260 5083
rect 10520 5080 10548 5111
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 10744 5120 11253 5148
rect 10744 5108 10750 5120
rect 11241 5117 11253 5120
rect 11287 5117 11299 5151
rect 12618 5148 12624 5160
rect 12579 5120 12624 5148
rect 11241 5111 11299 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12802 5148 12808 5160
rect 12763 5120 12808 5148
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 10962 5080 10968 5092
rect 10520 5052 10968 5080
rect 7202 5043 7260 5049
rect 10962 5040 10968 5052
rect 11020 5080 11026 5092
rect 11606 5080 11612 5092
rect 11020 5052 11612 5080
rect 11020 5040 11026 5052
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 12250 5040 12256 5092
rect 12308 5080 12314 5092
rect 12636 5080 12664 5108
rect 12308 5052 12664 5080
rect 12308 5040 12314 5052
rect 6089 5015 6147 5021
rect 6089 4981 6101 5015
rect 6135 4981 6147 5015
rect 6089 4975 6147 4981
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 6972 4984 8125 5012
rect 6972 4972 6978 4984
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 13004 5012 13032 5179
rect 17218 5176 17224 5188
rect 17276 5216 17282 5228
rect 18046 5216 18052 5228
rect 17276 5188 18052 5216
rect 17276 5176 17282 5188
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 18248 5225 18276 5312
rect 18598 5244 18604 5296
rect 18656 5284 18662 5296
rect 20714 5284 20720 5296
rect 18656 5256 20720 5284
rect 18656 5244 18662 5256
rect 20714 5244 20720 5256
rect 20772 5244 20778 5296
rect 22572 5284 22600 5324
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25593 5355 25651 5361
rect 25593 5352 25605 5355
rect 25004 5324 25605 5352
rect 25004 5312 25010 5324
rect 25593 5321 25605 5324
rect 25639 5321 25651 5355
rect 25593 5315 25651 5321
rect 27062 5312 27068 5364
rect 27120 5352 27126 5364
rect 27798 5352 27804 5364
rect 27120 5324 27804 5352
rect 27120 5312 27126 5324
rect 27798 5312 27804 5324
rect 27856 5352 27862 5364
rect 28169 5355 28227 5361
rect 28169 5352 28181 5355
rect 27856 5324 28181 5352
rect 27856 5312 27862 5324
rect 28169 5321 28181 5324
rect 28215 5321 28227 5355
rect 28718 5352 28724 5364
rect 28679 5324 28724 5352
rect 28169 5315 28227 5321
rect 28718 5312 28724 5324
rect 28776 5312 28782 5364
rect 29641 5355 29699 5361
rect 29641 5321 29653 5355
rect 29687 5352 29699 5355
rect 30006 5352 30012 5364
rect 29687 5324 30012 5352
rect 29687 5321 29699 5324
rect 29641 5315 29699 5321
rect 30006 5312 30012 5324
rect 30064 5312 30070 5364
rect 30650 5352 30656 5364
rect 30563 5324 30656 5352
rect 30650 5312 30656 5324
rect 30708 5352 30714 5364
rect 31110 5352 31116 5364
rect 30708 5324 31116 5352
rect 30708 5312 30714 5324
rect 31110 5312 31116 5324
rect 31168 5312 31174 5364
rect 24578 5284 24584 5296
rect 22572 5256 24584 5284
rect 18227 5219 18285 5225
rect 18227 5185 18239 5219
rect 18273 5185 18285 5219
rect 20990 5216 20996 5228
rect 18227 5179 18285 5185
rect 18524 5188 20996 5216
rect 13170 5148 13176 5160
rect 13131 5120 13176 5148
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14332 5120 14381 5148
rect 14332 5108 14338 5120
rect 14369 5117 14381 5120
rect 14415 5148 14427 5151
rect 15746 5148 15752 5160
rect 14415 5120 15752 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 16485 5151 16543 5157
rect 16485 5117 16497 5151
rect 16531 5117 16543 5151
rect 16485 5111 16543 5117
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 17037 5151 17095 5157
rect 17037 5117 17049 5151
rect 17083 5148 17095 5151
rect 17402 5148 17408 5160
rect 17083 5120 17408 5148
rect 17083 5117 17095 5120
rect 17037 5111 17095 5117
rect 14636 5083 14694 5089
rect 14636 5049 14648 5083
rect 14682 5080 14694 5083
rect 15010 5080 15016 5092
rect 14682 5052 15016 5080
rect 14682 5049 14694 5052
rect 14636 5043 14694 5049
rect 15010 5040 15016 5052
rect 15068 5040 15074 5092
rect 13078 5012 13084 5024
rect 11940 4984 13084 5012
rect 11940 4972 11946 4984
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 14366 5012 14372 5024
rect 13403 4984 14372 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 15654 4972 15660 5024
rect 15712 5012 15718 5024
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15712 4984 15761 5012
rect 15712 4972 15718 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 16500 5012 16528 5111
rect 16684 5080 16712 5111
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 17954 5148 17960 5160
rect 17915 5120 17960 5148
rect 17954 5108 17960 5120
rect 18012 5108 18018 5160
rect 18138 5148 18144 5160
rect 18099 5120 18144 5148
rect 18138 5108 18144 5120
rect 18196 5108 18202 5160
rect 18524 5157 18552 5188
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5216 22155 5219
rect 22370 5216 22376 5228
rect 22143 5188 22376 5216
rect 22143 5185 22155 5188
rect 22097 5179 22155 5185
rect 22370 5176 22376 5188
rect 22428 5176 22434 5228
rect 22572 5225 22600 5256
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 26050 5284 26056 5296
rect 25976 5256 26056 5284
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5185 22615 5219
rect 22830 5216 22836 5228
rect 22791 5188 22836 5216
rect 22557 5179 22615 5185
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 22922 5176 22928 5228
rect 22980 5216 22986 5228
rect 24486 5216 24492 5228
rect 22980 5188 24492 5216
rect 22980 5176 22986 5188
rect 24486 5176 24492 5188
rect 24544 5216 24550 5228
rect 25976 5225 26004 5256
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 27430 5244 27436 5296
rect 27488 5284 27494 5296
rect 30282 5284 30288 5296
rect 27488 5256 30288 5284
rect 27488 5244 27494 5256
rect 30282 5244 30288 5256
rect 30340 5244 30346 5296
rect 24765 5219 24823 5225
rect 24765 5216 24777 5219
rect 24544 5188 24777 5216
rect 24544 5176 24550 5188
rect 24765 5185 24777 5188
rect 24811 5185 24823 5219
rect 24765 5179 24823 5185
rect 25961 5219 26019 5225
rect 25961 5185 25973 5219
rect 26007 5185 26019 5219
rect 25961 5179 26019 5185
rect 26878 5176 26884 5228
rect 26936 5216 26942 5228
rect 27258 5219 27316 5225
rect 27258 5216 27270 5219
rect 26936 5188 27270 5216
rect 26936 5176 26942 5188
rect 27258 5185 27270 5188
rect 27304 5185 27316 5219
rect 27258 5179 27316 5185
rect 18371 5151 18429 5157
rect 18371 5117 18383 5151
rect 18417 5117 18429 5151
rect 18371 5111 18429 5117
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 16684 5052 16896 5080
rect 16868 5024 16896 5052
rect 18046 5040 18052 5092
rect 18104 5080 18110 5092
rect 18386 5080 18414 5111
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 19245 5151 19303 5157
rect 19245 5148 19257 5151
rect 18656 5120 19257 5148
rect 18656 5108 18662 5120
rect 19245 5117 19257 5120
rect 19291 5148 19303 5151
rect 19337 5151 19395 5157
rect 19337 5148 19349 5151
rect 19291 5120 19349 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 19337 5117 19349 5120
rect 19383 5117 19395 5151
rect 19337 5111 19395 5117
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5148 19671 5151
rect 19794 5148 19800 5160
rect 19659 5120 19800 5148
rect 19659 5117 19671 5120
rect 19613 5111 19671 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 23474 5108 23480 5160
rect 23532 5148 23538 5160
rect 24581 5151 24639 5157
rect 24581 5148 24593 5151
rect 23532 5120 24593 5148
rect 23532 5108 23538 5120
rect 24581 5117 24593 5120
rect 24627 5117 24639 5151
rect 24854 5148 24860 5160
rect 24815 5120 24860 5148
rect 24581 5111 24639 5117
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 24949 5151 25007 5157
rect 24949 5117 24961 5151
rect 24995 5117 25007 5151
rect 25130 5148 25136 5160
rect 25091 5120 25136 5148
rect 24949 5111 25007 5117
rect 21818 5080 21824 5092
rect 21876 5089 21882 5092
rect 18104 5052 18414 5080
rect 21788 5052 21824 5080
rect 18104 5040 18110 5052
rect 21818 5040 21824 5052
rect 21876 5043 21888 5089
rect 21876 5040 21882 5043
rect 23658 5040 23664 5092
rect 23716 5080 23722 5092
rect 24964 5080 24992 5111
rect 25130 5108 25136 5120
rect 25188 5108 25194 5160
rect 25777 5151 25835 5157
rect 25777 5117 25789 5151
rect 25823 5117 25835 5151
rect 26050 5148 26056 5160
rect 26011 5120 26056 5148
rect 25777 5111 25835 5117
rect 23716 5052 24992 5080
rect 23716 5040 23722 5052
rect 16758 5012 16764 5024
rect 16500 4984 16764 5012
rect 15749 4975 15807 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 16850 4972 16856 5024
rect 16908 4972 16914 5024
rect 18874 4972 18880 5024
rect 18932 5012 18938 5024
rect 20714 5012 20720 5024
rect 18932 4984 20720 5012
rect 18932 4972 18938 4984
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 24302 4972 24308 5024
rect 24360 5012 24366 5024
rect 24397 5015 24455 5021
rect 24397 5012 24409 5015
rect 24360 4984 24409 5012
rect 24360 4972 24366 4984
rect 24397 4981 24409 4984
rect 24443 4981 24455 5015
rect 25792 5012 25820 5111
rect 26050 5108 26056 5120
rect 26108 5108 26114 5160
rect 26145 5151 26203 5157
rect 26145 5117 26157 5151
rect 26191 5148 26203 5151
rect 26234 5148 26240 5160
rect 26191 5120 26240 5148
rect 26191 5117 26203 5120
rect 26145 5111 26203 5117
rect 26234 5108 26240 5120
rect 26292 5108 26298 5160
rect 26329 5151 26387 5157
rect 26329 5117 26341 5151
rect 26375 5117 26387 5151
rect 26329 5111 26387 5117
rect 26973 5151 27031 5157
rect 26973 5117 26985 5151
rect 27019 5148 27031 5151
rect 27062 5148 27068 5160
rect 27019 5120 27068 5148
rect 27019 5117 27031 5120
rect 26973 5111 27031 5117
rect 26344 5080 26372 5111
rect 27062 5108 27068 5120
rect 27120 5108 27126 5160
rect 27157 5151 27215 5157
rect 27157 5117 27169 5151
rect 27203 5117 27215 5151
rect 27157 5111 27215 5117
rect 27341 5151 27399 5157
rect 27341 5117 27353 5151
rect 27387 5150 27399 5151
rect 27430 5150 27436 5160
rect 27387 5122 27436 5150
rect 27387 5117 27399 5122
rect 27341 5111 27399 5117
rect 27172 5080 27200 5111
rect 27430 5108 27436 5122
rect 27488 5108 27494 5160
rect 27525 5151 27583 5157
rect 27525 5117 27537 5151
rect 27571 5148 27583 5151
rect 27614 5148 27620 5160
rect 27571 5120 27620 5148
rect 27571 5117 27583 5120
rect 27525 5111 27583 5117
rect 27614 5108 27620 5120
rect 27672 5108 27678 5160
rect 31113 5151 31171 5157
rect 31113 5117 31125 5151
rect 31159 5148 31171 5151
rect 31294 5148 31300 5160
rect 31159 5120 31300 5148
rect 31159 5117 31171 5120
rect 31113 5111 31171 5117
rect 31294 5108 31300 5120
rect 31352 5108 31358 5160
rect 32320 5148 33120 5162
rect 31726 5120 33120 5148
rect 27246 5080 27252 5092
rect 26344 5052 27108 5080
rect 27172 5052 27252 5080
rect 26326 5012 26332 5024
rect 25792 4984 26332 5012
rect 24397 4975 24455 4981
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 27080 5012 27108 5052
rect 27246 5040 27252 5052
rect 27304 5040 27310 5092
rect 27430 5012 27436 5024
rect 27080 4984 27436 5012
rect 27430 4972 27436 4984
rect 27488 4972 27494 5024
rect 27706 5012 27712 5024
rect 27667 4984 27712 5012
rect 27706 4972 27712 4984
rect 27764 4972 27770 5024
rect 31297 5015 31355 5021
rect 31297 4981 31309 5015
rect 31343 5012 31355 5015
rect 31726 5012 31754 5120
rect 32320 5106 33120 5120
rect 31343 4984 31754 5012
rect 31343 4981 31355 4984
rect 31297 4975 31355 4981
rect 1104 4922 32016 4944
rect 1104 4870 11253 4922
rect 11305 4870 11317 4922
rect 11369 4870 11381 4922
rect 11433 4870 11445 4922
rect 11497 4870 11509 4922
rect 11561 4870 21557 4922
rect 21609 4870 21621 4922
rect 21673 4870 21685 4922
rect 21737 4870 21749 4922
rect 21801 4870 21813 4922
rect 21865 4870 32016 4922
rect 1104 4848 32016 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2130 4808 2136 4820
rect 1995 4780 2136 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2593 4811 2651 4817
rect 2593 4777 2605 4811
rect 2639 4808 2651 4811
rect 2682 4808 2688 4820
rect 2639 4780 2688 4808
rect 2639 4777 2651 4780
rect 2593 4771 2651 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 3050 4808 3056 4820
rect 3011 4780 3056 4808
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 3694 4808 3700 4820
rect 3655 4780 3700 4808
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 7098 4808 7104 4820
rect 4672 4780 6684 4808
rect 7059 4780 7104 4808
rect 4672 4768 4678 4780
rect 1857 4743 1915 4749
rect 1857 4740 1869 4743
rect 768 4712 1869 4740
rect 1857 4709 1869 4712
rect 1903 4740 1915 4743
rect 3234 4740 3240 4752
rect 1903 4712 3240 4740
rect 1903 4709 1915 4712
rect 1857 4703 1915 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 4632 4712 6592 4740
rect 3142 4632 3148 4684
rect 3200 4672 3206 4684
rect 3878 4672 3884 4684
rect 3200 4644 3884 4672
rect 3200 4632 3206 4644
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 4632 4681 4660 4712
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 4488 4644 4629 4672
rect 4488 4632 4494 4644
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4764 4644 4813 4672
rect 4764 4632 4770 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 5000 4604 5028 4635
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 6564 4681 6592 4712
rect 5169 4675 5227 4681
rect 5169 4672 5181 4675
rect 5132 4644 5181 4672
rect 5132 4632 5138 4644
rect 5169 4641 5181 4644
rect 5215 4672 5227 4675
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 5215 4644 6377 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 6365 4641 6377 4644
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4641 6607 4675
rect 6656 4672 6684 4780
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9122 4808 9128 4820
rect 9079 4780 9128 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 13998 4808 14004 4820
rect 12299 4780 14004 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 15562 4808 15568 4820
rect 14415 4780 15568 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 19242 4808 19248 4820
rect 18708 4780 19248 4808
rect 12526 4740 12532 4752
rect 11716 4712 12532 4740
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6656 4644 6745 4672
rect 6549 4635 6607 4641
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6733 4635 6791 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4672 7711 4675
rect 7742 4672 7748 4684
rect 7699 4644 7748 4672
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 7920 4675 7978 4681
rect 7920 4641 7932 4675
rect 7966 4672 7978 4675
rect 9122 4672 9128 4684
rect 7966 4644 9128 4672
rect 7966 4641 7978 4644
rect 7920 4635 7978 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 11054 4672 11060 4684
rect 10643 4644 11060 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11716 4681 11744 4712
rect 12526 4700 12532 4712
rect 12584 4700 12590 4752
rect 13170 4700 13176 4752
rect 13228 4740 13234 4752
rect 15194 4740 15200 4752
rect 13228 4712 15200 4740
rect 13228 4700 13234 4712
rect 11517 4675 11575 4681
rect 11517 4641 11529 4675
rect 11563 4672 11575 4675
rect 11701 4675 11759 4681
rect 11563 4644 11652 4672
rect 11563 4641 11575 4644
rect 11517 4635 11575 4641
rect 5258 4604 5264 4616
rect 5000 4576 5264 4604
rect 4893 4567 4951 4573
rect 4908 4536 4936 4567
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5684 4576 5733 4604
rect 5684 4564 5690 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 6454 4536 6460 4548
rect 4908 4508 6460 4536
rect 6454 4496 6460 4508
rect 6512 4536 6518 4548
rect 6656 4536 6684 4567
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 10284 4576 10333 4604
rect 10284 4564 10290 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 6512 4508 6684 4536
rect 11624 4536 11652 4644
rect 11701 4641 11713 4675
rect 11747 4641 11759 4675
rect 11882 4672 11888 4684
rect 11843 4644 11888 4672
rect 11701 4635 11759 4641
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12069 4675 12127 4681
rect 12069 4641 12081 4675
rect 12115 4672 12127 4675
rect 12802 4672 12808 4684
rect 12115 4644 12808 4672
rect 12115 4641 12127 4644
rect 12069 4635 12127 4641
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4641 12955 4675
rect 13078 4672 13084 4684
rect 13039 4644 13084 4672
rect 12897 4635 12955 4641
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 11839 4576 12388 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12360 4548 12388 4576
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12912 4604 12940 4635
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13280 4681 13308 4712
rect 15194 4700 15200 4712
rect 15252 4700 15258 4752
rect 18141 4743 18199 4749
rect 18141 4709 18153 4743
rect 18187 4740 18199 4743
rect 18598 4740 18604 4752
rect 18187 4712 18604 4740
rect 18187 4709 18199 4712
rect 18141 4703 18199 4709
rect 18598 4700 18604 4712
rect 18656 4700 18662 4752
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 13446 4672 13452 4684
rect 13407 4644 13452 4672
rect 13265 4635 13323 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 15470 4672 15476 4684
rect 15528 4681 15534 4684
rect 15440 4644 15476 4672
rect 15470 4632 15476 4644
rect 15528 4635 15540 4681
rect 15746 4672 15752 4684
rect 15707 4644 15752 4672
rect 15528 4632 15534 4635
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 17494 4672 17500 4684
rect 17455 4644 17500 4672
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 18708 4681 18736 4780
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 19429 4811 19487 4817
rect 19429 4777 19441 4811
rect 19475 4808 19487 4811
rect 19610 4808 19616 4820
rect 19475 4780 19616 4808
rect 19475 4777 19487 4780
rect 19429 4771 19487 4777
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 21821 4811 21879 4817
rect 21821 4777 21833 4811
rect 21867 4808 21879 4811
rect 21910 4808 21916 4820
rect 21867 4780 21916 4808
rect 21867 4777 21879 4780
rect 21821 4771 21879 4777
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 23017 4811 23075 4817
rect 23017 4777 23029 4811
rect 23063 4808 23075 4811
rect 23474 4808 23480 4820
rect 23063 4780 23480 4808
rect 23063 4777 23075 4780
rect 23017 4771 23075 4777
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 26510 4768 26516 4820
rect 26568 4808 26574 4820
rect 27065 4811 27123 4817
rect 27065 4808 27077 4811
rect 26568 4780 27077 4808
rect 26568 4768 26574 4780
rect 27065 4777 27077 4780
rect 27111 4777 27123 4811
rect 27614 4808 27620 4820
rect 27065 4771 27123 4777
rect 27172 4780 27620 4808
rect 19058 4700 19064 4752
rect 19116 4740 19122 4752
rect 20438 4740 20444 4752
rect 19116 4712 19288 4740
rect 19116 4700 19122 4712
rect 18693 4675 18751 4681
rect 18693 4641 18705 4675
rect 18739 4641 18751 4675
rect 18874 4672 18880 4684
rect 18835 4644 18880 4672
rect 18693 4635 18751 4641
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 19260 4681 19288 4712
rect 19904 4712 20444 4740
rect 19904 4681 19932 4712
rect 20438 4700 20444 4712
rect 20496 4700 20502 4752
rect 22186 4700 22192 4752
rect 22244 4740 22250 4752
rect 22244 4712 22416 4740
rect 22244 4700 22250 4712
rect 20162 4681 20168 4684
rect 18969 4675 19027 4681
rect 18969 4641 18981 4675
rect 19015 4672 19027 4675
rect 19245 4675 19303 4681
rect 19015 4644 19196 4672
rect 19015 4641 19027 4644
rect 18969 4635 19027 4641
rect 12492 4576 12940 4604
rect 13173 4607 13231 4613
rect 12492 4564 12498 4576
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 12250 4536 12256 4548
rect 11624 4508 12256 4536
rect 6512 4496 6518 4508
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 13188 4536 13216 4567
rect 16298 4564 16304 4616
rect 16356 4604 16362 4616
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 16356 4576 17233 4604
rect 16356 4564 16362 4576
rect 17221 4573 17233 4576
rect 17267 4604 17279 4607
rect 17402 4604 17408 4616
rect 17267 4576 17408 4604
rect 17267 4573 17279 4576
rect 17221 4567 17279 4573
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 19058 4604 19064 4616
rect 19019 4576 19064 4604
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19168 4604 19196 4644
rect 19245 4641 19257 4675
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 19889 4675 19947 4681
rect 19889 4641 19901 4675
rect 19935 4641 19947 4675
rect 20156 4672 20168 4681
rect 20123 4644 20168 4672
rect 19889 4635 19947 4641
rect 20156 4635 20168 4644
rect 20162 4632 20168 4635
rect 20220 4632 20226 4684
rect 20714 4632 20720 4684
rect 20772 4672 20778 4684
rect 22388 4681 22416 4712
rect 23934 4700 23940 4752
rect 23992 4740 23998 4752
rect 23992 4712 24440 4740
rect 23992 4700 23998 4712
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 20772 4644 22017 4672
rect 20772 4632 20778 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22005 4635 22063 4641
rect 22373 4675 22431 4681
rect 22373 4641 22385 4675
rect 22419 4641 22431 4675
rect 22554 4672 22560 4684
rect 22515 4644 22560 4672
rect 22373 4635 22431 4641
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 24141 4675 24199 4681
rect 24141 4641 24153 4675
rect 24187 4672 24199 4675
rect 24302 4672 24308 4684
rect 24187 4644 24308 4672
rect 24187 4641 24199 4644
rect 24141 4635 24199 4641
rect 24302 4632 24308 4644
rect 24360 4632 24366 4684
rect 24412 4681 24440 4712
rect 26050 4700 26056 4752
rect 26108 4740 26114 4752
rect 26878 4740 26884 4752
rect 26108 4712 26884 4740
rect 26108 4700 26114 4712
rect 26878 4700 26884 4712
rect 26936 4700 26942 4752
rect 24397 4675 24455 4681
rect 24397 4641 24409 4675
rect 24443 4672 24455 4675
rect 24762 4672 24768 4684
rect 24443 4644 24768 4672
rect 24443 4641 24455 4644
rect 24397 4635 24455 4641
rect 24762 4632 24768 4644
rect 24820 4632 24826 4684
rect 24857 4675 24915 4681
rect 24857 4641 24869 4675
rect 24903 4672 24915 4675
rect 25038 4672 25044 4684
rect 24903 4644 25044 4672
rect 24903 4641 24915 4644
rect 24857 4635 24915 4641
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 26142 4672 26148 4684
rect 26103 4644 26148 4672
rect 26142 4632 26148 4644
rect 26200 4632 26206 4684
rect 27172 4681 27200 4780
rect 27614 4768 27620 4780
rect 27672 4768 27678 4820
rect 29917 4811 29975 4817
rect 29917 4777 29929 4811
rect 29963 4808 29975 4811
rect 30006 4808 30012 4820
rect 29963 4780 30012 4808
rect 29963 4777 29975 4780
rect 29917 4771 29975 4777
rect 30006 4768 30012 4780
rect 30064 4808 30070 4820
rect 30558 4808 30564 4820
rect 30064 4780 30564 4808
rect 30064 4768 30070 4780
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 31018 4808 31024 4820
rect 30979 4780 31024 4808
rect 31018 4768 31024 4780
rect 31076 4768 31082 4820
rect 27706 4700 27712 4752
rect 27764 4740 27770 4752
rect 28730 4743 28788 4749
rect 28730 4740 28742 4743
rect 27764 4712 28742 4740
rect 27764 4700 27770 4712
rect 28730 4709 28742 4712
rect 28776 4709 28788 4743
rect 30466 4740 30472 4752
rect 30379 4712 30472 4740
rect 28730 4703 28788 4709
rect 30466 4700 30472 4712
rect 30524 4740 30530 4752
rect 31202 4740 31208 4752
rect 30524 4712 31208 4740
rect 30524 4700 30530 4712
rect 31202 4700 31208 4712
rect 31260 4700 31266 4752
rect 27157 4675 27215 4681
rect 27157 4641 27169 4675
rect 27203 4641 27215 4675
rect 28994 4672 29000 4684
rect 28955 4644 29000 4672
rect 27157 4635 27215 4641
rect 19794 4604 19800 4616
rect 19168 4576 19800 4604
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 22186 4604 22192 4616
rect 22066 4576 22192 4604
rect 17954 4536 17960 4548
rect 12400 4508 13216 4536
rect 17915 4508 17960 4536
rect 12400 4496 12406 4508
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 22066 4536 22094 4576
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4604 22339 4607
rect 22830 4604 22836 4616
rect 22327 4576 22836 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 25130 4604 25136 4616
rect 25091 4576 25136 4604
rect 25130 4564 25136 4576
rect 25188 4564 25194 4616
rect 25958 4564 25964 4616
rect 26016 4604 26022 4616
rect 27172 4604 27200 4635
rect 28994 4632 29000 4644
rect 29052 4632 29058 4684
rect 26016 4576 27200 4604
rect 26016 4564 26022 4576
rect 20824 4508 22094 4536
rect 26237 4539 26295 4545
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4468 4491 4471
rect 5534 4468 5540 4480
rect 4479 4440 5540 4468
rect 4479 4437 4491 4440
rect 4433 4431 4491 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 12710 4468 12716 4480
rect 12671 4440 12716 4468
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 19886 4428 19892 4480
rect 19944 4468 19950 4480
rect 20824 4468 20852 4508
rect 26237 4505 26249 4539
rect 26283 4536 26295 4539
rect 27982 4536 27988 4548
rect 26283 4508 27988 4536
rect 26283 4505 26295 4508
rect 26237 4499 26295 4505
rect 27982 4496 27988 4508
rect 28040 4496 28046 4548
rect 19944 4440 20852 4468
rect 19944 4428 19950 4440
rect 21082 4428 21088 4480
rect 21140 4468 21146 4480
rect 21269 4471 21327 4477
rect 21269 4468 21281 4471
rect 21140 4440 21281 4468
rect 21140 4428 21146 4440
rect 21269 4437 21281 4440
rect 21315 4437 21327 4471
rect 21269 4431 21327 4437
rect 26418 4428 26424 4480
rect 26476 4468 26482 4480
rect 28350 4468 28356 4480
rect 26476 4440 28356 4468
rect 26476 4428 26482 4440
rect 28350 4428 28356 4440
rect 28408 4428 28414 4480
rect 1104 4378 32016 4400
rect 1104 4326 6102 4378
rect 6154 4326 6166 4378
rect 6218 4326 6230 4378
rect 6282 4326 6294 4378
rect 6346 4326 6358 4378
rect 6410 4326 16405 4378
rect 16457 4326 16469 4378
rect 16521 4326 16533 4378
rect 16585 4326 16597 4378
rect 16649 4326 16661 4378
rect 16713 4326 26709 4378
rect 26761 4326 26773 4378
rect 26825 4326 26837 4378
rect 26889 4326 26901 4378
rect 26953 4326 26965 4378
rect 27017 4326 32016 4378
rect 1104 4304 32016 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4264 1734 4276
rect 2866 4264 2872 4276
rect 1728 4236 2872 4264
rect 1728 4224 1734 4236
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 4430 4264 4436 4276
rect 4391 4236 4436 4264
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7009 4267 7067 4273
rect 7009 4264 7021 4267
rect 6972 4236 7021 4264
rect 6972 4224 6978 4236
rect 7009 4233 7021 4236
rect 7055 4233 7067 4267
rect 7009 4227 7067 4233
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 12400 4236 12572 4264
rect 12400 4224 12406 4236
rect 4338 4196 4344 4208
rect 3896 4168 4344 4196
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 3789 4131 3847 4137
rect 3789 4128 3801 4131
rect 1912 4100 3801 4128
rect 1912 4088 1918 4100
rect 3789 4097 3801 4100
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 3896 4060 3924 4168
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 7742 4156 7748 4208
rect 7800 4156 7806 4208
rect 10686 4196 10692 4208
rect 10336 4168 10692 4196
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 7760 4128 7788 4156
rect 8294 4128 8300 4140
rect 5859 4100 7788 4128
rect 8255 4100 8300 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9456 4100 9505 4128
rect 9456 4088 9462 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4128 9643 4131
rect 10226 4128 10232 4140
rect 9631 4100 10232 4128
rect 9631 4097 9643 4100
rect 9585 4091 9643 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 2363 4032 3924 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 5534 4020 5540 4072
rect 5592 4069 5598 4072
rect 5592 4060 5604 4069
rect 7745 4063 7803 4069
rect 5592 4032 5637 4060
rect 5592 4023 5604 4032
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 7926 4060 7932 4072
rect 7791 4032 7932 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 5592 4020 5598 4023
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 8570 4060 8576 4072
rect 8435 4032 8576 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 9309 4063 9367 4069
rect 9309 4060 9321 4063
rect 9272 4032 9321 4060
rect 9272 4020 9278 4032
rect 9309 4029 9321 4032
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 10042 4060 10048 4072
rect 9907 4032 10048 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 4890 3992 4896 4004
rect 2915 3964 4896 3992
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 7944 3992 7972 4020
rect 9692 3992 9720 4023
rect 10042 4020 10048 4032
rect 10100 4060 10106 4072
rect 10336 4060 10364 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 12544 4137 12572 4236
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 12860 4236 13461 4264
rect 12860 4224 12866 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 13449 4227 13507 4233
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 14185 4267 14243 4273
rect 14185 4264 14197 4267
rect 13872 4236 14197 4264
rect 13872 4224 13878 4236
rect 14185 4233 14197 4236
rect 14231 4233 14243 4267
rect 15470 4264 15476 4276
rect 15431 4236 15476 4264
rect 14185 4227 14243 4233
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 17954 4264 17960 4276
rect 15948 4236 17960 4264
rect 12618 4156 12624 4208
rect 12676 4196 12682 4208
rect 14090 4196 14096 4208
rect 12676 4168 14096 4196
rect 12676 4156 12682 4168
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 12529 4131 12587 4137
rect 10520 4100 12388 4128
rect 10520 4069 10548 4100
rect 10100 4032 10364 4060
rect 10505 4063 10563 4069
rect 10100 4020 10106 4032
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10962 4060 10968 4072
rect 10923 4032 10968 4060
rect 10505 4023 10563 4029
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 12250 4060 12256 4072
rect 12211 4032 12256 4060
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 12360 4060 12388 4100
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 13630 4088 13636 4140
rect 13688 4128 13694 4140
rect 13688 4100 14412 4128
rect 13688 4088 13694 4100
rect 12434 4060 12440 4072
rect 12360 4032 12440 4060
rect 12434 4020 12440 4032
rect 12492 4060 12498 4072
rect 12621 4063 12679 4069
rect 12492 4032 12537 4060
rect 12492 4020 12498 4032
rect 12621 4029 12633 4063
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13170 4060 13176 4072
rect 12851 4032 13176 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 9950 3992 9956 4004
rect 7944 3964 9956 3992
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10318 3992 10324 4004
rect 10060 3964 10324 3992
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3924 6607 3927
rect 7282 3924 7288 3936
rect 6595 3896 7288 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 7653 3927 7711 3933
rect 7653 3893 7665 3927
rect 7699 3924 7711 3927
rect 10060 3924 10088 3964
rect 10318 3952 10324 3964
rect 10376 3952 10382 4004
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 12526 3992 12532 4004
rect 10459 3964 12532 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 7699 3896 10088 3924
rect 7699 3893 7711 3896
rect 7653 3887 7711 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10594 3924 10600 3936
rect 10192 3896 10600 3924
rect 10192 3884 10198 3896
rect 10594 3884 10600 3896
rect 10652 3924 10658 3936
rect 11195 3927 11253 3933
rect 11195 3924 11207 3927
rect 10652 3896 11207 3924
rect 10652 3884 10658 3896
rect 11195 3893 11207 3896
rect 11241 3924 11253 3927
rect 12636 3924 12664 4023
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 14090 4060 14096 4072
rect 14051 4032 14096 4060
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 14384 4069 14412 4100
rect 14550 4088 14556 4140
rect 14608 4128 14614 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14608 4100 14657 4128
rect 14608 4088 14614 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 15378 4088 15384 4140
rect 15436 4128 15442 4140
rect 15948 4137 15976 4236
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 18138 4224 18144 4276
rect 18196 4264 18202 4276
rect 20625 4267 20683 4273
rect 20625 4264 20637 4267
rect 18196 4236 20637 4264
rect 18196 4224 18202 4236
rect 20625 4233 20637 4236
rect 20671 4233 20683 4267
rect 20625 4227 20683 4233
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 22465 4267 22523 4273
rect 22465 4264 22477 4267
rect 22428 4236 22477 4264
rect 22428 4224 22434 4236
rect 22465 4233 22477 4236
rect 22511 4233 22523 4267
rect 22465 4227 22523 4233
rect 27430 4224 27436 4276
rect 27488 4264 27494 4276
rect 28077 4267 28135 4273
rect 28077 4264 28089 4267
rect 27488 4236 28089 4264
rect 27488 4224 27494 4236
rect 28077 4233 28089 4236
rect 28123 4233 28135 4267
rect 28077 4227 28135 4233
rect 17218 4156 17224 4208
rect 17276 4196 17282 4208
rect 18230 4196 18236 4208
rect 17276 4168 18236 4196
rect 17276 4156 17282 4168
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 15436 4100 15853 4128
rect 15436 4088 15442 4100
rect 15841 4097 15853 4100
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 16758 4128 16764 4140
rect 16715 4100 16764 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17586 4128 17592 4140
rect 17175 4100 17592 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 17972 4137 18000 4168
rect 18230 4156 18236 4168
rect 18288 4156 18294 4208
rect 19242 4156 19248 4208
rect 19300 4196 19306 4208
rect 19300 4156 19334 4196
rect 17957 4131 18015 4137
rect 17957 4097 17969 4131
rect 18003 4097 18015 4131
rect 17957 4091 18015 4097
rect 18046 4088 18052 4140
rect 18104 4128 18110 4140
rect 18104 4100 18149 4128
rect 18104 4088 18110 4100
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 18417 4131 18475 4137
rect 18417 4128 18429 4131
rect 18380 4100 18429 4128
rect 18380 4088 18386 4100
rect 18417 4097 18429 4100
rect 18463 4097 18475 4131
rect 19306 4128 19334 4156
rect 27908 4168 28212 4196
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 19306 4100 19533 4128
rect 18417 4091 18475 4097
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 19521 4091 19579 4097
rect 23753 4131 23811 4137
rect 23753 4097 23765 4131
rect 23799 4128 23811 4131
rect 24670 4128 24676 4140
rect 23799 4100 24676 4128
rect 23799 4097 23811 4100
rect 23753 4091 23811 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 27154 4088 27160 4140
rect 27212 4128 27218 4140
rect 27522 4128 27528 4140
rect 27212 4100 27384 4128
rect 27483 4100 27528 4128
rect 27212 4088 27218 4100
rect 14369 4063 14427 4069
rect 14369 4029 14381 4063
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 14476 3992 14504 4023
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15620 4032 15669 4060
rect 15620 4020 15626 4032
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 16022 4020 16028 4072
rect 16080 4060 16086 4072
rect 16209 4063 16267 4069
rect 16080 4032 16125 4060
rect 16080 4020 16086 4032
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 16298 4060 16304 4072
rect 16255 4032 16304 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 16853 4063 16911 4069
rect 16853 4029 16865 4063
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 14332 3964 14504 3992
rect 16868 3992 16896 4023
rect 16942 4020 16948 4072
rect 17000 4060 17006 4072
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 17000 4032 17045 4060
rect 17144 4032 17233 4060
rect 17000 4020 17006 4032
rect 17034 3992 17040 4004
rect 16868 3964 17040 3992
rect 14332 3952 14338 3964
rect 17034 3952 17040 3964
rect 17092 3952 17098 4004
rect 11241 3896 12664 3924
rect 11241 3893 11253 3896
rect 11195 3887 11253 3893
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 12952 3896 13001 3924
rect 12952 3884 12958 3896
rect 12989 3893 13001 3896
rect 13035 3893 13047 3927
rect 12989 3887 13047 3893
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 17144 3924 17172 4032
rect 17221 4029 17233 4032
rect 17267 4029 17279 4063
rect 17678 4060 17684 4072
rect 17639 4032 17684 4060
rect 17221 4023 17279 4029
rect 17678 4020 17684 4032
rect 17736 4020 17742 4072
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4029 17923 4063
rect 18230 4060 18236 4072
rect 18191 4032 18236 4060
rect 17865 4023 17923 4029
rect 17880 3992 17908 4023
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 19061 4063 19119 4069
rect 19061 4029 19073 4063
rect 19107 4060 19119 4063
rect 19245 4063 19303 4069
rect 19245 4060 19257 4063
rect 19107 4032 19257 4060
rect 19107 4029 19119 4032
rect 19061 4023 19119 4029
rect 19245 4029 19257 4032
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 19702 4020 19708 4072
rect 19760 4060 19766 4072
rect 20533 4063 20591 4069
rect 20533 4060 20545 4063
rect 19760 4032 20545 4060
rect 19760 4020 19766 4032
rect 20533 4029 20545 4032
rect 20579 4029 20591 4063
rect 21174 4060 21180 4072
rect 21135 4032 21180 4060
rect 20533 4023 20591 4029
rect 21174 4020 21180 4032
rect 21232 4020 21238 4072
rect 23658 4060 23664 4072
rect 23619 4032 23664 4060
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 24578 4060 24584 4072
rect 24539 4032 24584 4060
rect 24578 4020 24584 4032
rect 24636 4020 24642 4072
rect 24857 4063 24915 4069
rect 24857 4029 24869 4063
rect 24903 4060 24915 4063
rect 26050 4060 26056 4072
rect 24903 4032 26056 4060
rect 24903 4029 24915 4032
rect 24857 4023 24915 4029
rect 26050 4020 26056 4032
rect 26108 4020 26114 4072
rect 27356 4060 27384 4100
rect 27522 4088 27528 4100
rect 27580 4088 27586 4140
rect 27908 4060 27936 4168
rect 28184 4128 28212 4168
rect 28537 4131 28595 4137
rect 28537 4128 28549 4131
rect 28184 4100 28549 4128
rect 28537 4097 28549 4100
rect 28583 4128 28595 4131
rect 28718 4128 28724 4140
rect 28583 4100 28724 4128
rect 28583 4097 28595 4100
rect 28537 4091 28595 4097
rect 28718 4088 28724 4100
rect 28776 4088 28782 4140
rect 29641 4131 29699 4137
rect 29641 4097 29653 4131
rect 29687 4128 29699 4131
rect 30193 4131 30251 4137
rect 30193 4128 30205 4131
rect 29687 4100 30205 4128
rect 29687 4097 29699 4100
rect 29641 4091 29699 4097
rect 30193 4097 30205 4100
rect 30239 4128 30251 4131
rect 30650 4128 30656 4140
rect 30239 4100 30656 4128
rect 30239 4097 30251 4100
rect 30193 4091 30251 4097
rect 30650 4088 30656 4100
rect 30708 4088 30714 4140
rect 30926 4128 30932 4140
rect 30887 4100 30932 4128
rect 30926 4088 30932 4100
rect 30984 4088 30990 4140
rect 27356 4032 27936 4060
rect 27982 4020 27988 4072
rect 28040 4060 28046 4072
rect 28261 4063 28319 4069
rect 28261 4060 28273 4063
rect 28040 4032 28273 4060
rect 28040 4020 28046 4032
rect 28261 4029 28273 4032
rect 28307 4029 28319 4063
rect 28261 4023 28319 4029
rect 28350 4020 28356 4072
rect 28408 4060 28414 4072
rect 28629 4063 28687 4069
rect 28408 4032 28453 4060
rect 28408 4020 28414 4032
rect 28629 4029 28641 4063
rect 28675 4060 28687 4063
rect 29546 4060 29552 4072
rect 28675 4032 29552 4060
rect 28675 4029 28687 4032
rect 28629 4023 28687 4029
rect 29546 4020 29552 4032
rect 29604 4020 29610 4072
rect 30374 4020 30380 4072
rect 30432 4060 30438 4072
rect 30558 4060 30564 4072
rect 30432 4032 30564 4060
rect 30432 4020 30438 4032
rect 30558 4020 30564 4032
rect 30616 4020 30622 4072
rect 19334 3992 19340 4004
rect 17880 3964 19340 3992
rect 19334 3952 19340 3964
rect 19392 3952 19398 4004
rect 21192 3992 21220 4020
rect 25869 3995 25927 4001
rect 25869 3992 25881 3995
rect 21192 3964 25881 3992
rect 25869 3961 25881 3964
rect 25915 3992 25927 3995
rect 28994 3992 29000 4004
rect 25915 3964 29000 3992
rect 25915 3961 25927 3964
rect 25869 3955 25927 3961
rect 28994 3952 29000 3964
rect 29052 3952 29058 4004
rect 16172 3896 17172 3924
rect 16172 3884 16178 3896
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 19061 3927 19119 3933
rect 19061 3924 19073 3927
rect 17552 3896 19073 3924
rect 17552 3884 17558 3896
rect 19061 3893 19073 3896
rect 19107 3893 19119 3927
rect 19061 3887 19119 3893
rect 1104 3834 32016 3856
rect 1104 3782 11253 3834
rect 11305 3782 11317 3834
rect 11369 3782 11381 3834
rect 11433 3782 11445 3834
rect 11497 3782 11509 3834
rect 11561 3782 21557 3834
rect 21609 3782 21621 3834
rect 21673 3782 21685 3834
rect 21737 3782 21749 3834
rect 21801 3782 21813 3834
rect 21865 3782 32016 3834
rect 1104 3760 32016 3782
rect 2866 3720 2872 3732
rect 2827 3692 2872 3720
rect 2866 3680 2872 3692
rect 2924 3720 2930 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 2924 3692 3893 3720
rect 2924 3680 2930 3692
rect 3881 3689 3893 3692
rect 3927 3689 3939 3723
rect 3881 3683 3939 3689
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 4212 3692 4445 3720
rect 4212 3680 4218 3692
rect 4433 3689 4445 3692
rect 4479 3720 4491 3723
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 4479 3692 5733 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 5721 3689 5733 3692
rect 5767 3689 5779 3723
rect 5721 3683 5779 3689
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3720 6515 3723
rect 6730 3720 6736 3732
rect 6503 3692 6736 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6730 3680 6736 3692
rect 6788 3720 6794 3732
rect 7098 3720 7104 3732
rect 6788 3692 7104 3720
rect 6788 3680 6794 3692
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 7926 3720 7932 3732
rect 7887 3692 7932 3720
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 11517 3723 11575 3729
rect 11517 3720 11529 3723
rect 11112 3692 11529 3720
rect 11112 3680 11118 3692
rect 11517 3689 11529 3692
rect 11563 3689 11575 3723
rect 11517 3683 11575 3689
rect 15194 3680 15200 3732
rect 15252 3720 15258 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 15252 3692 15669 3720
rect 15252 3680 15258 3692
rect 15657 3689 15669 3692
rect 15703 3720 15715 3723
rect 17678 3720 17684 3732
rect 15703 3692 16712 3720
rect 17639 3692 17684 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 5077 3655 5135 3661
rect 5077 3621 5089 3655
rect 5123 3652 5135 3655
rect 5810 3652 5816 3664
rect 5123 3624 5816 3652
rect 5123 3621 5135 3624
rect 5077 3615 5135 3621
rect 5810 3612 5816 3624
rect 5868 3612 5874 3664
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 7469 3655 7527 3661
rect 7469 3652 7481 3655
rect 7432 3624 7481 3652
rect 7432 3612 7438 3624
rect 7469 3621 7481 3624
rect 7515 3652 7527 3655
rect 8478 3652 8484 3664
rect 7515 3624 8484 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 9766 3652 9772 3664
rect 9324 3624 9772 3652
rect 9324 3593 9352 3624
rect 9766 3612 9772 3624
rect 9824 3652 9830 3664
rect 10870 3652 10876 3664
rect 9824 3624 10876 3652
rect 9824 3612 9830 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 14182 3652 14188 3664
rect 12406 3624 14188 3652
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 768 3556 1869 3584
rect 768 3244 796 3556
rect 1857 3553 1869 3556
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 9053 3587 9111 3593
rect 9053 3553 9065 3587
rect 9099 3584 9111 3587
rect 9309 3587 9367 3593
rect 9099 3556 9260 3584
rect 9099 3553 9111 3556
rect 9053 3547 9111 3553
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 7466 3516 7472 3528
rect 2179 3488 7472 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 9232 3516 9260 3556
rect 9309 3553 9321 3587
rect 9355 3553 9367 3587
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9309 3547 9367 3553
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10226 3584 10232 3596
rect 10187 3556 10232 3584
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3584 10563 3587
rect 10686 3584 10692 3596
rect 10551 3556 10692 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9232 3488 9781 3516
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 9769 3479 9827 3485
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10336 3392 10364 3547
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 12066 3584 12072 3596
rect 12027 3556 12072 3584
rect 12066 3544 12072 3556
rect 12124 3584 12130 3596
rect 12406 3584 12434 3624
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 14366 3612 14372 3664
rect 14424 3652 14430 3664
rect 14522 3655 14580 3661
rect 14522 3652 14534 3655
rect 14424 3624 14534 3652
rect 14424 3612 14430 3624
rect 14522 3621 14534 3624
rect 14568 3621 14580 3655
rect 14522 3615 14580 3621
rect 16684 3593 16712 3692
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 19242 3720 19248 3732
rect 18748 3692 19248 3720
rect 18748 3680 18754 3692
rect 19242 3680 19248 3692
rect 19300 3720 19306 3732
rect 19429 3723 19487 3729
rect 19429 3720 19441 3723
rect 19300 3692 19441 3720
rect 19300 3680 19306 3692
rect 19429 3689 19441 3692
rect 19475 3689 19487 3723
rect 19429 3683 19487 3689
rect 23566 3680 23572 3732
rect 23624 3720 23630 3732
rect 24578 3720 24584 3732
rect 23624 3692 24584 3720
rect 23624 3680 23630 3692
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 24670 3680 24676 3732
rect 24728 3720 24734 3732
rect 24728 3692 26188 3720
rect 24728 3680 24734 3692
rect 16942 3612 16948 3664
rect 17000 3652 17006 3664
rect 25222 3652 25228 3664
rect 17000 3624 18000 3652
rect 17000 3612 17006 3624
rect 12124 3556 12434 3584
rect 16669 3587 16727 3593
rect 12124 3544 12130 3556
rect 16669 3553 16681 3587
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 16758 3544 16764 3596
rect 16816 3584 16822 3596
rect 17972 3593 18000 3624
rect 19260 3624 20116 3652
rect 19260 3596 19288 3624
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 16816 3556 17877 3584
rect 16816 3544 16822 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 18877 3587 18935 3593
rect 18877 3584 18889 3587
rect 18279 3556 18889 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 18877 3553 18889 3556
rect 18923 3553 18935 3587
rect 18877 3547 18935 3553
rect 18969 3587 19027 3593
rect 18969 3553 18981 3587
rect 19015 3584 19027 3587
rect 19242 3584 19248 3596
rect 19015 3556 19248 3584
rect 19015 3553 19027 3556
rect 18969 3547 19027 3553
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19429 3587 19487 3593
rect 19429 3553 19441 3587
rect 19475 3584 19487 3587
rect 19521 3587 19579 3593
rect 19521 3584 19533 3587
rect 19475 3556 19533 3584
rect 19475 3553 19487 3556
rect 19429 3547 19487 3553
rect 19521 3553 19533 3556
rect 19567 3553 19579 3587
rect 19702 3584 19708 3596
rect 19663 3556 19708 3584
rect 19521 3547 19579 3553
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 19794 3544 19800 3596
rect 19852 3584 19858 3596
rect 20088 3593 20116 3624
rect 23860 3624 25228 3652
rect 20073 3587 20131 3593
rect 19852 3556 19897 3584
rect 19852 3544 19858 3556
rect 20073 3553 20085 3587
rect 20119 3553 20131 3587
rect 20073 3547 20131 3553
rect 22373 3587 22431 3593
rect 22373 3553 22385 3587
rect 22419 3584 22431 3587
rect 22830 3584 22836 3596
rect 22419 3556 22836 3584
rect 22419 3553 22431 3556
rect 22373 3547 22431 3553
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 23860 3593 23888 3624
rect 25222 3612 25228 3624
rect 25280 3612 25286 3664
rect 23845 3587 23903 3593
rect 23845 3584 23857 3587
rect 23492 3556 23857 3584
rect 13814 3516 13820 3528
rect 13775 3488 13820 3516
rect 13814 3476 13820 3488
rect 13872 3516 13878 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13872 3488 14289 3516
rect 13872 3476 13878 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17644 3488 18153 3516
rect 17644 3476 17650 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 19058 3516 19064 3528
rect 18380 3488 19064 3516
rect 18380 3476 18386 3488
rect 19058 3476 19064 3488
rect 19116 3516 19122 3528
rect 19886 3516 19892 3528
rect 19116 3488 19892 3516
rect 19116 3476 19122 3488
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3516 20315 3519
rect 20714 3516 20720 3528
rect 20303 3488 20720 3516
rect 20303 3485 20315 3488
rect 20257 3479 20315 3485
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 21910 3476 21916 3528
rect 21968 3516 21974 3528
rect 23492 3516 23520 3556
rect 23845 3553 23857 3556
rect 23891 3553 23903 3587
rect 24578 3584 24584 3596
rect 24539 3556 24584 3584
rect 23845 3547 23903 3553
rect 24578 3544 24584 3556
rect 24636 3544 24642 3596
rect 24670 3544 24676 3596
rect 24728 3584 24734 3596
rect 24949 3587 25007 3593
rect 24949 3584 24961 3587
rect 24728 3556 24961 3584
rect 24728 3544 24734 3556
rect 24949 3553 24961 3556
rect 24995 3553 25007 3587
rect 25130 3584 25136 3596
rect 25091 3556 25136 3584
rect 24949 3547 25007 3553
rect 25130 3544 25136 3556
rect 25188 3584 25194 3596
rect 25593 3587 25651 3593
rect 25593 3584 25605 3587
rect 25188 3556 25605 3584
rect 25188 3544 25194 3556
rect 25593 3553 25605 3556
rect 25639 3553 25651 3587
rect 25593 3547 25651 3553
rect 25682 3544 25688 3596
rect 25740 3584 25746 3596
rect 26160 3593 26188 3692
rect 26234 3680 26240 3732
rect 26292 3720 26298 3732
rect 27157 3723 27215 3729
rect 27157 3720 27169 3723
rect 26292 3692 27169 3720
rect 26292 3680 26298 3692
rect 27157 3689 27169 3692
rect 27203 3689 27215 3723
rect 27157 3683 27215 3689
rect 27246 3680 27252 3732
rect 27304 3720 27310 3732
rect 27798 3720 27804 3732
rect 27304 3692 27804 3720
rect 27304 3680 27310 3692
rect 27798 3680 27804 3692
rect 27856 3680 27862 3732
rect 28258 3680 28264 3732
rect 28316 3720 28322 3732
rect 30374 3720 30380 3732
rect 28316 3692 30380 3720
rect 28316 3680 28322 3692
rect 30374 3680 30380 3692
rect 30432 3680 30438 3732
rect 30558 3720 30564 3732
rect 30519 3692 30564 3720
rect 30558 3680 30564 3692
rect 30616 3680 30622 3732
rect 29641 3655 29699 3661
rect 29641 3621 29653 3655
rect 29687 3652 29699 3655
rect 30466 3652 30472 3664
rect 29687 3624 30472 3652
rect 29687 3621 29699 3624
rect 29641 3615 29699 3621
rect 30466 3612 30472 3624
rect 30524 3612 30530 3664
rect 25777 3587 25835 3593
rect 25777 3584 25789 3587
rect 25740 3556 25789 3584
rect 25740 3544 25746 3556
rect 25777 3553 25789 3556
rect 25823 3553 25835 3587
rect 25777 3547 25835 3553
rect 26145 3587 26203 3593
rect 26145 3553 26157 3587
rect 26191 3584 26203 3587
rect 27065 3587 27123 3593
rect 27065 3584 27077 3587
rect 26191 3556 27077 3584
rect 26191 3553 26203 3556
rect 26145 3547 26203 3553
rect 27065 3553 27077 3556
rect 27111 3553 27123 3587
rect 27065 3547 27123 3553
rect 27522 3544 27528 3596
rect 27580 3584 27586 3596
rect 27709 3587 27767 3593
rect 27709 3584 27721 3587
rect 27580 3556 27721 3584
rect 27580 3544 27586 3556
rect 27709 3553 27721 3556
rect 27755 3553 27767 3587
rect 27709 3547 27767 3553
rect 27798 3544 27804 3596
rect 27856 3584 27862 3596
rect 27965 3587 28023 3593
rect 27965 3584 27977 3587
rect 27856 3556 27977 3584
rect 27856 3544 27862 3556
rect 27965 3553 27977 3556
rect 28011 3553 28023 3587
rect 27965 3547 28023 3553
rect 28350 3544 28356 3596
rect 28408 3584 28414 3596
rect 28810 3584 28816 3596
rect 28408 3556 28816 3584
rect 28408 3544 28414 3556
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 30282 3544 30288 3596
rect 30340 3584 30346 3596
rect 31113 3587 31171 3593
rect 31113 3584 31125 3587
rect 30340 3556 31125 3584
rect 30340 3544 30346 3556
rect 31113 3553 31125 3556
rect 31159 3553 31171 3587
rect 31113 3547 31171 3553
rect 21968 3488 23520 3516
rect 23569 3519 23627 3525
rect 21968 3476 21974 3488
rect 23569 3485 23581 3519
rect 23615 3516 23627 3519
rect 24486 3516 24492 3528
rect 23615 3488 24492 3516
rect 23615 3485 23627 3488
rect 23569 3479 23627 3485
rect 24486 3476 24492 3488
rect 24544 3476 24550 3528
rect 24762 3516 24768 3528
rect 24723 3488 24768 3516
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3516 24915 3519
rect 25038 3516 25044 3528
rect 24903 3488 25044 3516
rect 24903 3485 24915 3488
rect 24857 3479 24915 3485
rect 25038 3476 25044 3488
rect 25096 3516 25102 3528
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 25096 3488 25881 3516
rect 25096 3476 25102 3488
rect 25869 3485 25881 3488
rect 25915 3485 25927 3519
rect 25869 3479 25927 3485
rect 25961 3519 26019 3525
rect 25961 3485 25973 3519
rect 26007 3485 26019 3519
rect 25961 3479 26019 3485
rect 18506 3408 18512 3460
rect 18564 3448 18570 3460
rect 21082 3448 21088 3460
rect 18564 3420 21088 3448
rect 18564 3408 18570 3420
rect 21082 3408 21088 3420
rect 21140 3408 21146 3460
rect 24780 3448 24808 3476
rect 25976 3448 26004 3479
rect 24780 3420 26004 3448
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 10318 3380 10324 3392
rect 8628 3352 10324 3380
rect 8628 3340 8634 3352
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 16761 3383 16819 3389
rect 16761 3380 16773 3383
rect 11848 3352 16773 3380
rect 11848 3340 11854 3352
rect 16761 3349 16773 3352
rect 16807 3349 16819 3383
rect 16761 3343 16819 3349
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 20717 3383 20775 3389
rect 20717 3380 20729 3383
rect 17920 3352 20729 3380
rect 17920 3340 17926 3352
rect 20717 3349 20729 3352
rect 20763 3349 20775 3383
rect 20717 3343 20775 3349
rect 22281 3383 22339 3389
rect 22281 3349 22293 3383
rect 22327 3380 22339 3383
rect 24302 3380 24308 3392
rect 22327 3352 24308 3380
rect 22327 3349 22339 3352
rect 22281 3343 22339 3349
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 24397 3383 24455 3389
rect 24397 3349 24409 3383
rect 24443 3380 24455 3383
rect 25038 3380 25044 3392
rect 24443 3352 25044 3380
rect 24443 3349 24455 3352
rect 24397 3343 24455 3349
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 25866 3340 25872 3392
rect 25924 3380 25930 3392
rect 26329 3383 26387 3389
rect 26329 3380 26341 3383
rect 25924 3352 26341 3380
rect 25924 3340 25930 3352
rect 26329 3349 26341 3352
rect 26375 3349 26387 3383
rect 26329 3343 26387 3349
rect 26602 3340 26608 3392
rect 26660 3380 26666 3392
rect 29089 3383 29147 3389
rect 29089 3380 29101 3383
rect 26660 3352 29101 3380
rect 26660 3340 26666 3352
rect 29089 3349 29101 3352
rect 29135 3349 29147 3383
rect 29089 3343 29147 3349
rect 31297 3383 31355 3389
rect 31297 3349 31309 3383
rect 31343 3380 31355 3383
rect 31343 3352 32352 3380
rect 31343 3349 31355 3352
rect 31297 3343 31355 3349
rect 1104 3290 32016 3312
rect 768 3216 888 3244
rect 1104 3238 6102 3290
rect 6154 3238 6166 3290
rect 6218 3238 6230 3290
rect 6282 3238 6294 3290
rect 6346 3238 6358 3290
rect 6410 3238 16405 3290
rect 16457 3238 16469 3290
rect 16521 3238 16533 3290
rect 16585 3238 16597 3290
rect 16649 3238 16661 3290
rect 16713 3238 26709 3290
rect 26761 3238 26773 3290
rect 26825 3238 26837 3290
rect 26889 3238 26901 3290
rect 26953 3238 26965 3290
rect 27017 3238 32016 3290
rect 32324 3244 32352 3352
rect 1104 3216 32016 3238
rect 32232 3216 32352 3244
rect 0 3108 800 3122
rect 860 3108 888 3216
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 2866 3176 2872 3188
rect 2731 3148 2872 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 2866 3136 2872 3148
rect 2924 3176 2930 3188
rect 3145 3179 3203 3185
rect 3145 3176 3157 3179
rect 2924 3148 3157 3176
rect 2924 3136 2930 3148
rect 3145 3145 3157 3148
rect 3191 3176 3203 3179
rect 3789 3179 3847 3185
rect 3789 3176 3801 3179
rect 3191 3148 3801 3176
rect 3191 3145 3203 3148
rect 3145 3139 3203 3145
rect 3789 3145 3801 3148
rect 3835 3176 3847 3179
rect 4154 3176 4160 3188
rect 3835 3148 4160 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 4154 3136 4160 3148
rect 4212 3176 4218 3188
rect 4341 3179 4399 3185
rect 4341 3176 4353 3179
rect 4212 3148 4353 3176
rect 4212 3136 4218 3148
rect 4341 3145 4353 3148
rect 4387 3176 4399 3179
rect 5442 3176 5448 3188
rect 4387 3148 5448 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 5442 3136 5448 3148
rect 5500 3176 5506 3188
rect 5537 3179 5595 3185
rect 5537 3176 5549 3179
rect 5500 3148 5549 3176
rect 5500 3136 5506 3148
rect 5537 3145 5549 3148
rect 5583 3176 5595 3179
rect 6089 3179 6147 3185
rect 6089 3176 6101 3179
rect 5583 3148 6101 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 6089 3145 6101 3148
rect 6135 3145 6147 3179
rect 7282 3176 7288 3188
rect 7243 3148 7288 3176
rect 6089 3139 6147 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 8478 3176 8484 3188
rect 8435 3148 8484 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9309 3179 9367 3185
rect 9309 3145 9321 3179
rect 9355 3176 9367 3179
rect 9858 3176 9864 3188
rect 9355 3148 9864 3176
rect 9355 3145 9367 3148
rect 9309 3139 9367 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 11204 3148 11621 3176
rect 11204 3136 11210 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 11609 3139 11667 3145
rect 12161 3179 12219 3185
rect 12161 3145 12173 3179
rect 12207 3176 12219 3179
rect 12434 3176 12440 3188
rect 12207 3148 12440 3176
rect 12207 3145 12219 3148
rect 12161 3139 12219 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3176 15991 3179
rect 16022 3176 16028 3188
rect 15979 3148 16028 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 16758 3176 16764 3188
rect 16719 3148 16764 3176
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 18230 3176 18236 3188
rect 17451 3148 18236 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 19334 3176 19340 3188
rect 19295 3148 19340 3176
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 24302 3136 24308 3188
rect 24360 3176 24366 3188
rect 26513 3179 26571 3185
rect 24360 3148 26464 3176
rect 24360 3136 24366 3148
rect 1489 3111 1547 3117
rect 1489 3108 1501 3111
rect 0 3080 1501 3108
rect 0 3066 800 3080
rect 1489 3077 1501 3080
rect 1535 3077 1547 3111
rect 1489 3071 1547 3077
rect 2774 3068 2780 3120
rect 2832 3108 2838 3120
rect 9030 3108 9036 3120
rect 2832 3080 9036 3108
rect 2832 3068 2838 3080
rect 9030 3068 9036 3080
rect 9088 3068 9094 3120
rect 10042 3068 10048 3120
rect 10100 3068 10106 3120
rect 10226 3108 10232 3120
rect 10152 3080 10232 3108
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5350 3040 5356 3052
rect 5123 3012 5356 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 7466 3040 7472 3052
rect 6871 3012 7472 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 10060 3040 10088 3068
rect 10152 3049 10180 3080
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 22186 3108 22192 3120
rect 22147 3080 22192 3108
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 24946 3108 24952 3120
rect 23400 3080 24952 3108
rect 9876 3012 10088 3040
rect 10137 3043 10195 3049
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 9674 2972 9680 2984
rect 9447 2944 9680 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9876 2981 9904 3012
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10594 3040 10600 3052
rect 10137 3003 10195 3009
rect 10244 3012 10600 3040
rect 10244 2984 10272 3012
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 13541 3043 13599 3049
rect 13541 3009 13553 3043
rect 13587 3040 13599 3043
rect 13814 3040 13820 3052
rect 13587 3012 13820 3040
rect 13587 3009 13599 3012
rect 13541 3003 13599 3009
rect 13814 3000 13820 3012
rect 13872 3040 13878 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 13872 3012 14565 3040
rect 13872 3000 13878 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 17957 3043 18015 3049
rect 17957 3009 17969 3043
rect 18003 3040 18015 3043
rect 18417 3043 18475 3049
rect 18003 3012 18276 3040
rect 18003 3009 18015 3012
rect 17957 3003 18015 3009
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2941 9919 2975
rect 10042 2972 10048 2984
rect 10003 2944 10048 2972
rect 9861 2935 9919 2941
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10424 2975 10482 2981
rect 10284 2944 10377 2972
rect 10284 2932 10290 2944
rect 10424 2941 10436 2975
rect 10470 2972 10482 2975
rect 10778 2972 10784 2984
rect 10470 2944 10784 2972
rect 10470 2941 10482 2944
rect 10424 2935 10482 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 2133 2907 2191 2913
rect 2133 2873 2145 2907
rect 2179 2904 2191 2907
rect 5994 2904 6000 2916
rect 2179 2876 6000 2904
rect 2179 2873 2191 2876
rect 2133 2867 2191 2873
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 10060 2904 10088 2932
rect 11716 2904 11744 2935
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13274 2975 13332 2981
rect 13274 2972 13286 2975
rect 12768 2944 13286 2972
rect 12768 2932 12774 2944
rect 13274 2941 13286 2944
rect 13320 2941 13332 2975
rect 13274 2935 13332 2941
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2941 16911 2975
rect 17310 2972 17316 2984
rect 17271 2944 17316 2972
rect 16853 2935 16911 2941
rect 11974 2904 11980 2916
rect 10060 2876 11980 2904
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 14820 2907 14878 2913
rect 14820 2873 14832 2907
rect 14866 2904 14878 2907
rect 16666 2904 16672 2916
rect 14866 2876 16672 2904
rect 14866 2873 14878 2876
rect 14820 2867 14878 2873
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 16868 2904 16896 2935
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2941 18199 2975
rect 18141 2935 18199 2941
rect 18046 2904 18052 2916
rect 16868 2876 18052 2904
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 10594 2836 10600 2848
rect 10555 2808 10600 2836
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 10962 2796 10968 2848
rect 11020 2836 11026 2848
rect 12710 2836 12716 2848
rect 11020 2808 12716 2836
rect 11020 2796 11026 2808
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 18156 2836 18184 2935
rect 18248 2904 18276 3012
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 19794 3040 19800 3052
rect 18463 3012 19800 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 23400 2984 23428 3080
rect 24762 3040 24768 3052
rect 24723 3012 24768 3040
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 24872 3049 24900 3080
rect 24946 3068 24952 3080
rect 25004 3068 25010 3120
rect 26436 3108 26464 3148
rect 26513 3145 26525 3179
rect 26559 3176 26571 3179
rect 27798 3176 27804 3188
rect 26559 3148 27804 3176
rect 26559 3145 26571 3148
rect 26513 3139 26571 3145
rect 27798 3136 27804 3148
rect 27856 3136 27862 3188
rect 28718 3136 28724 3188
rect 28776 3176 28782 3188
rect 29641 3179 29699 3185
rect 29641 3176 29653 3179
rect 28776 3148 29653 3176
rect 28776 3136 28782 3148
rect 29641 3145 29653 3148
rect 29687 3145 29699 3179
rect 30098 3176 30104 3188
rect 30059 3148 30104 3176
rect 29641 3139 29699 3145
rect 30098 3136 30104 3148
rect 30156 3136 30162 3188
rect 31018 3176 31024 3188
rect 30931 3148 31024 3176
rect 31018 3136 31024 3148
rect 31076 3176 31082 3188
rect 31294 3176 31300 3188
rect 31076 3148 31300 3176
rect 31076 3136 31082 3148
rect 31294 3136 31300 3148
rect 31352 3136 31358 3188
rect 32232 3108 32260 3216
rect 32320 3108 33120 3122
rect 26436 3080 29868 3108
rect 32232 3080 33120 3108
rect 24857 3043 24915 3049
rect 24857 3009 24869 3043
rect 24903 3009 24915 3043
rect 26050 3040 26056 3052
rect 26011 3012 26056 3040
rect 24857 3003 24915 3009
rect 26050 3000 26056 3012
rect 26108 3000 26114 3052
rect 26234 3000 26240 3052
rect 26292 3040 26298 3052
rect 28626 3040 28632 3052
rect 26292 3012 28488 3040
rect 28587 3012 28632 3040
rect 26292 3000 26298 3012
rect 18322 2932 18328 2984
rect 18380 2972 18386 2984
rect 18506 2972 18512 2984
rect 18380 2944 18425 2972
rect 18467 2944 18512 2972
rect 18380 2932 18386 2944
rect 18506 2932 18512 2944
rect 18564 2932 18570 2984
rect 18690 2972 18696 2984
rect 18651 2944 18696 2972
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19245 2975 19303 2981
rect 19245 2972 19257 2975
rect 19116 2944 19257 2972
rect 19116 2932 19122 2944
rect 19245 2941 19257 2944
rect 19291 2941 19303 2975
rect 19245 2935 19303 2941
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 22094 2972 22100 2984
rect 21499 2944 22100 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 22094 2932 22100 2944
rect 22152 2972 22158 2984
rect 22370 2972 22376 2984
rect 22152 2944 22376 2972
rect 22152 2932 22158 2944
rect 22370 2932 22376 2944
rect 22428 2932 22434 2984
rect 23382 2972 23388 2984
rect 23343 2944 23388 2972
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23624 2944 23673 2972
rect 23624 2932 23630 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 23750 2932 23756 2984
rect 23808 2972 23814 2984
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 23808 2944 24593 2972
rect 23808 2932 23814 2944
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 24949 2975 25007 2981
rect 24949 2941 24961 2975
rect 24995 2941 25007 2975
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 24949 2935 25007 2941
rect 21186 2907 21244 2913
rect 21186 2904 21198 2907
rect 18248 2876 21198 2904
rect 21186 2873 21198 2876
rect 21232 2873 21244 2907
rect 21186 2867 21244 2873
rect 21358 2864 21364 2916
rect 21416 2904 21422 2916
rect 21910 2904 21916 2916
rect 21416 2876 21916 2904
rect 21416 2864 21422 2876
rect 21910 2864 21916 2876
rect 21968 2904 21974 2916
rect 22005 2907 22063 2913
rect 22005 2904 22017 2907
rect 21968 2876 22017 2904
rect 21968 2864 21974 2876
rect 22005 2873 22017 2876
rect 22051 2873 22063 2907
rect 22005 2867 22063 2873
rect 22830 2864 22836 2916
rect 22888 2904 22894 2916
rect 24964 2904 24992 2935
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 25777 2975 25835 2981
rect 25777 2941 25789 2975
rect 25823 2941 25835 2975
rect 25958 2972 25964 2984
rect 25919 2944 25964 2972
rect 25777 2935 25835 2941
rect 22888 2876 24992 2904
rect 22888 2864 22894 2876
rect 19702 2836 19708 2848
rect 18156 2808 19708 2836
rect 19702 2796 19708 2808
rect 19760 2836 19766 2848
rect 20073 2839 20131 2845
rect 20073 2836 20085 2839
rect 19760 2808 20085 2836
rect 19760 2796 19766 2808
rect 20073 2805 20085 2808
rect 20119 2805 20131 2839
rect 20073 2799 20131 2805
rect 22186 2796 22192 2848
rect 22244 2836 22250 2848
rect 24397 2839 24455 2845
rect 24397 2836 24409 2839
rect 22244 2808 24409 2836
rect 22244 2796 22250 2808
rect 24397 2805 24409 2808
rect 24443 2805 24455 2839
rect 25792 2836 25820 2935
rect 25958 2932 25964 2944
rect 26016 2932 26022 2984
rect 26145 2975 26203 2981
rect 26145 2941 26157 2975
rect 26191 2941 26203 2975
rect 26145 2935 26203 2941
rect 26329 2975 26387 2981
rect 26329 2941 26341 2975
rect 26375 2972 26387 2975
rect 26602 2972 26608 2984
rect 26375 2944 26608 2972
rect 26375 2941 26387 2944
rect 26329 2935 26387 2941
rect 26160 2904 26188 2935
rect 26602 2932 26608 2944
rect 26660 2932 26666 2984
rect 26973 2975 27031 2981
rect 26973 2941 26985 2975
rect 27019 2972 27031 2975
rect 27154 2972 27160 2984
rect 27019 2944 27160 2972
rect 27019 2941 27031 2944
rect 26973 2935 27031 2941
rect 27154 2932 27160 2944
rect 27212 2932 27218 2984
rect 28460 2981 28488 3012
rect 28626 3000 28632 3012
rect 28684 3000 28690 3052
rect 29840 3040 29868 3080
rect 32320 3066 33120 3080
rect 29840 3012 29960 3040
rect 28445 2975 28503 2981
rect 28445 2941 28457 2975
rect 28491 2941 28503 2975
rect 28445 2935 28503 2941
rect 28534 2932 28540 2984
rect 28592 2972 28598 2984
rect 28712 2975 28770 2981
rect 28712 2972 28724 2975
rect 28592 2944 28724 2972
rect 28592 2932 28598 2944
rect 28712 2941 28724 2944
rect 28758 2941 28770 2975
rect 28712 2935 28770 2941
rect 28813 2975 28871 2981
rect 28813 2941 28825 2975
rect 28859 2972 28871 2975
rect 28902 2972 28908 2984
rect 28859 2944 28908 2972
rect 28859 2941 28871 2944
rect 28813 2935 28871 2941
rect 28902 2932 28908 2944
rect 28960 2932 28966 2984
rect 28997 2975 29055 2981
rect 28997 2941 29009 2975
rect 29043 2941 29055 2975
rect 28997 2935 29055 2941
rect 27338 2904 27344 2916
rect 26160 2876 27344 2904
rect 27338 2864 27344 2876
rect 27396 2864 27402 2916
rect 29012 2904 29040 2935
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29932 2981 29960 3012
rect 29549 2975 29607 2981
rect 29549 2972 29561 2975
rect 29144 2944 29561 2972
rect 29144 2932 29150 2944
rect 29549 2941 29561 2944
rect 29595 2941 29607 2975
rect 29549 2935 29607 2941
rect 29825 2975 29883 2981
rect 29825 2941 29837 2975
rect 29871 2941 29883 2975
rect 29825 2935 29883 2941
rect 29917 2975 29975 2981
rect 29917 2941 29929 2975
rect 29963 2941 29975 2975
rect 29917 2935 29975 2941
rect 29178 2904 29184 2916
rect 29012 2876 29184 2904
rect 29178 2864 29184 2876
rect 29236 2864 29242 2916
rect 26234 2836 26240 2848
rect 25792 2808 26240 2836
rect 24397 2799 24455 2805
rect 26234 2796 26240 2808
rect 26292 2836 26298 2848
rect 27062 2836 27068 2848
rect 26292 2808 27068 2836
rect 26292 2796 26298 2808
rect 27062 2796 27068 2808
rect 27120 2836 27126 2848
rect 27203 2839 27261 2845
rect 27203 2836 27215 2839
rect 27120 2808 27215 2836
rect 27120 2796 27126 2808
rect 27203 2805 27215 2808
rect 27249 2836 27261 2839
rect 28074 2836 28080 2848
rect 27249 2808 28080 2836
rect 27249 2805 27261 2808
rect 27203 2799 27261 2805
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 28166 2796 28172 2848
rect 28224 2836 28230 2848
rect 28261 2839 28319 2845
rect 28261 2836 28273 2839
rect 28224 2808 28273 2836
rect 28224 2796 28230 2808
rect 28261 2805 28273 2808
rect 28307 2805 28319 2839
rect 28261 2799 28319 2805
rect 28810 2796 28816 2848
rect 28868 2836 28874 2848
rect 29840 2836 29868 2935
rect 28868 2808 29868 2836
rect 28868 2796 28874 2808
rect 1104 2746 32016 2768
rect 1104 2694 11253 2746
rect 11305 2694 11317 2746
rect 11369 2694 11381 2746
rect 11433 2694 11445 2746
rect 11497 2694 11509 2746
rect 11561 2694 21557 2746
rect 21609 2694 21621 2746
rect 21673 2694 21685 2746
rect 21737 2694 21749 2746
rect 21801 2694 21813 2746
rect 21865 2694 32016 2746
rect 1104 2672 32016 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 3142 2632 3148 2644
rect 2731 2604 3148 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 4154 2632 4160 2644
rect 3292 2604 3337 2632
rect 4115 2604 4160 2632
rect 3292 2592 3298 2604
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 5629 2635 5687 2641
rect 5629 2632 5641 2635
rect 5500 2604 5641 2632
rect 5500 2592 5506 2604
rect 5629 2601 5641 2604
rect 5675 2632 5687 2635
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 5675 2604 6377 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7156 2604 7389 2632
rect 7156 2592 7162 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 8570 2632 8576 2644
rect 8435 2604 8576 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 12710 2632 12716 2644
rect 9732 2604 10649 2632
rect 12671 2604 12716 2632
rect 9732 2592 9738 2604
rect 9524 2567 9582 2573
rect 9524 2533 9536 2567
rect 9570 2564 9582 2567
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9570 2536 10241 2564
rect 9570 2533 9582 2536
rect 9524 2527 9582 2533
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 10376 2468 10425 2496
rect 10376 2456 10382 2468
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 10621 2496 10649 2604
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 14185 2635 14243 2641
rect 14185 2601 14197 2635
rect 14231 2632 14243 2635
rect 14274 2632 14280 2644
rect 14231 2604 14280 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 16666 2632 16672 2644
rect 16627 2604 16672 2632
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 17218 2632 17224 2644
rect 17052 2604 17224 2632
rect 10686 2524 10692 2576
rect 10744 2564 10750 2576
rect 13170 2564 13176 2576
rect 10744 2536 11008 2564
rect 10744 2524 10750 2536
rect 10778 2496 10784 2508
rect 10621 2468 10784 2496
rect 10413 2459 10471 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 10980 2505 11008 2536
rect 11716 2536 13176 2564
rect 11716 2508 11744 2536
rect 13170 2524 13176 2536
rect 13228 2564 13234 2576
rect 15930 2564 15936 2576
rect 13228 2536 14136 2564
rect 13228 2524 13234 2536
rect 10965 2499 11023 2505
rect 10965 2465 10977 2499
rect 11011 2496 11023 2499
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11011 2468 11529 2496
rect 11011 2465 11023 2468
rect 10965 2459 11023 2465
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11698 2496 11704 2508
rect 11659 2468 11704 2496
rect 11517 2459 11575 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 14108 2505 14136 2536
rect 14568 2536 15936 2564
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 12032 2468 12081 2496
rect 12032 2456 12038 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 13633 2499 13691 2505
rect 13633 2465 13645 2499
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10284 2400 10609 2428
rect 10284 2388 10290 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10612 2360 10640 2391
rect 10686 2388 10692 2440
rect 10744 2428 10750 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 10744 2400 11805 2428
rect 10744 2388 10750 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 13648 2428 13676 2459
rect 14568 2428 14596 2536
rect 15930 2524 15936 2536
rect 15988 2564 15994 2576
rect 15988 2536 16896 2564
rect 15988 2524 15994 2536
rect 15004 2499 15062 2505
rect 15004 2465 15016 2499
rect 15050 2496 15062 2499
rect 15378 2496 15384 2508
rect 15050 2468 15384 2496
rect 15050 2465 15062 2468
rect 15004 2459 15062 2465
rect 15378 2456 15384 2468
rect 15436 2456 15442 2508
rect 16868 2505 16896 2536
rect 17052 2505 17080 2604
rect 17218 2592 17224 2604
rect 17276 2632 17282 2644
rect 22002 2632 22008 2644
rect 17276 2604 18000 2632
rect 17276 2592 17282 2604
rect 17770 2564 17776 2576
rect 17144 2536 17776 2564
rect 17144 2505 17172 2536
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 17972 2564 18000 2604
rect 21836 2604 22008 2632
rect 19794 2564 19800 2576
rect 17972 2536 18276 2564
rect 17402 2505 17408 2508
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 17221 2499 17279 2505
rect 17221 2465 17233 2499
rect 17267 2496 17279 2499
rect 17267 2468 17356 2496
rect 17267 2465 17279 2468
rect 17221 2459 17279 2465
rect 14734 2428 14740 2440
rect 13648 2400 14596 2428
rect 14695 2400 14740 2428
rect 11885 2391 11943 2397
rect 11900 2360 11928 2391
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 17144 2428 17172 2459
rect 16080 2400 17172 2428
rect 16080 2388 16086 2400
rect 10612 2332 11928 2360
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 16117 2363 16175 2369
rect 16117 2360 16129 2363
rect 15988 2332 16129 2360
rect 15988 2320 15994 2332
rect 16117 2329 16129 2332
rect 16163 2360 16175 2363
rect 17328 2360 17356 2468
rect 17401 2459 17408 2505
rect 17460 2496 17466 2508
rect 17865 2499 17923 2505
rect 17865 2496 17877 2499
rect 17460 2468 17877 2496
rect 17402 2456 17408 2459
rect 17460 2456 17466 2468
rect 17865 2465 17877 2468
rect 17911 2465 17923 2499
rect 18046 2496 18052 2508
rect 18007 2468 18052 2496
rect 17865 2459 17923 2465
rect 18046 2456 18052 2468
rect 18104 2456 18110 2508
rect 18248 2505 18276 2536
rect 19352 2536 19800 2564
rect 18233 2499 18291 2505
rect 18233 2465 18245 2499
rect 18279 2496 18291 2499
rect 18414 2496 18420 2508
rect 18279 2465 18312 2496
rect 18375 2468 18420 2496
rect 18233 2459 18312 2465
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18141 2431 18199 2437
rect 18141 2428 18153 2431
rect 18012 2400 18153 2428
rect 18012 2388 18018 2400
rect 18141 2397 18153 2400
rect 18187 2397 18199 2431
rect 18284 2428 18312 2459
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 18690 2456 18696 2508
rect 18748 2496 18754 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18748 2468 19073 2496
rect 18748 2456 18754 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19242 2496 19248 2508
rect 19203 2468 19248 2496
rect 19061 2459 19119 2465
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 19352 2505 19380 2536
rect 19794 2524 19800 2536
rect 19852 2524 19858 2576
rect 19337 2499 19395 2505
rect 19337 2465 19349 2499
rect 19383 2465 19395 2499
rect 19337 2459 19395 2465
rect 19429 2499 19487 2505
rect 19429 2465 19441 2499
rect 19475 2496 19487 2499
rect 19518 2496 19524 2508
rect 19475 2468 19524 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 19444 2428 19472 2459
rect 19518 2456 19524 2468
rect 19576 2456 19582 2508
rect 19613 2499 19671 2505
rect 19613 2465 19625 2499
rect 19659 2465 19671 2499
rect 19613 2459 19671 2465
rect 19628 2428 19656 2459
rect 20254 2456 20260 2508
rect 20312 2496 20318 2508
rect 21836 2505 21864 2604
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 23201 2635 23259 2641
rect 23201 2601 23213 2635
rect 23247 2632 23259 2635
rect 23658 2632 23664 2644
rect 23247 2604 23664 2632
rect 23247 2601 23259 2604
rect 23201 2595 23259 2601
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 23753 2635 23811 2641
rect 23753 2601 23765 2635
rect 23799 2632 23811 2635
rect 24578 2632 24584 2644
rect 23799 2604 24584 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 24854 2592 24860 2644
rect 24912 2592 24918 2644
rect 26050 2592 26056 2644
rect 26108 2632 26114 2644
rect 28534 2632 28540 2644
rect 26108 2604 28540 2632
rect 26108 2592 26114 2604
rect 28534 2592 28540 2604
rect 28592 2592 28598 2644
rect 29546 2632 29552 2644
rect 29507 2604 29552 2632
rect 29546 2592 29552 2604
rect 29604 2592 29610 2644
rect 30377 2635 30435 2641
rect 30377 2601 30389 2635
rect 30423 2632 30435 2635
rect 30926 2632 30932 2644
rect 30423 2604 30932 2632
rect 30423 2601 30435 2604
rect 30377 2595 30435 2601
rect 30926 2592 30932 2604
rect 30984 2592 30990 2644
rect 22088 2567 22146 2573
rect 22088 2533 22100 2567
rect 22134 2564 22146 2567
rect 22186 2564 22192 2576
rect 22134 2536 22192 2564
rect 22134 2533 22146 2536
rect 22088 2527 22146 2533
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 24872 2564 24900 2592
rect 24872 2536 25176 2564
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 20312 2468 21833 2496
rect 20312 2456 20318 2468
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 24877 2499 24935 2505
rect 24877 2465 24889 2499
rect 24923 2496 24935 2499
rect 25038 2496 25044 2508
rect 24923 2468 25044 2496
rect 24923 2465 24935 2468
rect 24877 2459 24935 2465
rect 25038 2456 25044 2468
rect 25096 2456 25102 2508
rect 25148 2505 25176 2536
rect 26602 2524 26608 2576
rect 26660 2564 26666 2576
rect 26660 2536 28488 2564
rect 26660 2524 26666 2536
rect 25133 2499 25191 2505
rect 25133 2465 25145 2499
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 25222 2456 25228 2508
rect 25280 2496 25286 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 25280 2468 25605 2496
rect 25280 2456 25286 2468
rect 25593 2465 25605 2468
rect 25639 2496 25651 2499
rect 26973 2499 27031 2505
rect 26973 2496 26985 2499
rect 25639 2468 26985 2496
rect 25639 2465 25651 2468
rect 25593 2459 25651 2465
rect 26973 2465 26985 2468
rect 27019 2465 27031 2499
rect 26973 2459 27031 2465
rect 27249 2499 27307 2505
rect 27249 2465 27261 2499
rect 27295 2496 27307 2499
rect 27338 2496 27344 2508
rect 27295 2468 27344 2496
rect 27295 2465 27307 2468
rect 27249 2459 27307 2465
rect 27338 2456 27344 2468
rect 27396 2456 27402 2508
rect 28074 2456 28080 2508
rect 28132 2496 28138 2508
rect 28258 2496 28264 2508
rect 28132 2468 28264 2496
rect 28132 2456 28138 2468
rect 28258 2456 28264 2468
rect 28316 2456 28322 2508
rect 28460 2505 28488 2536
rect 28552 2505 28580 2592
rect 28445 2499 28503 2505
rect 28445 2465 28457 2499
rect 28491 2465 28503 2499
rect 28445 2459 28503 2465
rect 28537 2499 28595 2505
rect 28537 2465 28549 2499
rect 28583 2465 28595 2499
rect 28810 2496 28816 2508
rect 28771 2468 28816 2496
rect 28537 2459 28595 2465
rect 28810 2456 28816 2468
rect 28868 2496 28874 2508
rect 29457 2499 29515 2505
rect 29457 2496 29469 2499
rect 28868 2468 29469 2496
rect 28868 2456 28874 2468
rect 29457 2465 29469 2468
rect 29503 2465 29515 2499
rect 29457 2459 29515 2465
rect 18284 2400 19472 2428
rect 19518 2400 19656 2428
rect 20993 2431 21051 2437
rect 18141 2391 18199 2397
rect 16163 2332 17356 2360
rect 16163 2329 16175 2332
rect 16117 2323 16175 2329
rect 18046 2320 18052 2372
rect 18104 2360 18110 2372
rect 18874 2360 18880 2372
rect 18104 2332 18880 2360
rect 18104 2320 18110 2332
rect 18874 2320 18880 2332
rect 18932 2360 18938 2372
rect 18932 2332 19334 2360
rect 18932 2320 18938 2332
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 10686 2292 10692 2304
rect 10192 2264 10692 2292
rect 10192 2252 10198 2264
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 12250 2292 12256 2304
rect 12211 2264 12256 2292
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 13541 2295 13599 2301
rect 13541 2261 13553 2295
rect 13587 2292 13599 2295
rect 17034 2292 17040 2304
rect 13587 2264 17040 2292
rect 13587 2261 13599 2264
rect 13541 2255 13599 2261
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 18598 2292 18604 2304
rect 18559 2264 18604 2292
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 19306 2292 19334 2332
rect 19518 2292 19546 2400
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 21358 2428 21364 2440
rect 21315 2400 21364 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 19610 2320 19616 2372
rect 19668 2360 19674 2372
rect 21008 2360 21036 2391
rect 21358 2388 21364 2400
rect 21416 2388 21422 2440
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2397 25927 2431
rect 27356 2428 27384 2456
rect 28626 2428 28632 2440
rect 27356 2400 28632 2428
rect 25869 2391 25927 2397
rect 19668 2332 21036 2360
rect 19668 2320 19674 2332
rect 19794 2292 19800 2304
rect 19306 2264 19546 2292
rect 19755 2264 19800 2292
rect 19794 2252 19800 2264
rect 19852 2252 19858 2304
rect 24762 2252 24768 2304
rect 24820 2292 24826 2304
rect 25774 2292 25780 2304
rect 24820 2264 25780 2292
rect 24820 2252 24826 2264
rect 25774 2252 25780 2264
rect 25832 2292 25838 2304
rect 25884 2292 25912 2391
rect 28626 2388 28632 2400
rect 28684 2388 28690 2440
rect 28258 2320 28264 2372
rect 28316 2360 28322 2372
rect 29178 2360 29184 2372
rect 28316 2332 29184 2360
rect 28316 2320 28322 2332
rect 29178 2320 29184 2332
rect 29236 2320 29242 2372
rect 30098 2320 30104 2372
rect 30156 2360 30162 2372
rect 30837 2363 30895 2369
rect 30837 2360 30849 2363
rect 30156 2332 30849 2360
rect 30156 2320 30162 2332
rect 30837 2329 30849 2332
rect 30883 2329 30895 2363
rect 30837 2323 30895 2329
rect 25832 2264 25912 2292
rect 25832 2252 25838 2264
rect 27338 2252 27344 2304
rect 27396 2292 27402 2304
rect 28997 2295 29055 2301
rect 28997 2292 29009 2295
rect 27396 2264 29009 2292
rect 27396 2252 27402 2264
rect 28997 2261 29009 2264
rect 29043 2261 29055 2295
rect 28997 2255 29055 2261
rect 1104 2202 32016 2224
rect 1104 2150 6102 2202
rect 6154 2150 6166 2202
rect 6218 2150 6230 2202
rect 6282 2150 6294 2202
rect 6346 2150 6358 2202
rect 6410 2150 16405 2202
rect 16457 2150 16469 2202
rect 16521 2150 16533 2202
rect 16585 2150 16597 2202
rect 16649 2150 16661 2202
rect 16713 2150 26709 2202
rect 26761 2150 26773 2202
rect 26825 2150 26837 2202
rect 26889 2150 26901 2202
rect 26953 2150 26965 2202
rect 27017 2150 32016 2202
rect 1104 2128 32016 2150
rect 1486 2088 1492 2100
rect 1447 2060 1492 2088
rect 1486 2048 1492 2060
rect 1544 2048 1550 2100
rect 2130 2048 2136 2100
rect 2188 2088 2194 2100
rect 2501 2091 2559 2097
rect 2501 2088 2513 2091
rect 2188 2060 2513 2088
rect 2188 2048 2194 2060
rect 2501 2057 2513 2060
rect 2547 2057 2559 2091
rect 2501 2051 2559 2057
rect 3145 2091 3203 2097
rect 3145 2057 3157 2091
rect 3191 2088 3203 2091
rect 3326 2088 3332 2100
rect 3191 2060 3332 2088
rect 3191 2057 3203 2060
rect 3145 2051 3203 2057
rect 3326 2048 3332 2060
rect 3384 2048 3390 2100
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 3789 2091 3847 2097
rect 3789 2088 3801 2091
rect 3476 2060 3801 2088
rect 3476 2048 3482 2060
rect 3789 2057 3801 2060
rect 3835 2057 3847 2091
rect 5994 2088 6000 2100
rect 5955 2060 6000 2088
rect 3789 2051 3847 2057
rect 5994 2048 6000 2060
rect 6052 2088 6058 2100
rect 9582 2088 9588 2100
rect 6052 2060 8432 2088
rect 9543 2060 9588 2088
rect 6052 2048 6058 2060
rect 8404 2032 8432 2060
rect 9582 2048 9588 2060
rect 9640 2048 9646 2100
rect 12066 2088 12072 2100
rect 9692 2060 12072 2088
rect 2041 2023 2099 2029
rect 2041 1989 2053 2023
rect 2087 2020 2099 2023
rect 2590 2020 2596 2032
rect 2087 1992 2596 2020
rect 2087 1989 2099 1992
rect 2041 1983 2099 1989
rect 2590 1980 2596 1992
rect 2648 1980 2654 2032
rect 5442 1980 5448 2032
rect 5500 2020 5506 2032
rect 6825 2023 6883 2029
rect 6825 2020 6837 2023
rect 5500 1992 6837 2020
rect 5500 1980 5506 1992
rect 6825 1989 6837 1992
rect 6871 2020 6883 2023
rect 7377 2023 7435 2029
rect 7377 2020 7389 2023
rect 6871 1992 7389 2020
rect 6871 1989 6883 1992
rect 6825 1983 6883 1989
rect 7377 1989 7389 1992
rect 7423 1989 7435 2023
rect 8386 2020 8392 2032
rect 8299 1992 8392 2020
rect 7377 1983 7435 1989
rect 8386 1980 8392 1992
rect 8444 2020 8450 2032
rect 9033 2023 9091 2029
rect 9033 2020 9045 2023
rect 8444 1992 9045 2020
rect 8444 1980 8450 1992
rect 9033 1989 9045 1992
rect 9079 2020 9091 2023
rect 9122 2020 9128 2032
rect 9079 1992 9128 2020
rect 9079 1989 9091 1992
rect 9033 1983 9091 1989
rect 9122 1980 9128 1992
rect 9180 2020 9186 2032
rect 9692 2020 9720 2060
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 12713 2091 12771 2097
rect 12713 2057 12725 2091
rect 12759 2088 12771 2091
rect 12986 2088 12992 2100
rect 12759 2060 12992 2088
rect 12759 2057 12771 2060
rect 12713 2051 12771 2057
rect 12986 2048 12992 2060
rect 13044 2048 13050 2100
rect 13262 2088 13268 2100
rect 13223 2060 13268 2088
rect 13262 2048 13268 2060
rect 13320 2048 13326 2100
rect 16761 2091 16819 2097
rect 16761 2057 16773 2091
rect 16807 2088 16819 2091
rect 16850 2088 16856 2100
rect 16807 2060 16856 2088
rect 16807 2057 16819 2060
rect 16761 2051 16819 2057
rect 16850 2048 16856 2060
rect 16908 2048 16914 2100
rect 18782 2088 18788 2100
rect 17144 2060 18788 2088
rect 9180 1992 9720 2020
rect 9180 1980 9186 1992
rect 10042 1980 10048 2032
rect 10100 2020 10106 2032
rect 10597 2023 10655 2029
rect 10597 2020 10609 2023
rect 10100 1992 10609 2020
rect 10100 1980 10106 1992
rect 10597 1989 10609 1992
rect 10643 1989 10655 2023
rect 10597 1983 10655 1989
rect 15657 2023 15715 2029
rect 15657 1989 15669 2023
rect 15703 2020 15715 2023
rect 17144 2020 17172 2060
rect 18782 2048 18788 2060
rect 18840 2048 18846 2100
rect 19242 2048 19248 2100
rect 19300 2088 19306 2100
rect 19613 2091 19671 2097
rect 19613 2088 19625 2091
rect 19300 2060 19625 2088
rect 19300 2048 19306 2060
rect 19613 2057 19625 2060
rect 19659 2057 19671 2091
rect 22830 2088 22836 2100
rect 22791 2060 22836 2088
rect 19613 2051 19671 2057
rect 22830 2048 22836 2060
rect 22888 2048 22894 2100
rect 23106 2048 23112 2100
rect 23164 2088 23170 2100
rect 23293 2091 23351 2097
rect 23293 2088 23305 2091
rect 23164 2060 23305 2088
rect 23164 2048 23170 2060
rect 23293 2057 23305 2060
rect 23339 2057 23351 2091
rect 23293 2051 23351 2057
rect 24397 2091 24455 2097
rect 24397 2057 24409 2091
rect 24443 2088 24455 2091
rect 24670 2088 24676 2100
rect 24443 2060 24676 2088
rect 24443 2057 24455 2060
rect 24397 2051 24455 2057
rect 24670 2048 24676 2060
rect 24728 2048 24734 2100
rect 24854 2048 24860 2100
rect 24912 2088 24918 2100
rect 26326 2088 26332 2100
rect 24912 2060 25820 2088
rect 26287 2060 26332 2088
rect 24912 2048 24918 2060
rect 15703 1992 17172 2020
rect 15703 1989 15715 1992
rect 15657 1983 15715 1989
rect 13814 1912 13820 1964
rect 13872 1952 13878 1964
rect 14093 1955 14151 1961
rect 14093 1952 14105 1955
rect 13872 1924 14105 1952
rect 13872 1912 13878 1924
rect 14093 1921 14105 1924
rect 14139 1952 14151 1955
rect 14734 1952 14740 1964
rect 14139 1924 14740 1952
rect 14139 1921 14151 1924
rect 14093 1915 14151 1921
rect 14734 1912 14740 1924
rect 14792 1912 14798 1964
rect 25792 1961 25820 2060
rect 26326 2048 26332 2060
rect 26384 2048 26390 2100
rect 28445 2091 28503 2097
rect 28445 2057 28457 2091
rect 28491 2088 28503 2091
rect 28810 2088 28816 2100
rect 28491 2060 28816 2088
rect 28491 2057 28503 2060
rect 28445 2051 28503 2057
rect 28810 2048 28816 2060
rect 28868 2048 28874 2100
rect 28997 2091 29055 2097
rect 28997 2057 29009 2091
rect 29043 2088 29055 2091
rect 30006 2088 30012 2100
rect 29043 2060 30012 2088
rect 29043 2057 29055 2060
rect 28997 2051 29055 2057
rect 30006 2048 30012 2060
rect 30064 2048 30070 2100
rect 25777 1955 25835 1961
rect 25777 1921 25789 1955
rect 25823 1952 25835 1955
rect 26418 1952 26424 1964
rect 25823 1924 26424 1952
rect 25823 1921 25835 1924
rect 25777 1915 25835 1921
rect 26418 1912 26424 1924
rect 26476 1952 26482 1964
rect 26476 1924 27108 1952
rect 26476 1912 26482 1924
rect 10870 1844 10876 1896
rect 10928 1884 10934 1896
rect 11977 1887 12035 1893
rect 11977 1884 11989 1887
rect 10928 1856 11989 1884
rect 10928 1844 10934 1856
rect 11977 1853 11989 1856
rect 12023 1853 12035 1887
rect 14366 1884 14372 1896
rect 14327 1856 14372 1884
rect 11977 1847 12035 1853
rect 14366 1844 14372 1856
rect 14424 1844 14430 1896
rect 15746 1844 15752 1896
rect 15804 1884 15810 1896
rect 16669 1887 16727 1893
rect 16669 1884 16681 1887
rect 15804 1856 16681 1884
rect 15804 1844 15810 1856
rect 16669 1853 16681 1856
rect 16715 1853 16727 1887
rect 16669 1847 16727 1853
rect 18437 1887 18495 1893
rect 18437 1853 18449 1887
rect 18483 1884 18495 1887
rect 18598 1884 18604 1896
rect 18483 1856 18604 1884
rect 18483 1853 18495 1856
rect 18437 1847 18495 1853
rect 18598 1844 18604 1856
rect 18656 1844 18662 1896
rect 18693 1887 18751 1893
rect 18693 1853 18705 1887
rect 18739 1884 18751 1887
rect 20254 1884 20260 1896
rect 18739 1856 20260 1884
rect 18739 1853 18751 1856
rect 18693 1847 18751 1853
rect 20254 1844 20260 1856
rect 20312 1884 20318 1896
rect 20993 1887 21051 1893
rect 20993 1884 21005 1887
rect 20312 1856 21005 1884
rect 20312 1844 20318 1856
rect 20993 1853 21005 1856
rect 21039 1884 21051 1887
rect 21453 1887 21511 1893
rect 21453 1884 21465 1887
rect 21039 1856 21465 1884
rect 21039 1853 21051 1856
rect 20993 1847 21051 1853
rect 21453 1853 21465 1856
rect 21499 1853 21511 1887
rect 21453 1847 21511 1853
rect 25521 1887 25579 1893
rect 25521 1853 25533 1887
rect 25567 1884 25579 1887
rect 25866 1884 25872 1896
rect 25567 1856 25872 1884
rect 25567 1853 25579 1856
rect 25521 1847 25579 1853
rect 25866 1844 25872 1856
rect 25924 1844 25930 1896
rect 27080 1893 27108 1924
rect 26237 1887 26295 1893
rect 26237 1853 26249 1887
rect 26283 1853 26295 1887
rect 26237 1847 26295 1853
rect 27065 1887 27123 1893
rect 27065 1853 27077 1887
rect 27111 1884 27123 1887
rect 27111 1856 27568 1884
rect 27111 1853 27123 1856
rect 27065 1847 27123 1853
rect 11732 1819 11790 1825
rect 11732 1785 11744 1819
rect 11778 1816 11790 1819
rect 12250 1816 12256 1828
rect 11778 1788 12256 1816
rect 11778 1785 11790 1788
rect 11732 1779 11790 1785
rect 12250 1776 12256 1788
rect 12308 1776 12314 1828
rect 20714 1816 20720 1828
rect 20772 1825 20778 1828
rect 20684 1788 20720 1816
rect 20714 1776 20720 1788
rect 20772 1779 20784 1825
rect 21720 1819 21778 1825
rect 21720 1785 21732 1819
rect 21766 1816 21778 1819
rect 22646 1816 22652 1828
rect 21766 1788 22652 1816
rect 21766 1785 21778 1788
rect 21720 1779 21778 1785
rect 20772 1776 20778 1779
rect 22646 1776 22652 1788
rect 22704 1776 22710 1828
rect 25682 1776 25688 1828
rect 25740 1816 25746 1828
rect 26252 1816 26280 1847
rect 27540 1828 27568 1856
rect 27338 1825 27344 1828
rect 27332 1816 27344 1825
rect 25740 1788 26280 1816
rect 27299 1788 27344 1816
rect 25740 1776 25746 1788
rect 27332 1779 27344 1788
rect 27338 1776 27344 1779
rect 27396 1776 27402 1828
rect 27522 1776 27528 1828
rect 27580 1776 27586 1828
rect 28994 1776 29000 1828
rect 29052 1816 29058 1828
rect 29549 1819 29607 1825
rect 29549 1816 29561 1819
rect 29052 1788 29561 1816
rect 29052 1776 29058 1788
rect 29549 1785 29561 1788
rect 29595 1816 29607 1819
rect 30098 1816 30104 1828
rect 29595 1788 30104 1816
rect 29595 1785 29607 1788
rect 29549 1779 29607 1785
rect 30098 1776 30104 1788
rect 30156 1776 30162 1828
rect 10137 1751 10195 1757
rect 10137 1717 10149 1751
rect 10183 1748 10195 1751
rect 16206 1748 16212 1760
rect 10183 1720 16212 1748
rect 10183 1717 10195 1720
rect 10137 1711 10195 1717
rect 16206 1708 16212 1720
rect 16264 1708 16270 1760
rect 16942 1708 16948 1760
rect 17000 1748 17006 1760
rect 17310 1748 17316 1760
rect 17000 1720 17316 1748
rect 17000 1708 17006 1720
rect 17310 1708 17316 1720
rect 17368 1748 17374 1760
rect 18414 1748 18420 1760
rect 17368 1720 18420 1748
rect 17368 1708 17374 1720
rect 18414 1708 18420 1720
rect 18472 1708 18478 1760
rect 30926 1748 30932 1760
rect 30887 1720 30932 1748
rect 30926 1708 30932 1720
rect 30984 1708 30990 1760
rect 1104 1658 32016 1680
rect 1104 1606 11253 1658
rect 11305 1606 11317 1658
rect 11369 1606 11381 1658
rect 11433 1606 11445 1658
rect 11497 1606 11509 1658
rect 11561 1606 21557 1658
rect 21609 1606 21621 1658
rect 21673 1606 21685 1658
rect 21737 1606 21749 1658
rect 21801 1606 21813 1658
rect 21865 1606 32016 1658
rect 1104 1584 32016 1606
rect 8021 1547 8079 1553
rect 8021 1513 8033 1547
rect 8067 1544 8079 1547
rect 8386 1544 8392 1556
rect 8067 1516 8392 1544
rect 8067 1513 8079 1516
rect 8021 1507 8079 1513
rect 8386 1504 8392 1516
rect 8444 1544 8450 1556
rect 8573 1547 8631 1553
rect 8573 1544 8585 1547
rect 8444 1516 8585 1544
rect 8444 1504 8450 1516
rect 8573 1513 8585 1516
rect 8619 1544 8631 1547
rect 9122 1544 9128 1556
rect 8619 1516 9128 1544
rect 8619 1513 8631 1516
rect 8573 1507 8631 1513
rect 9122 1504 9128 1516
rect 9180 1504 9186 1556
rect 9585 1547 9643 1553
rect 9585 1513 9597 1547
rect 9631 1544 9643 1547
rect 9674 1544 9680 1556
rect 9631 1516 9680 1544
rect 9631 1513 9643 1516
rect 9585 1507 9643 1513
rect 9674 1504 9680 1516
rect 9732 1504 9738 1556
rect 12713 1547 12771 1553
rect 12713 1513 12725 1547
rect 12759 1544 12771 1547
rect 13354 1544 13360 1556
rect 12759 1516 13360 1544
rect 12759 1513 12771 1516
rect 12713 1507 12771 1513
rect 13354 1504 13360 1516
rect 13412 1504 13418 1556
rect 14366 1504 14372 1556
rect 14424 1544 14430 1556
rect 14553 1547 14611 1553
rect 14553 1544 14565 1547
rect 14424 1516 14565 1544
rect 14424 1504 14430 1516
rect 14553 1513 14565 1516
rect 14599 1513 14611 1547
rect 15930 1544 15936 1556
rect 14553 1507 14611 1513
rect 15580 1516 15936 1544
rect 10594 1436 10600 1488
rect 10652 1476 10658 1488
rect 10698 1479 10756 1485
rect 10698 1476 10710 1479
rect 10652 1448 10710 1476
rect 10652 1436 10658 1448
rect 10698 1445 10710 1448
rect 10744 1445 10756 1479
rect 13814 1476 13820 1488
rect 10698 1439 10756 1445
rect 13188 1448 13820 1476
rect 1854 1408 1860 1420
rect 1815 1380 1860 1408
rect 1854 1368 1860 1380
rect 1912 1368 1918 1420
rect 10870 1368 10876 1420
rect 10928 1408 10934 1420
rect 10965 1411 11023 1417
rect 10965 1408 10977 1411
rect 10928 1380 10977 1408
rect 10928 1368 10934 1380
rect 10965 1377 10977 1380
rect 11011 1377 11023 1411
rect 10965 1371 11023 1377
rect 2777 1343 2835 1349
rect 2777 1309 2789 1343
rect 2823 1340 2835 1343
rect 2958 1340 2964 1352
rect 2823 1312 2964 1340
rect 2823 1309 2835 1312
rect 2777 1303 2835 1309
rect 2958 1300 2964 1312
rect 3016 1300 3022 1352
rect 10980 1340 11008 1371
rect 13188 1352 13216 1448
rect 13814 1436 13820 1448
rect 13872 1436 13878 1488
rect 13440 1411 13498 1417
rect 13440 1377 13452 1411
rect 13486 1408 13498 1411
rect 13998 1408 14004 1420
rect 13486 1380 14004 1408
rect 13486 1377 13498 1380
rect 13440 1371 13498 1377
rect 13998 1368 14004 1380
rect 14056 1368 14062 1420
rect 15580 1417 15608 1516
rect 15930 1504 15936 1516
rect 15988 1504 15994 1556
rect 16761 1547 16819 1553
rect 16761 1513 16773 1547
rect 16807 1513 16819 1547
rect 18874 1544 18880 1556
rect 18835 1516 18880 1544
rect 16761 1507 16819 1513
rect 16776 1476 16804 1507
rect 18874 1504 18880 1516
rect 18932 1504 18938 1556
rect 21450 1504 21456 1556
rect 21508 1544 21514 1556
rect 21821 1547 21879 1553
rect 21821 1544 21833 1547
rect 21508 1516 21833 1544
rect 21508 1504 21514 1516
rect 21821 1513 21833 1516
rect 21867 1513 21879 1547
rect 21821 1507 21879 1513
rect 24489 1547 24547 1553
rect 24489 1513 24501 1547
rect 24535 1544 24547 1547
rect 28994 1544 29000 1556
rect 24535 1516 26234 1544
rect 28955 1516 29000 1544
rect 24535 1513 24547 1516
rect 24489 1507 24547 1513
rect 17310 1476 17316 1488
rect 15948 1448 17316 1476
rect 15948 1417 15976 1448
rect 17310 1436 17316 1448
rect 17368 1476 17374 1488
rect 19058 1476 19064 1488
rect 17368 1448 19064 1476
rect 17368 1436 17374 1448
rect 19058 1436 19064 1448
rect 19116 1436 19122 1488
rect 19794 1436 19800 1488
rect 19852 1476 19858 1488
rect 19990 1479 20048 1485
rect 19990 1476 20002 1479
rect 19852 1448 20002 1476
rect 19852 1436 19858 1448
rect 19990 1445 20002 1448
rect 20036 1445 20048 1479
rect 26206 1476 26234 1516
rect 28994 1504 29000 1516
rect 29052 1544 29058 1556
rect 29457 1547 29515 1553
rect 29457 1544 29469 1547
rect 29052 1516 29469 1544
rect 29052 1504 29058 1516
rect 29457 1513 29469 1516
rect 29503 1513 29515 1547
rect 30006 1544 30012 1556
rect 29967 1516 30012 1544
rect 29457 1507 29515 1513
rect 30006 1504 30012 1516
rect 30064 1504 30070 1556
rect 29086 1476 29092 1488
rect 19990 1439 20048 1445
rect 23308 1448 24440 1476
rect 26206 1448 29092 1476
rect 15565 1411 15623 1417
rect 15565 1377 15577 1411
rect 15611 1377 15623 1411
rect 15565 1371 15623 1377
rect 15933 1411 15991 1417
rect 15933 1377 15945 1411
rect 15979 1377 15991 1411
rect 15933 1371 15991 1377
rect 16117 1411 16175 1417
rect 16117 1377 16129 1411
rect 16163 1408 16175 1411
rect 16758 1408 16764 1420
rect 16163 1380 16764 1408
rect 16163 1377 16175 1380
rect 16117 1371 16175 1377
rect 16758 1368 16764 1380
rect 16816 1408 16822 1420
rect 17402 1408 17408 1420
rect 16816 1380 17408 1408
rect 16816 1368 16822 1380
rect 17402 1368 17408 1380
rect 17460 1368 17466 1420
rect 17494 1368 17500 1420
rect 17552 1408 17558 1420
rect 17874 1411 17932 1417
rect 17874 1408 17886 1411
rect 17552 1380 17886 1408
rect 17552 1368 17558 1380
rect 17874 1377 17886 1380
rect 17920 1377 17932 1411
rect 17874 1371 17932 1377
rect 22830 1368 22836 1420
rect 22888 1408 22894 1420
rect 23308 1417 23336 1448
rect 24412 1417 24440 1448
rect 29086 1436 29092 1448
rect 29144 1436 29150 1488
rect 22925 1411 22983 1417
rect 22925 1408 22937 1411
rect 22888 1380 22937 1408
rect 22888 1368 22894 1380
rect 22925 1377 22937 1380
rect 22971 1377 22983 1411
rect 22925 1371 22983 1377
rect 23293 1411 23351 1417
rect 23293 1377 23305 1411
rect 23339 1377 23351 1411
rect 23293 1371 23351 1377
rect 23477 1411 23535 1417
rect 23477 1377 23489 1411
rect 23523 1408 23535 1411
rect 24397 1411 24455 1417
rect 23523 1380 24348 1408
rect 23523 1377 23535 1380
rect 23477 1371 23535 1377
rect 13170 1340 13176 1352
rect 10980 1312 13176 1340
rect 13170 1300 13176 1312
rect 13228 1300 13234 1352
rect 15378 1340 15384 1352
rect 15339 1312 15384 1340
rect 15378 1300 15384 1312
rect 15436 1300 15442 1352
rect 15749 1343 15807 1349
rect 15749 1309 15761 1343
rect 15795 1309 15807 1343
rect 15749 1303 15807 1309
rect 15841 1343 15899 1349
rect 15841 1309 15853 1343
rect 15887 1340 15899 1343
rect 16022 1340 16028 1352
rect 15887 1312 16028 1340
rect 15887 1309 15899 1312
rect 15841 1303 15899 1309
rect 2133 1275 2191 1281
rect 2133 1241 2145 1275
rect 2179 1272 2191 1275
rect 7374 1272 7380 1284
rect 2179 1244 7380 1272
rect 2179 1241 2191 1244
rect 2133 1235 2191 1241
rect 7374 1232 7380 1244
rect 7432 1232 7438 1284
rect 11609 1275 11667 1281
rect 11609 1241 11621 1275
rect 11655 1272 11667 1275
rect 12158 1272 12164 1284
rect 11655 1244 12164 1272
rect 11655 1241 11667 1244
rect 11609 1235 11667 1241
rect 12158 1232 12164 1244
rect 12216 1232 12222 1284
rect 15764 1272 15792 1303
rect 16022 1300 16028 1312
rect 16080 1300 16086 1352
rect 18141 1343 18199 1349
rect 18141 1309 18153 1343
rect 18187 1340 18199 1343
rect 19150 1340 19156 1352
rect 18187 1312 19156 1340
rect 18187 1309 18199 1312
rect 18141 1303 18199 1309
rect 19150 1300 19156 1312
rect 19208 1300 19214 1352
rect 20254 1340 20260 1352
rect 20215 1312 20260 1340
rect 20254 1300 20260 1312
rect 20312 1300 20318 1352
rect 22646 1300 22652 1352
rect 22704 1340 22710 1352
rect 22741 1343 22799 1349
rect 22741 1340 22753 1343
rect 22704 1312 22753 1340
rect 22704 1300 22710 1312
rect 22741 1309 22753 1312
rect 22787 1309 22799 1343
rect 22741 1303 22799 1309
rect 23109 1343 23167 1349
rect 23109 1309 23121 1343
rect 23155 1309 23167 1343
rect 23109 1303 23167 1309
rect 23201 1343 23259 1349
rect 23201 1309 23213 1343
rect 23247 1340 23259 1343
rect 23382 1340 23388 1352
rect 23247 1312 23388 1340
rect 23247 1309 23259 1312
rect 23201 1303 23259 1309
rect 17126 1272 17132 1284
rect 15764 1244 17132 1272
rect 17126 1232 17132 1244
rect 17184 1232 17190 1284
rect 23124 1272 23152 1303
rect 23382 1300 23388 1312
rect 23440 1300 23446 1352
rect 24320 1340 24348 1380
rect 24397 1377 24409 1411
rect 24443 1408 24455 1411
rect 24578 1408 24584 1420
rect 24443 1380 24584 1408
rect 24443 1377 24455 1380
rect 24397 1371 24455 1377
rect 24578 1368 24584 1380
rect 24636 1368 24642 1420
rect 25130 1408 25136 1420
rect 24688 1380 25136 1408
rect 24688 1340 24716 1380
rect 25130 1368 25136 1380
rect 25188 1368 25194 1420
rect 25590 1368 25596 1420
rect 25648 1408 25654 1420
rect 26154 1411 26212 1417
rect 26154 1408 26166 1411
rect 25648 1380 26166 1408
rect 25648 1368 25654 1380
rect 26154 1377 26166 1380
rect 26200 1377 26212 1411
rect 26418 1408 26424 1420
rect 26379 1380 26424 1408
rect 26154 1371 26212 1377
rect 26418 1368 26424 1380
rect 26476 1368 26482 1420
rect 28166 1368 28172 1420
rect 28224 1417 28230 1420
rect 28224 1408 28236 1417
rect 28224 1380 28269 1408
rect 28224 1371 28236 1380
rect 28224 1368 28230 1371
rect 30466 1368 30472 1420
rect 30524 1408 30530 1420
rect 31113 1411 31171 1417
rect 31113 1408 31125 1411
rect 30524 1380 31125 1408
rect 30524 1368 30530 1380
rect 31113 1377 31125 1380
rect 31159 1377 31171 1411
rect 31113 1371 31171 1377
rect 24320 1312 24716 1340
rect 28445 1343 28503 1349
rect 28445 1309 28457 1343
rect 28491 1309 28503 1343
rect 28445 1303 28503 1309
rect 24762 1272 24768 1284
rect 23124 1244 24768 1272
rect 24762 1232 24768 1244
rect 24820 1232 24826 1284
rect 10594 1164 10600 1216
rect 10652 1204 10658 1216
rect 12069 1207 12127 1213
rect 12069 1204 12081 1207
rect 10652 1176 12081 1204
rect 10652 1164 10658 1176
rect 12069 1173 12081 1176
rect 12115 1173 12127 1207
rect 12069 1167 12127 1173
rect 12986 1164 12992 1216
rect 13044 1204 13050 1216
rect 20717 1207 20775 1213
rect 20717 1204 20729 1207
rect 13044 1176 20729 1204
rect 13044 1164 13050 1176
rect 20717 1173 20729 1176
rect 20763 1173 20775 1207
rect 20717 1167 20775 1173
rect 25041 1207 25099 1213
rect 25041 1173 25053 1207
rect 25087 1204 25099 1207
rect 25498 1204 25504 1216
rect 25087 1176 25504 1204
rect 25087 1173 25099 1176
rect 25041 1167 25099 1173
rect 25498 1164 25504 1176
rect 25556 1204 25562 1216
rect 25682 1204 25688 1216
rect 25556 1176 25688 1204
rect 25556 1164 25562 1176
rect 25682 1164 25688 1176
rect 25740 1164 25746 1216
rect 26142 1164 26148 1216
rect 26200 1204 26206 1216
rect 27065 1207 27123 1213
rect 27065 1204 27077 1207
rect 26200 1176 27077 1204
rect 26200 1164 26206 1176
rect 27065 1173 27077 1176
rect 27111 1173 27123 1207
rect 27065 1167 27123 1173
rect 27522 1164 27528 1216
rect 27580 1204 27586 1216
rect 28460 1204 28488 1303
rect 27580 1176 28488 1204
rect 31297 1207 31355 1213
rect 27580 1164 27586 1176
rect 31297 1173 31309 1207
rect 31343 1204 31355 1207
rect 31343 1176 32076 1204
rect 31343 1173 31355 1176
rect 31297 1167 31355 1173
rect 1104 1114 32016 1136
rect 0 1068 800 1082
rect 0 1040 1072 1068
rect 1104 1062 6102 1114
rect 6154 1062 6166 1114
rect 6218 1062 6230 1114
rect 6282 1062 6294 1114
rect 6346 1062 6358 1114
rect 6410 1062 16405 1114
rect 16457 1062 16469 1114
rect 16521 1062 16533 1114
rect 16585 1062 16597 1114
rect 16649 1062 16661 1114
rect 16713 1062 26709 1114
rect 26761 1062 26773 1114
rect 26825 1062 26837 1114
rect 26889 1062 26901 1114
rect 26953 1062 26965 1114
rect 27017 1062 32016 1114
rect 1104 1040 32016 1062
rect 32048 1068 32076 1176
rect 32320 1068 33120 1082
rect 32048 1040 33120 1068
rect 0 1026 800 1040
rect 1044 1000 1072 1040
rect 32320 1026 33120 1040
rect 1581 1003 1639 1009
rect 1581 1000 1593 1003
rect 1044 972 1593 1000
rect 1581 969 1593 972
rect 1627 1000 1639 1003
rect 1854 1000 1860 1012
rect 1627 972 1860 1000
rect 1627 969 1639 972
rect 1581 963 1639 969
rect 1854 960 1860 972
rect 1912 960 1918 1012
rect 8386 1000 8392 1012
rect 8347 972 8392 1000
rect 8386 960 8392 972
rect 8444 960 8450 1012
rect 10413 1003 10471 1009
rect 10413 969 10425 1003
rect 10459 1000 10471 1003
rect 14458 1000 14464 1012
rect 10459 972 14464 1000
rect 10459 969 10471 972
rect 10413 963 10471 969
rect 14458 960 14464 972
rect 14516 960 14522 1012
rect 15289 1003 15347 1009
rect 15289 969 15301 1003
rect 15335 1000 15347 1003
rect 15838 1000 15844 1012
rect 15335 972 15844 1000
rect 15335 969 15347 972
rect 15289 963 15347 969
rect 15838 960 15844 972
rect 15896 960 15902 1012
rect 16025 1003 16083 1009
rect 16025 969 16037 1003
rect 16071 1000 16083 1003
rect 16114 1000 16120 1012
rect 16071 972 16120 1000
rect 16071 969 16083 972
rect 16025 963 16083 969
rect 16114 960 16120 972
rect 16172 960 16178 1012
rect 17494 1000 17500 1012
rect 17455 972 17500 1000
rect 17494 960 17500 972
rect 17552 960 17558 1012
rect 18049 1003 18107 1009
rect 18049 969 18061 1003
rect 18095 1000 18107 1003
rect 18506 1000 18512 1012
rect 18095 972 18512 1000
rect 18095 969 18107 972
rect 18049 963 18107 969
rect 18506 960 18512 972
rect 18564 960 18570 1012
rect 18601 1003 18659 1009
rect 18601 969 18613 1003
rect 18647 1000 18659 1003
rect 18966 1000 18972 1012
rect 18647 972 18972 1000
rect 18647 969 18659 972
rect 18601 963 18659 969
rect 18966 960 18972 972
rect 19024 960 19030 1012
rect 19426 1000 19432 1012
rect 19387 972 19432 1000
rect 19426 960 19432 972
rect 19484 960 19490 1012
rect 20717 1003 20775 1009
rect 20717 969 20729 1003
rect 20763 1000 20775 1003
rect 20806 1000 20812 1012
rect 20763 972 20812 1000
rect 20763 969 20775 972
rect 20717 963 20775 969
rect 20806 960 20812 972
rect 20864 960 20870 1012
rect 20898 960 20904 1012
rect 20956 1000 20962 1012
rect 21821 1003 21879 1009
rect 21821 1000 21833 1003
rect 20956 972 21833 1000
rect 20956 960 20962 972
rect 21821 969 21833 972
rect 21867 969 21879 1003
rect 21821 963 21879 969
rect 22278 960 22284 1012
rect 22336 1000 22342 1012
rect 22373 1003 22431 1009
rect 22373 1000 22385 1003
rect 22336 972 22385 1000
rect 22336 960 22342 972
rect 22373 969 22385 972
rect 22419 969 22431 1003
rect 22373 963 22431 969
rect 22738 960 22744 1012
rect 22796 1000 22802 1012
rect 27617 1003 27675 1009
rect 27617 1000 27629 1003
rect 22796 972 27629 1000
rect 22796 960 22802 972
rect 27617 969 27629 972
rect 27663 1000 27675 1003
rect 28077 1003 28135 1009
rect 28077 1000 28089 1003
rect 27663 972 28089 1000
rect 27663 969 27675 972
rect 27617 963 27675 969
rect 28077 969 28089 972
rect 28123 969 28135 1003
rect 28077 963 28135 969
rect 28721 1003 28779 1009
rect 28721 969 28733 1003
rect 28767 1000 28779 1003
rect 28994 1000 29000 1012
rect 28767 972 29000 1000
rect 28767 969 28779 972
rect 28721 963 28779 969
rect 28994 960 29000 972
rect 29052 960 29058 1012
rect 7837 935 7895 941
rect 7837 901 7849 935
rect 7883 932 7895 935
rect 8294 932 8300 944
rect 7883 904 8300 932
rect 7883 901 7895 904
rect 7837 895 7895 901
rect 8294 892 8300 904
rect 8352 892 8358 944
rect 11698 892 11704 944
rect 11756 932 11762 944
rect 11793 935 11851 941
rect 11793 932 11805 935
rect 11756 904 11805 932
rect 11756 892 11762 904
rect 11793 901 11805 904
rect 11839 901 11851 935
rect 11793 895 11851 901
rect 13998 892 14004 944
rect 14056 932 14062 944
rect 14093 935 14151 941
rect 14093 932 14105 935
rect 14056 904 14105 932
rect 14056 892 14062 904
rect 14093 901 14105 904
rect 14139 901 14151 935
rect 14093 895 14151 901
rect 20070 892 20076 944
rect 20128 932 20134 944
rect 21177 935 21235 941
rect 21177 932 21189 935
rect 20128 904 21189 932
rect 20128 892 20134 904
rect 21177 901 21189 904
rect 21223 901 21235 935
rect 23014 932 23020 944
rect 22975 904 23020 932
rect 21177 895 21235 901
rect 23014 892 23020 904
rect 23072 892 23078 944
rect 23198 892 23204 944
rect 23256 932 23262 944
rect 23477 935 23535 941
rect 23477 932 23489 935
rect 23256 904 23489 932
rect 23256 892 23262 904
rect 23477 901 23489 904
rect 23523 901 23535 935
rect 23477 895 23535 901
rect 25501 935 25559 941
rect 25501 901 25513 935
rect 25547 932 25559 935
rect 25590 932 25596 944
rect 25547 904 25596 932
rect 25547 901 25559 904
rect 25501 895 25559 901
rect 25590 892 25596 904
rect 25648 892 25654 944
rect 25682 892 25688 944
rect 25740 932 25746 944
rect 29549 935 29607 941
rect 29549 932 29561 935
rect 25740 904 29561 932
rect 25740 892 25746 904
rect 29549 901 29561 904
rect 29595 901 29607 935
rect 29549 895 29607 901
rect 8312 796 8340 892
rect 13170 864 13176 876
rect 13131 836 13176 864
rect 13170 824 13176 836
rect 13228 824 13234 876
rect 16022 824 16028 876
rect 16080 864 16086 876
rect 17037 867 17095 873
rect 17037 864 17049 867
rect 16080 836 17049 864
rect 16080 824 16086 836
rect 17037 833 17049 836
rect 17083 833 17095 867
rect 17037 827 17095 833
rect 17129 867 17187 873
rect 17129 833 17141 867
rect 17175 864 17187 867
rect 17218 864 17224 876
rect 17175 836 17224 864
rect 17175 833 17187 836
rect 17129 827 17187 833
rect 17218 824 17224 836
rect 17276 824 17282 876
rect 25958 864 25964 876
rect 25919 836 25964 864
rect 25958 824 25964 836
rect 26016 824 26022 876
rect 27065 867 27123 873
rect 27065 833 27077 867
rect 27111 864 27123 867
rect 27154 864 27160 876
rect 27111 836 27160 864
rect 27111 833 27123 836
rect 27065 827 27123 833
rect 27154 824 27160 836
rect 27212 824 27218 876
rect 9401 799 9459 805
rect 9401 796 9413 799
rect 8312 768 9413 796
rect 9401 765 9413 768
rect 9447 765 9459 799
rect 12894 796 12900 808
rect 12952 805 12958 808
rect 12864 768 12900 796
rect 9401 759 9459 765
rect 12894 756 12900 768
rect 12952 759 12964 805
rect 12952 756 12958 759
rect 13906 756 13912 808
rect 13964 796 13970 808
rect 14277 799 14335 805
rect 14277 796 14289 799
rect 13964 768 14289 796
rect 13964 756 13970 768
rect 14277 765 14289 768
rect 14323 765 14335 799
rect 15930 796 15936 808
rect 15891 768 15936 796
rect 14277 759 14335 765
rect 15930 756 15936 768
rect 15988 756 15994 808
rect 16758 796 16764 808
rect 16719 768 16764 796
rect 16758 756 16764 768
rect 16816 756 16822 808
rect 16942 796 16948 808
rect 16903 768 16948 796
rect 16942 756 16948 768
rect 17000 756 17006 808
rect 17310 796 17316 808
rect 17271 768 17316 796
rect 17310 756 17316 768
rect 17368 756 17374 808
rect 19426 756 19432 808
rect 19484 796 19490 808
rect 19613 799 19671 805
rect 19613 796 19625 799
rect 19484 768 19625 796
rect 19484 756 19490 768
rect 19613 765 19625 768
rect 19659 796 19671 799
rect 19659 768 22094 796
rect 19659 765 19671 768
rect 19613 759 19671 765
rect 7285 731 7343 737
rect 7285 697 7297 731
rect 7331 728 7343 731
rect 13924 728 13952 756
rect 7331 700 13952 728
rect 22066 728 22094 768
rect 24026 756 24032 808
rect 24084 796 24090 808
rect 24765 799 24823 805
rect 24765 796 24777 799
rect 24084 768 24777 796
rect 24084 756 24090 768
rect 24765 765 24777 768
rect 24811 765 24823 799
rect 24946 796 24952 808
rect 24907 768 24952 796
rect 24765 759 24823 765
rect 24946 756 24952 768
rect 25004 756 25010 808
rect 25498 756 25504 808
rect 25556 796 25562 808
rect 25685 799 25743 805
rect 25685 796 25697 799
rect 25556 768 25697 796
rect 25556 756 25562 768
rect 25685 765 25697 768
rect 25731 765 25743 799
rect 25685 759 25743 765
rect 25774 756 25780 808
rect 25832 805 25838 808
rect 25832 799 25881 805
rect 25832 765 25835 799
rect 25869 765 25881 799
rect 25832 759 25881 765
rect 26049 799 26107 805
rect 26049 765 26061 799
rect 26095 796 26107 799
rect 26142 796 26148 808
rect 26095 768 26148 796
rect 26095 765 26107 768
rect 26049 759 26107 765
rect 25832 756 25838 759
rect 26142 756 26148 768
rect 26200 756 26206 808
rect 26234 756 26240 808
rect 26292 796 26298 808
rect 26292 768 26337 796
rect 26292 756 26298 768
rect 26694 756 26700 808
rect 26752 796 26758 808
rect 30926 796 30932 808
rect 26752 768 30932 796
rect 26752 756 26758 768
rect 30926 756 30932 768
rect 30984 756 30990 808
rect 30101 731 30159 737
rect 30101 728 30113 731
rect 22066 700 24900 728
rect 7331 697 7343 700
rect 7285 691 7343 697
rect 9490 660 9496 672
rect 9451 632 9496 660
rect 9490 620 9496 632
rect 9548 620 9554 672
rect 10965 663 11023 669
rect 10965 629 10977 663
rect 11011 660 11023 663
rect 14642 660 14648 672
rect 11011 632 14648 660
rect 11011 629 11023 632
rect 10965 623 11023 629
rect 14642 620 14648 632
rect 14700 620 14706 672
rect 20162 660 20168 672
rect 20123 632 20168 660
rect 20162 620 20168 632
rect 20220 620 20226 672
rect 24872 660 24900 700
rect 26206 700 30113 728
rect 26206 672 26234 700
rect 30101 697 30113 700
rect 30147 697 30159 731
rect 30101 691 30159 697
rect 25682 660 25688 672
rect 24872 632 25688 660
rect 25682 620 25688 632
rect 25740 620 25746 672
rect 26142 620 26148 672
rect 26200 632 26234 672
rect 26200 620 26206 632
rect 1104 570 32016 592
rect 1104 518 11253 570
rect 11305 518 11317 570
rect 11369 518 11381 570
rect 11433 518 11445 570
rect 11497 518 11509 570
rect 11561 518 21557 570
rect 21609 518 21621 570
rect 21673 518 21685 570
rect 21737 518 21749 570
rect 21801 518 21813 570
rect 21865 518 32016 570
rect 1104 496 32016 518
rect 9490 416 9496 468
rect 9548 456 9554 468
rect 23014 456 23020 468
rect 9548 428 23020 456
rect 9548 416 9554 428
rect 23014 416 23020 428
rect 23072 416 23078 468
rect 24946 416 24952 468
rect 25004 456 25010 468
rect 26142 456 26148 468
rect 25004 428 26148 456
rect 25004 416 25010 428
rect 26142 416 26148 428
rect 26200 416 26206 468
rect 20162 348 20168 400
rect 20220 388 20226 400
rect 26694 388 26700 400
rect 20220 360 26700 388
rect 20220 348 20226 360
rect 26694 348 26700 360
rect 26752 348 26758 400
<< via1 >>
rect 11253 48390 11305 48442
rect 11317 48390 11369 48442
rect 11381 48390 11433 48442
rect 11445 48390 11497 48442
rect 11509 48390 11561 48442
rect 21557 48390 21609 48442
rect 21621 48390 21673 48442
rect 21685 48390 21737 48442
rect 21749 48390 21801 48442
rect 21813 48390 21865 48442
rect 8484 48152 8536 48204
rect 15844 48195 15896 48204
rect 15844 48161 15853 48195
rect 15853 48161 15887 48195
rect 15887 48161 15896 48195
rect 15844 48152 15896 48161
rect 24768 48152 24820 48204
rect 31300 48152 31352 48204
rect 8300 48016 8352 48068
rect 14924 48016 14976 48068
rect 5724 47948 5776 48000
rect 11612 47948 11664 48000
rect 15936 47991 15988 48000
rect 15936 47957 15945 47991
rect 15945 47957 15979 47991
rect 15979 47957 15988 47991
rect 15936 47948 15988 47957
rect 16764 47948 16816 48000
rect 24860 48016 24912 48068
rect 20076 47991 20128 48000
rect 20076 47957 20085 47991
rect 20085 47957 20119 47991
rect 20119 47957 20128 47991
rect 20076 47948 20128 47957
rect 6102 47846 6154 47898
rect 6166 47846 6218 47898
rect 6230 47846 6282 47898
rect 6294 47846 6346 47898
rect 6358 47846 6410 47898
rect 16405 47846 16457 47898
rect 16469 47846 16521 47898
rect 16533 47846 16585 47898
rect 16597 47846 16649 47898
rect 16661 47846 16713 47898
rect 26709 47846 26761 47898
rect 26773 47846 26825 47898
rect 26837 47846 26889 47898
rect 26901 47846 26953 47898
rect 26965 47846 27017 47898
rect 18328 47744 18380 47796
rect 11612 47676 11664 47728
rect 14924 47719 14976 47728
rect 14924 47685 14933 47719
rect 14933 47685 14967 47719
rect 14967 47685 14976 47719
rect 14924 47676 14976 47685
rect 12900 47608 12952 47660
rect 10416 47540 10468 47592
rect 8024 47515 8076 47524
rect 8024 47481 8042 47515
rect 8042 47481 8076 47515
rect 8024 47472 8076 47481
rect 10968 47472 11020 47524
rect 6920 47447 6972 47456
rect 6920 47413 6929 47447
rect 6929 47413 6963 47447
rect 6963 47413 6972 47447
rect 6920 47404 6972 47413
rect 10876 47404 10928 47456
rect 12808 47447 12860 47456
rect 12808 47413 12817 47447
rect 12817 47413 12851 47447
rect 12851 47413 12860 47447
rect 12808 47404 12860 47413
rect 13084 47540 13136 47592
rect 13728 47540 13780 47592
rect 14372 47540 14424 47592
rect 18052 47540 18104 47592
rect 21916 47540 21968 47592
rect 13820 47472 13872 47524
rect 15752 47472 15804 47524
rect 17868 47472 17920 47524
rect 20996 47472 21048 47524
rect 22560 47472 22612 47524
rect 13544 47404 13596 47456
rect 16120 47404 16172 47456
rect 17684 47404 17736 47456
rect 19708 47447 19760 47456
rect 19708 47413 19717 47447
rect 19717 47413 19751 47447
rect 19751 47413 19760 47447
rect 19708 47404 19760 47413
rect 22376 47404 22428 47456
rect 24492 47404 24544 47456
rect 11253 47302 11305 47354
rect 11317 47302 11369 47354
rect 11381 47302 11433 47354
rect 11445 47302 11497 47354
rect 11509 47302 11561 47354
rect 21557 47302 21609 47354
rect 21621 47302 21673 47354
rect 21685 47302 21737 47354
rect 21749 47302 21801 47354
rect 21813 47302 21865 47354
rect 15384 47243 15436 47252
rect 15384 47209 15393 47243
rect 15393 47209 15427 47243
rect 15427 47209 15436 47243
rect 15384 47200 15436 47209
rect 15844 47200 15896 47252
rect 22560 47243 22612 47252
rect 22560 47209 22569 47243
rect 22569 47209 22603 47243
rect 22603 47209 22612 47243
rect 22560 47200 22612 47209
rect 24768 47243 24820 47252
rect 24768 47209 24777 47243
rect 24777 47209 24811 47243
rect 24811 47209 24820 47243
rect 24768 47200 24820 47209
rect 31300 47243 31352 47252
rect 31300 47209 31309 47243
rect 31309 47209 31343 47243
rect 31343 47209 31352 47243
rect 31300 47200 31352 47209
rect 7748 47107 7800 47116
rect 7748 47073 7757 47107
rect 7757 47073 7791 47107
rect 7791 47073 7800 47107
rect 7748 47064 7800 47073
rect 7840 47064 7892 47116
rect 10416 47132 10468 47184
rect 12808 47132 12860 47184
rect 9864 47107 9916 47116
rect 9864 47073 9898 47107
rect 9898 47073 9916 47107
rect 9864 47064 9916 47073
rect 13360 47064 13412 47116
rect 16120 47107 16172 47116
rect 16120 47073 16129 47107
rect 16129 47073 16163 47107
rect 16163 47073 16172 47107
rect 16120 47064 16172 47073
rect 17408 47064 17460 47116
rect 18052 47107 18104 47116
rect 18052 47073 18061 47107
rect 18061 47073 18095 47107
rect 18095 47073 18104 47107
rect 20720 47132 20772 47184
rect 23848 47132 23900 47184
rect 18052 47064 18104 47073
rect 18788 47064 18840 47116
rect 19708 47064 19760 47116
rect 20168 47064 20220 47116
rect 21456 47064 21508 47116
rect 22008 47107 22060 47116
rect 22008 47073 22017 47107
rect 22017 47073 22051 47107
rect 22051 47073 22060 47107
rect 22008 47064 22060 47073
rect 22376 47107 22428 47116
rect 22376 47073 22385 47107
rect 22385 47073 22419 47107
rect 22419 47073 22428 47107
rect 22376 47064 22428 47073
rect 30656 47064 30708 47116
rect 12164 47039 12216 47048
rect 12164 47005 12173 47039
rect 12173 47005 12207 47039
rect 12207 47005 12216 47039
rect 12164 46996 12216 47005
rect 11612 46971 11664 46980
rect 11612 46937 11621 46971
rect 11621 46937 11655 46971
rect 11655 46937 11664 46971
rect 11612 46928 11664 46937
rect 9220 46860 9272 46912
rect 10876 46860 10928 46912
rect 13544 46903 13596 46912
rect 13544 46869 13553 46903
rect 13553 46869 13587 46903
rect 13587 46869 13596 46903
rect 13544 46860 13596 46869
rect 21272 46996 21324 47048
rect 22560 46996 22612 47048
rect 16028 46971 16080 46980
rect 16028 46937 16037 46971
rect 16037 46937 16071 46971
rect 16071 46937 16080 46971
rect 16028 46928 16080 46937
rect 20628 46971 20680 46980
rect 20628 46937 20637 46971
rect 20637 46937 20671 46971
rect 20671 46937 20680 46971
rect 20628 46928 20680 46937
rect 21364 46928 21416 46980
rect 21916 46928 21968 46980
rect 14372 46860 14424 46912
rect 17316 46860 17368 46912
rect 18972 46860 19024 46912
rect 21088 46860 21140 46912
rect 30656 46903 30708 46912
rect 30656 46869 30665 46903
rect 30665 46869 30699 46903
rect 30699 46869 30708 46903
rect 30656 46860 30708 46869
rect 6102 46758 6154 46810
rect 6166 46758 6218 46810
rect 6230 46758 6282 46810
rect 6294 46758 6346 46810
rect 6358 46758 6410 46810
rect 16405 46758 16457 46810
rect 16469 46758 16521 46810
rect 16533 46758 16585 46810
rect 16597 46758 16649 46810
rect 16661 46758 16713 46810
rect 26709 46758 26761 46810
rect 26773 46758 26825 46810
rect 26837 46758 26889 46810
rect 26901 46758 26953 46810
rect 26965 46758 27017 46810
rect 7840 46656 7892 46708
rect 13820 46656 13872 46708
rect 17868 46699 17920 46708
rect 17868 46665 17877 46699
rect 17877 46665 17911 46699
rect 17911 46665 17920 46699
rect 17868 46656 17920 46665
rect 18328 46699 18380 46708
rect 18328 46665 18337 46699
rect 18337 46665 18371 46699
rect 18371 46665 18380 46699
rect 18328 46656 18380 46665
rect 6920 46520 6972 46572
rect 23756 46588 23808 46640
rect 7288 46452 7340 46504
rect 7840 46495 7892 46504
rect 7840 46461 7849 46495
rect 7849 46461 7883 46495
rect 7883 46461 7892 46495
rect 7840 46452 7892 46461
rect 9220 46520 9272 46572
rect 9496 46563 9548 46572
rect 9496 46529 9505 46563
rect 9505 46529 9539 46563
rect 9539 46529 9548 46563
rect 9496 46520 9548 46529
rect 13544 46520 13596 46572
rect 7564 46384 7616 46436
rect 9036 46452 9088 46504
rect 9404 46495 9456 46504
rect 9404 46461 9413 46495
rect 9413 46461 9447 46495
rect 9447 46461 9456 46495
rect 9680 46495 9732 46504
rect 9404 46452 9456 46461
rect 9680 46461 9689 46495
rect 9689 46461 9723 46495
rect 9723 46461 9732 46495
rect 9680 46452 9732 46461
rect 10416 46452 10468 46504
rect 12164 46495 12216 46504
rect 12164 46461 12173 46495
rect 12173 46461 12207 46495
rect 12207 46461 12216 46495
rect 12164 46452 12216 46461
rect 12808 46452 12860 46504
rect 14372 46495 14424 46504
rect 14372 46461 14381 46495
rect 14381 46461 14415 46495
rect 14415 46461 14424 46495
rect 14372 46452 14424 46461
rect 21916 46520 21968 46572
rect 23480 46520 23532 46572
rect 16672 46452 16724 46504
rect 17132 46495 17184 46504
rect 17132 46461 17141 46495
rect 17141 46461 17175 46495
rect 17175 46461 17184 46495
rect 17132 46452 17184 46461
rect 17316 46495 17368 46504
rect 17316 46461 17325 46495
rect 17325 46461 17359 46495
rect 17359 46461 17368 46495
rect 17316 46452 17368 46461
rect 17684 46495 17736 46504
rect 9772 46384 9824 46436
rect 14096 46384 14148 46436
rect 14648 46427 14700 46436
rect 14648 46393 14682 46427
rect 14682 46393 14700 46427
rect 14648 46384 14700 46393
rect 11704 46359 11756 46368
rect 11704 46325 11713 46359
rect 11713 46325 11747 46359
rect 11747 46325 11756 46359
rect 11704 46316 11756 46325
rect 12624 46316 12676 46368
rect 13728 46316 13780 46368
rect 15108 46316 15160 46368
rect 16304 46359 16356 46368
rect 16304 46325 16313 46359
rect 16313 46325 16347 46359
rect 16347 46325 16356 46359
rect 16304 46316 16356 46325
rect 17684 46461 17693 46495
rect 17693 46461 17727 46495
rect 17727 46461 17736 46495
rect 17684 46452 17736 46461
rect 18328 46452 18380 46504
rect 24216 46452 24268 46504
rect 17592 46384 17644 46436
rect 19616 46384 19668 46436
rect 20076 46384 20128 46436
rect 20812 46384 20864 46436
rect 23112 46384 23164 46436
rect 24492 46452 24544 46504
rect 17500 46316 17552 46368
rect 19984 46316 20036 46368
rect 20720 46316 20772 46368
rect 21916 46316 21968 46368
rect 22008 46316 22060 46368
rect 23664 46316 23716 46368
rect 24308 46316 24360 46368
rect 25136 46359 25188 46368
rect 25136 46325 25145 46359
rect 25145 46325 25179 46359
rect 25179 46325 25188 46359
rect 25136 46316 25188 46325
rect 25688 46359 25740 46368
rect 25688 46325 25697 46359
rect 25697 46325 25731 46359
rect 25731 46325 25740 46359
rect 25688 46316 25740 46325
rect 11253 46214 11305 46266
rect 11317 46214 11369 46266
rect 11381 46214 11433 46266
rect 11445 46214 11497 46266
rect 11509 46214 11561 46266
rect 21557 46214 21609 46266
rect 21621 46214 21673 46266
rect 21685 46214 21737 46266
rect 21749 46214 21801 46266
rect 21813 46214 21865 46266
rect 1400 46019 1452 46028
rect 1400 45985 1431 46019
rect 1431 45985 1452 46019
rect 1400 45976 1452 45985
rect 7748 46044 7800 46096
rect 7196 45976 7248 46028
rect 9036 46019 9088 46028
rect 7472 45840 7524 45892
rect 9036 45985 9045 46019
rect 9045 45985 9079 46019
rect 9079 45985 9088 46019
rect 9036 45976 9088 45985
rect 9220 46019 9272 46028
rect 9220 45985 9229 46019
rect 9229 45985 9263 46019
rect 9263 45985 9272 46019
rect 9220 45976 9272 45985
rect 9404 46112 9456 46164
rect 9864 46112 9916 46164
rect 10968 46155 11020 46164
rect 10968 46121 10977 46155
rect 10977 46121 11011 46155
rect 11011 46121 11020 46155
rect 10968 46112 11020 46121
rect 13360 46155 13412 46164
rect 13360 46121 13369 46155
rect 13369 46121 13403 46155
rect 13403 46121 13412 46155
rect 13360 46112 13412 46121
rect 14648 46112 14700 46164
rect 15752 46155 15804 46164
rect 15752 46121 15761 46155
rect 15761 46121 15795 46155
rect 15795 46121 15804 46155
rect 15752 46112 15804 46121
rect 17408 46155 17460 46164
rect 17408 46121 17417 46155
rect 17417 46121 17451 46155
rect 17451 46121 17460 46155
rect 17408 46112 17460 46121
rect 18788 46155 18840 46164
rect 18788 46121 18797 46155
rect 18797 46121 18831 46155
rect 18831 46121 18840 46155
rect 18788 46112 18840 46121
rect 20812 46112 20864 46164
rect 9680 46044 9732 46096
rect 9496 45976 9548 46028
rect 9772 45976 9824 46028
rect 10232 46019 10284 46028
rect 10232 45985 10241 46019
rect 10241 45985 10275 46019
rect 10275 45985 10284 46019
rect 10232 45976 10284 45985
rect 10784 46019 10836 46028
rect 10784 45985 10793 46019
rect 10793 45985 10827 46019
rect 10827 45985 10836 46019
rect 10784 45976 10836 45985
rect 11704 46019 11756 46028
rect 11704 45985 11723 46019
rect 11723 45985 11756 46019
rect 11704 45976 11756 45985
rect 12624 46019 12676 46028
rect 12624 45985 12633 46019
rect 12633 45985 12667 46019
rect 12667 45985 12676 46019
rect 12624 45976 12676 45985
rect 12808 46019 12860 46028
rect 12808 45985 12817 46019
rect 12817 45985 12851 46019
rect 12851 45985 12860 46019
rect 12808 45976 12860 45985
rect 13728 45976 13780 46028
rect 15384 46044 15436 46096
rect 16120 46044 16172 46096
rect 4988 45772 5040 45824
rect 8392 45772 8444 45824
rect 10508 45951 10560 45960
rect 10508 45917 10517 45951
rect 10517 45917 10551 45951
rect 10551 45917 10560 45951
rect 10508 45908 10560 45917
rect 10600 45951 10652 45960
rect 10600 45917 10609 45951
rect 10609 45917 10643 45951
rect 10643 45917 10652 45951
rect 12900 45951 12952 45960
rect 10600 45908 10652 45917
rect 12900 45917 12909 45951
rect 12909 45917 12943 45951
rect 12943 45917 12952 45951
rect 12900 45908 12952 45917
rect 12992 45951 13044 45960
rect 12992 45917 13001 45951
rect 13001 45917 13035 45951
rect 13035 45917 13044 45951
rect 12992 45908 13044 45917
rect 9772 45840 9824 45892
rect 10876 45840 10928 45892
rect 10232 45772 10284 45824
rect 10968 45772 11020 45824
rect 13084 45840 13136 45892
rect 13728 45840 13780 45892
rect 14188 45951 14240 45960
rect 14188 45917 14197 45951
rect 14197 45917 14231 45951
rect 14231 45917 14240 45951
rect 14832 45976 14884 46028
rect 15108 45976 15160 46028
rect 16672 46019 16724 46028
rect 16672 45985 16681 46019
rect 16681 45985 16715 46019
rect 16715 45985 16724 46019
rect 16672 45976 16724 45985
rect 17500 46044 17552 46096
rect 22008 46112 22060 46164
rect 17316 45976 17368 46028
rect 18972 46019 19024 46028
rect 18972 45985 18981 46019
rect 18981 45985 19015 46019
rect 19015 45985 19024 46019
rect 18972 45976 19024 45985
rect 19340 46019 19392 46028
rect 19340 45985 19349 46019
rect 19349 45985 19383 46019
rect 19383 45985 19392 46019
rect 19340 45976 19392 45985
rect 15292 45951 15344 45960
rect 14188 45908 14240 45917
rect 13912 45840 13964 45892
rect 15292 45917 15301 45951
rect 15301 45917 15335 45951
rect 15335 45917 15344 45951
rect 15292 45908 15344 45917
rect 17592 45908 17644 45960
rect 20168 46019 20220 46028
rect 20168 45985 20177 46019
rect 20177 45985 20211 46019
rect 20211 45985 20220 46019
rect 20168 45976 20220 45985
rect 20352 45951 20404 45960
rect 14188 45772 14240 45824
rect 18052 45772 18104 45824
rect 20352 45917 20361 45951
rect 20361 45917 20395 45951
rect 20395 45917 20404 45951
rect 20352 45908 20404 45917
rect 20812 45976 20864 46028
rect 22284 46044 22336 46096
rect 25136 46044 25188 46096
rect 22100 46019 22152 46028
rect 22100 45985 22109 46019
rect 22109 45985 22143 46019
rect 22143 45985 22152 46019
rect 22376 46019 22428 46028
rect 22100 45976 22152 45985
rect 22376 45985 22385 46019
rect 22385 45985 22419 46019
rect 22419 45985 22428 46019
rect 22376 45976 22428 45985
rect 24032 45976 24084 46028
rect 24124 45976 24176 46028
rect 30656 46019 30708 46028
rect 30656 45985 30665 46019
rect 30665 45985 30699 46019
rect 30699 45985 30708 46019
rect 30656 45976 30708 45985
rect 31576 45976 31628 46028
rect 21272 45908 21324 45960
rect 21548 45908 21600 45960
rect 21916 45908 21968 45960
rect 26148 45951 26200 45960
rect 26148 45917 26157 45951
rect 26157 45917 26191 45951
rect 26191 45917 26200 45951
rect 26148 45908 26200 45917
rect 21456 45840 21508 45892
rect 24216 45840 24268 45892
rect 20352 45772 20404 45824
rect 20904 45772 20956 45824
rect 21088 45772 21140 45824
rect 21640 45772 21692 45824
rect 21916 45772 21968 45824
rect 24308 45815 24360 45824
rect 24308 45781 24317 45815
rect 24317 45781 24351 45815
rect 24351 45781 24360 45815
rect 24308 45772 24360 45781
rect 24400 45772 24452 45824
rect 26240 45772 26292 45824
rect 6102 45670 6154 45722
rect 6166 45670 6218 45722
rect 6230 45670 6282 45722
rect 6294 45670 6346 45722
rect 6358 45670 6410 45722
rect 16405 45670 16457 45722
rect 16469 45670 16521 45722
rect 16533 45670 16585 45722
rect 16597 45670 16649 45722
rect 16661 45670 16713 45722
rect 26709 45670 26761 45722
rect 26773 45670 26825 45722
rect 26837 45670 26889 45722
rect 26901 45670 26953 45722
rect 26965 45670 27017 45722
rect 1400 45611 1452 45620
rect 1400 45577 1409 45611
rect 1409 45577 1443 45611
rect 1443 45577 1452 45611
rect 1400 45568 1452 45577
rect 9496 45568 9548 45620
rect 10600 45568 10652 45620
rect 13728 45568 13780 45620
rect 8024 45543 8076 45552
rect 8024 45509 8033 45543
rect 8033 45509 8067 45543
rect 8067 45509 8076 45543
rect 8024 45500 8076 45509
rect 9864 45500 9916 45552
rect 11612 45500 11664 45552
rect 14188 45500 14240 45552
rect 14280 45500 14332 45552
rect 7564 45475 7616 45484
rect 7564 45441 7573 45475
rect 7573 45441 7607 45475
rect 7607 45441 7616 45475
rect 7564 45432 7616 45441
rect 12900 45432 12952 45484
rect 14096 45475 14148 45484
rect 14096 45441 14105 45475
rect 14105 45441 14139 45475
rect 14139 45441 14148 45475
rect 14096 45432 14148 45441
rect 15292 45568 15344 45620
rect 19616 45568 19668 45620
rect 16212 45500 16264 45552
rect 20996 45500 21048 45552
rect 21456 45500 21508 45552
rect 22284 45500 22336 45552
rect 23480 45500 23532 45552
rect 15752 45432 15804 45484
rect 6920 45364 6972 45416
rect 7288 45407 7340 45416
rect 7288 45373 7297 45407
rect 7297 45373 7331 45407
rect 7331 45373 7340 45407
rect 7288 45364 7340 45373
rect 7472 45407 7524 45416
rect 7472 45373 7485 45407
rect 7485 45373 7519 45407
rect 7519 45373 7524 45407
rect 7472 45364 7524 45373
rect 7840 45407 7892 45416
rect 7380 45296 7432 45348
rect 7840 45373 7849 45407
rect 7849 45373 7883 45407
rect 7883 45373 7892 45407
rect 7840 45364 7892 45373
rect 9220 45364 9272 45416
rect 10876 45407 10928 45416
rect 10876 45373 10885 45407
rect 10885 45373 10919 45407
rect 10919 45373 10928 45407
rect 10876 45364 10928 45373
rect 11980 45364 12032 45416
rect 12532 45407 12584 45416
rect 9496 45339 9548 45348
rect 9496 45305 9505 45339
rect 9505 45305 9539 45339
rect 9539 45305 9548 45339
rect 9496 45296 9548 45305
rect 12532 45373 12541 45407
rect 12541 45373 12575 45407
rect 12575 45373 12584 45407
rect 12532 45364 12584 45373
rect 13820 45364 13872 45416
rect 13912 45296 13964 45348
rect 14648 45407 14700 45416
rect 14648 45373 14657 45407
rect 14657 45373 14691 45407
rect 14691 45373 14700 45407
rect 14648 45364 14700 45373
rect 14832 45407 14884 45416
rect 14832 45373 14841 45407
rect 14841 45373 14875 45407
rect 14875 45373 14884 45407
rect 20904 45432 20956 45484
rect 14832 45364 14884 45373
rect 16672 45296 16724 45348
rect 8024 45228 8076 45280
rect 9772 45228 9824 45280
rect 10784 45271 10836 45280
rect 10784 45237 10793 45271
rect 10793 45237 10827 45271
rect 10827 45237 10836 45271
rect 10784 45228 10836 45237
rect 15108 45228 15160 45280
rect 15568 45228 15620 45280
rect 16856 45228 16908 45280
rect 20720 45364 20772 45416
rect 17960 45296 18012 45348
rect 21180 45296 21232 45348
rect 18512 45228 18564 45280
rect 18696 45271 18748 45280
rect 18696 45237 18705 45271
rect 18705 45237 18739 45271
rect 18739 45237 18748 45271
rect 18696 45228 18748 45237
rect 19340 45228 19392 45280
rect 19800 45228 19852 45280
rect 20168 45228 20220 45280
rect 21548 45373 21557 45394
rect 21557 45373 21591 45394
rect 21591 45373 21600 45394
rect 21548 45342 21600 45373
rect 21640 45407 21692 45416
rect 21640 45373 21649 45407
rect 21649 45373 21683 45407
rect 21683 45373 21692 45407
rect 21640 45364 21692 45373
rect 23112 45407 23164 45416
rect 23112 45373 23121 45407
rect 23121 45373 23155 45407
rect 23155 45373 23164 45407
rect 23112 45364 23164 45373
rect 23296 45409 23348 45416
rect 23296 45375 23305 45409
rect 23305 45375 23339 45409
rect 23339 45375 23348 45409
rect 23296 45364 23348 45375
rect 23756 45432 23808 45484
rect 26148 45568 26200 45620
rect 26240 45611 26292 45620
rect 26240 45577 26249 45611
rect 26249 45577 26283 45611
rect 26283 45577 26292 45611
rect 26240 45568 26292 45577
rect 26148 45432 26200 45484
rect 27620 45432 27672 45484
rect 27528 45364 27580 45416
rect 22192 45228 22244 45280
rect 23940 45228 23992 45280
rect 26056 45228 26108 45280
rect 11253 45126 11305 45178
rect 11317 45126 11369 45178
rect 11381 45126 11433 45178
rect 11445 45126 11497 45178
rect 11509 45126 11561 45178
rect 21557 45126 21609 45178
rect 21621 45126 21673 45178
rect 21685 45126 21737 45178
rect 21749 45126 21801 45178
rect 21813 45126 21865 45178
rect 7196 45067 7248 45076
rect 7196 45033 7205 45067
rect 7205 45033 7239 45067
rect 7239 45033 7248 45067
rect 7196 45024 7248 45033
rect 10692 45024 10744 45076
rect 7288 44956 7340 45008
rect 7564 44956 7616 45008
rect 7472 44888 7524 44940
rect 7748 44931 7800 44940
rect 7748 44897 7757 44931
rect 7757 44897 7791 44931
rect 7791 44897 7800 44931
rect 7748 44888 7800 44897
rect 11152 44956 11204 45008
rect 10232 44931 10284 44940
rect 10232 44897 10241 44931
rect 10241 44897 10275 44931
rect 10275 44897 10284 44931
rect 10232 44888 10284 44897
rect 10692 44888 10744 44940
rect 10876 44888 10928 44940
rect 13636 45024 13688 45076
rect 14832 45024 14884 45076
rect 7196 44820 7248 44872
rect 7656 44863 7708 44872
rect 7656 44829 7665 44863
rect 7665 44829 7699 44863
rect 7699 44829 7708 44863
rect 7656 44820 7708 44829
rect 9312 44820 9364 44872
rect 9956 44820 10008 44872
rect 10508 44863 10560 44872
rect 10508 44829 10517 44863
rect 10517 44829 10551 44863
rect 10551 44829 10560 44863
rect 10508 44820 10560 44829
rect 10600 44863 10652 44872
rect 10600 44829 10609 44863
rect 10609 44829 10643 44863
rect 10643 44829 10652 44863
rect 13636 44888 13688 44940
rect 14648 44931 14700 44940
rect 14648 44897 14657 44931
rect 14657 44897 14691 44931
rect 14691 44897 14700 44931
rect 14648 44888 14700 44897
rect 15752 45024 15804 45076
rect 17040 45024 17092 45076
rect 17960 45067 18012 45076
rect 15108 44956 15160 45008
rect 15476 44931 15528 44940
rect 10600 44820 10652 44829
rect 12624 44820 12676 44872
rect 13452 44820 13504 44872
rect 15476 44897 15485 44931
rect 15485 44897 15519 44931
rect 15519 44897 15528 44931
rect 15476 44888 15528 44897
rect 15752 44931 15804 44940
rect 15752 44897 15761 44931
rect 15761 44897 15795 44931
rect 15795 44897 15804 44931
rect 15752 44888 15804 44897
rect 15936 44888 15988 44940
rect 17132 44888 17184 44940
rect 17684 44888 17736 44940
rect 17960 45033 17969 45067
rect 17969 45033 18003 45067
rect 18003 45033 18012 45067
rect 17960 45024 18012 45033
rect 18512 45067 18564 45076
rect 18512 45033 18521 45067
rect 18521 45033 18555 45067
rect 18555 45033 18564 45067
rect 18512 45024 18564 45033
rect 21180 45024 21232 45076
rect 21272 44956 21324 45008
rect 15844 44820 15896 44872
rect 17500 44863 17552 44872
rect 17500 44829 17509 44863
rect 17509 44829 17543 44863
rect 17543 44829 17552 44863
rect 17500 44820 17552 44829
rect 17592 44863 17644 44872
rect 17592 44829 17601 44863
rect 17601 44829 17635 44863
rect 17635 44829 17644 44863
rect 17868 44888 17920 44940
rect 19800 44931 19852 44940
rect 17592 44820 17644 44829
rect 18696 44820 18748 44872
rect 19800 44897 19809 44931
rect 19809 44897 19843 44931
rect 19843 44897 19852 44931
rect 19800 44888 19852 44897
rect 22100 44956 22152 45008
rect 23388 45024 23440 45076
rect 23480 44956 23532 45008
rect 24124 45067 24176 45076
rect 24124 45033 24133 45067
rect 24133 45033 24167 45067
rect 24167 45033 24176 45067
rect 24124 45024 24176 45033
rect 12348 44752 12400 44804
rect 16120 44752 16172 44804
rect 16672 44752 16724 44804
rect 21088 44820 21140 44872
rect 21456 44888 21508 44940
rect 22008 44931 22060 44940
rect 22008 44897 22017 44931
rect 22017 44897 22051 44931
rect 22051 44897 22060 44931
rect 22008 44888 22060 44897
rect 22192 44931 22244 44940
rect 22192 44897 22201 44931
rect 22201 44897 22235 44931
rect 22235 44897 22244 44931
rect 22192 44888 22244 44897
rect 23112 44888 23164 44940
rect 24400 44888 24452 44940
rect 24492 44888 24544 44940
rect 25688 44888 25740 44940
rect 26424 44888 26476 44940
rect 23756 44863 23808 44872
rect 23756 44829 23765 44863
rect 23765 44829 23799 44863
rect 23799 44829 23808 44863
rect 23756 44820 23808 44829
rect 24216 44820 24268 44872
rect 24308 44752 24360 44804
rect 24768 44752 24820 44804
rect 7380 44684 7432 44736
rect 10140 44684 10192 44736
rect 15936 44727 15988 44736
rect 15936 44693 15945 44727
rect 15945 44693 15979 44727
rect 15979 44693 15988 44727
rect 15936 44684 15988 44693
rect 16212 44684 16264 44736
rect 16948 44684 17000 44736
rect 22376 44684 22428 44736
rect 24032 44684 24084 44736
rect 24860 44684 24912 44736
rect 26332 44684 26384 44736
rect 27620 44684 27672 44736
rect 30932 44727 30984 44736
rect 30932 44693 30941 44727
rect 30941 44693 30975 44727
rect 30975 44693 30984 44727
rect 30932 44684 30984 44693
rect 6102 44582 6154 44634
rect 6166 44582 6218 44634
rect 6230 44582 6282 44634
rect 6294 44582 6346 44634
rect 6358 44582 6410 44634
rect 16405 44582 16457 44634
rect 16469 44582 16521 44634
rect 16533 44582 16585 44634
rect 16597 44582 16649 44634
rect 16661 44582 16713 44634
rect 26709 44582 26761 44634
rect 26773 44582 26825 44634
rect 26837 44582 26889 44634
rect 26901 44582 26953 44634
rect 26965 44582 27017 44634
rect 2688 44480 2740 44532
rect 7012 44412 7064 44464
rect 7748 44412 7800 44464
rect 9496 44412 9548 44464
rect 12072 44412 12124 44464
rect 10600 44344 10652 44396
rect 14280 44344 14332 44396
rect 14464 44344 14516 44396
rect 5816 44319 5868 44328
rect 5816 44285 5825 44319
rect 5825 44285 5859 44319
rect 5859 44285 5868 44319
rect 5816 44276 5868 44285
rect 8024 44319 8076 44328
rect 8024 44285 8033 44319
rect 8033 44285 8067 44319
rect 8067 44285 8076 44319
rect 8024 44276 8076 44285
rect 8392 44319 8444 44328
rect 1860 44251 1912 44260
rect 1860 44217 1869 44251
rect 1869 44217 1903 44251
rect 1903 44217 1912 44251
rect 1860 44208 1912 44217
rect 6828 44208 6880 44260
rect 7932 44208 7984 44260
rect 8392 44285 8401 44319
rect 8401 44285 8435 44319
rect 8435 44285 8444 44319
rect 8392 44276 8444 44285
rect 10508 44276 10560 44328
rect 9864 44251 9916 44260
rect 9864 44217 9873 44251
rect 9873 44217 9907 44251
rect 9907 44217 9916 44251
rect 9864 44208 9916 44217
rect 11612 44251 11664 44260
rect 11612 44217 11621 44251
rect 11621 44217 11655 44251
rect 11655 44217 11664 44251
rect 12164 44276 12216 44328
rect 12348 44319 12400 44328
rect 12348 44285 12382 44319
rect 12382 44285 12400 44319
rect 12348 44276 12400 44285
rect 15476 44319 15528 44328
rect 15476 44285 15485 44319
rect 15485 44285 15519 44319
rect 15519 44285 15528 44319
rect 15476 44276 15528 44285
rect 18052 44480 18104 44532
rect 22560 44480 22612 44532
rect 23756 44480 23808 44532
rect 24124 44480 24176 44532
rect 16212 44344 16264 44396
rect 15752 44319 15804 44328
rect 15752 44285 15761 44319
rect 15761 44285 15795 44319
rect 15795 44285 15804 44319
rect 16028 44319 16080 44328
rect 15752 44276 15804 44285
rect 16028 44285 16037 44319
rect 16037 44285 16071 44319
rect 16071 44285 16080 44319
rect 16028 44276 16080 44285
rect 17132 44412 17184 44464
rect 17040 44319 17092 44328
rect 17040 44285 17049 44319
rect 17049 44285 17083 44319
rect 17083 44285 17092 44319
rect 17040 44276 17092 44285
rect 17592 44344 17644 44396
rect 18420 44344 18472 44396
rect 21456 44412 21508 44464
rect 22836 44412 22888 44464
rect 24216 44412 24268 44464
rect 24492 44455 24544 44464
rect 24492 44421 24501 44455
rect 24501 44421 24535 44455
rect 24535 44421 24544 44455
rect 24492 44412 24544 44421
rect 27068 44412 27120 44464
rect 27528 44412 27580 44464
rect 29368 44412 29420 44464
rect 22100 44344 22152 44396
rect 22192 44344 22244 44396
rect 11612 44208 11664 44217
rect 9128 44140 9180 44192
rect 9220 44183 9272 44192
rect 9220 44149 9229 44183
rect 9229 44149 9263 44183
rect 9263 44149 9272 44183
rect 9220 44140 9272 44149
rect 13912 44208 13964 44260
rect 16948 44208 17000 44260
rect 17960 44276 18012 44328
rect 17316 44208 17368 44260
rect 12256 44140 12308 44192
rect 16396 44140 16448 44192
rect 17224 44140 17276 44192
rect 17592 44183 17644 44192
rect 17592 44149 17601 44183
rect 17601 44149 17635 44183
rect 17635 44149 17644 44183
rect 17592 44140 17644 44149
rect 17684 44140 17736 44192
rect 21272 44276 21324 44328
rect 22008 44276 22060 44328
rect 22744 44319 22796 44328
rect 22744 44285 22753 44319
rect 22753 44285 22787 44319
rect 22787 44285 22796 44319
rect 22744 44276 22796 44285
rect 23020 44319 23072 44328
rect 23020 44285 23029 44319
rect 23029 44285 23063 44319
rect 23063 44285 23072 44319
rect 23020 44276 23072 44285
rect 23664 44319 23716 44328
rect 23664 44285 23673 44319
rect 23673 44285 23707 44319
rect 23707 44285 23716 44319
rect 23664 44276 23716 44285
rect 24216 44208 24268 44260
rect 19432 44140 19484 44192
rect 20628 44140 20680 44192
rect 20812 44140 20864 44192
rect 21456 44140 21508 44192
rect 22284 44183 22336 44192
rect 22284 44149 22293 44183
rect 22293 44149 22327 44183
rect 22327 44149 22336 44183
rect 22284 44140 22336 44149
rect 22376 44140 22428 44192
rect 24584 44276 24636 44328
rect 26608 44208 26660 44260
rect 27620 44276 27672 44328
rect 31116 44319 31168 44328
rect 31116 44285 31125 44319
rect 31125 44285 31159 44319
rect 31159 44285 31168 44319
rect 31116 44276 31168 44285
rect 27344 44208 27396 44260
rect 25320 44140 25372 44192
rect 25872 44140 25924 44192
rect 26240 44140 26292 44192
rect 30656 44183 30708 44192
rect 30656 44149 30665 44183
rect 30665 44149 30699 44183
rect 30699 44149 30708 44183
rect 30656 44140 30708 44149
rect 11253 44038 11305 44090
rect 11317 44038 11369 44090
rect 11381 44038 11433 44090
rect 11445 44038 11497 44090
rect 11509 44038 11561 44090
rect 21557 44038 21609 44090
rect 21621 44038 21673 44090
rect 21685 44038 21737 44090
rect 21749 44038 21801 44090
rect 21813 44038 21865 44090
rect 6828 43979 6880 43988
rect 6828 43945 6837 43979
rect 6837 43945 6871 43979
rect 6871 43945 6880 43979
rect 6828 43936 6880 43945
rect 14648 43936 14700 43988
rect 17224 43936 17276 43988
rect 1860 43868 1912 43920
rect 12256 43868 12308 43920
rect 7012 43843 7064 43852
rect 7012 43809 7021 43843
rect 7021 43809 7055 43843
rect 7055 43809 7064 43843
rect 7012 43800 7064 43809
rect 7472 43800 7524 43852
rect 7564 43843 7616 43852
rect 7564 43809 7573 43843
rect 7573 43809 7607 43843
rect 7607 43809 7616 43843
rect 7564 43800 7616 43809
rect 9496 43800 9548 43852
rect 10876 43843 10928 43852
rect 10876 43809 10885 43843
rect 10885 43809 10919 43843
rect 10919 43809 10928 43843
rect 10876 43800 10928 43809
rect 14556 43868 14608 43920
rect 15752 43868 15804 43920
rect 14924 43843 14976 43852
rect 7196 43775 7248 43784
rect 7196 43741 7205 43775
rect 7205 43741 7239 43775
rect 7239 43741 7248 43775
rect 7196 43732 7248 43741
rect 7288 43775 7340 43784
rect 7288 43741 7297 43775
rect 7297 43741 7331 43775
rect 7331 43741 7340 43775
rect 8576 43775 8628 43784
rect 7288 43732 7340 43741
rect 8576 43741 8585 43775
rect 8585 43741 8619 43775
rect 8619 43741 8628 43775
rect 8576 43732 8628 43741
rect 9312 43775 9364 43784
rect 9312 43741 9321 43775
rect 9321 43741 9355 43775
rect 9355 43741 9364 43775
rect 9312 43732 9364 43741
rect 9956 43732 10008 43784
rect 11612 43732 11664 43784
rect 14464 43732 14516 43784
rect 14924 43809 14933 43843
rect 14933 43809 14967 43843
rect 14967 43809 14976 43843
rect 14924 43800 14976 43809
rect 15568 43843 15620 43852
rect 15568 43809 15577 43843
rect 15577 43809 15611 43843
rect 15611 43809 15620 43843
rect 15568 43800 15620 43809
rect 16304 43868 16356 43920
rect 17592 43868 17644 43920
rect 17960 43936 18012 43988
rect 20352 43936 20404 43988
rect 24216 43936 24268 43988
rect 26424 43979 26476 43988
rect 26424 43945 26433 43979
rect 26433 43945 26467 43979
rect 26467 43945 26476 43979
rect 26424 43936 26476 43945
rect 29368 43979 29420 43988
rect 29368 43945 29377 43979
rect 29377 43945 29411 43979
rect 29411 43945 29420 43979
rect 29368 43936 29420 43945
rect 16120 43843 16172 43852
rect 16120 43809 16129 43843
rect 16129 43809 16163 43843
rect 16163 43809 16172 43843
rect 16120 43800 16172 43809
rect 18972 43800 19024 43852
rect 20260 43800 20312 43852
rect 20536 43843 20588 43852
rect 20536 43809 20545 43843
rect 20545 43809 20579 43843
rect 20579 43809 20588 43843
rect 20536 43800 20588 43809
rect 21272 43800 21324 43852
rect 21364 43800 21416 43852
rect 22376 43843 22428 43852
rect 22376 43809 22385 43843
rect 22385 43809 22419 43843
rect 22419 43809 22428 43843
rect 22376 43800 22428 43809
rect 24860 43868 24912 43920
rect 23112 43800 23164 43852
rect 24400 43800 24452 43852
rect 25688 43843 25740 43852
rect 25688 43809 25697 43843
rect 25697 43809 25731 43843
rect 25731 43809 25740 43843
rect 25688 43800 25740 43809
rect 25872 43843 25924 43852
rect 25872 43809 25881 43843
rect 25881 43809 25915 43843
rect 25915 43809 25924 43843
rect 25872 43800 25924 43809
rect 26240 43843 26292 43852
rect 26240 43809 26249 43843
rect 26249 43809 26283 43843
rect 26283 43809 26292 43843
rect 26240 43800 26292 43809
rect 27160 43800 27212 43852
rect 15200 43732 15252 43784
rect 16212 43732 16264 43784
rect 15936 43664 15988 43716
rect 16396 43664 16448 43716
rect 2136 43639 2188 43648
rect 2136 43605 2145 43639
rect 2145 43605 2179 43639
rect 2179 43605 2188 43639
rect 2136 43596 2188 43605
rect 6736 43596 6788 43648
rect 10692 43596 10744 43648
rect 14464 43596 14516 43648
rect 15292 43596 15344 43648
rect 20444 43732 20496 43784
rect 21088 43732 21140 43784
rect 22192 43775 22244 43784
rect 22192 43741 22201 43775
rect 22201 43741 22235 43775
rect 22235 43741 22244 43775
rect 22192 43732 22244 43741
rect 22744 43732 22796 43784
rect 22928 43732 22980 43784
rect 22100 43664 22152 43716
rect 23296 43732 23348 43784
rect 26332 43732 26384 43784
rect 26148 43664 26200 43716
rect 18512 43596 18564 43648
rect 20168 43596 20220 43648
rect 23204 43596 23256 43648
rect 25228 43639 25280 43648
rect 25228 43605 25237 43639
rect 25237 43605 25271 43639
rect 25271 43605 25280 43639
rect 25228 43596 25280 43605
rect 27620 43596 27672 43648
rect 28724 43596 28776 43648
rect 31024 43639 31076 43648
rect 31024 43605 31033 43639
rect 31033 43605 31067 43639
rect 31067 43605 31076 43639
rect 31024 43596 31076 43605
rect 6102 43494 6154 43546
rect 6166 43494 6218 43546
rect 6230 43494 6282 43546
rect 6294 43494 6346 43546
rect 6358 43494 6410 43546
rect 16405 43494 16457 43546
rect 16469 43494 16521 43546
rect 16533 43494 16585 43546
rect 16597 43494 16649 43546
rect 16661 43494 16713 43546
rect 26709 43494 26761 43546
rect 26773 43494 26825 43546
rect 26837 43494 26889 43546
rect 26901 43494 26953 43546
rect 26965 43494 27017 43546
rect 5632 43392 5684 43444
rect 9312 43392 9364 43444
rect 10324 43324 10376 43376
rect 5816 43256 5868 43308
rect 9864 43256 9916 43308
rect 9956 43256 10008 43308
rect 15660 43392 15712 43444
rect 17776 43392 17828 43444
rect 24676 43392 24728 43444
rect 27160 43435 27212 43444
rect 27160 43401 27169 43435
rect 27169 43401 27203 43435
rect 27203 43401 27212 43435
rect 27160 43392 27212 43401
rect 30932 43392 30984 43444
rect 31116 43392 31168 43444
rect 21088 43324 21140 43376
rect 12532 43256 12584 43308
rect 14464 43256 14516 43308
rect 16948 43256 17000 43308
rect 17132 43256 17184 43308
rect 18420 43299 18472 43308
rect 18420 43265 18429 43299
rect 18429 43265 18463 43299
rect 18463 43265 18472 43299
rect 18420 43256 18472 43265
rect 1584 43052 1636 43104
rect 1768 43052 1820 43104
rect 2872 43052 2924 43104
rect 2964 43052 3016 43104
rect 4160 43052 4212 43104
rect 7288 43120 7340 43172
rect 9220 43188 9272 43240
rect 10232 43188 10284 43240
rect 10876 43231 10928 43240
rect 10876 43197 10885 43231
rect 10885 43197 10919 43231
rect 10919 43197 10928 43231
rect 10876 43188 10928 43197
rect 11060 43231 11112 43240
rect 11060 43197 11069 43231
rect 11069 43197 11103 43231
rect 11103 43197 11112 43231
rect 11060 43188 11112 43197
rect 11704 43120 11756 43172
rect 14372 43188 14424 43240
rect 15476 43231 15528 43240
rect 15476 43197 15485 43231
rect 15485 43197 15519 43231
rect 15519 43197 15528 43231
rect 15476 43188 15528 43197
rect 15568 43188 15620 43240
rect 19340 43188 19392 43240
rect 26148 43324 26200 43376
rect 20352 43188 20404 43240
rect 23480 43256 23532 43308
rect 23756 43256 23808 43308
rect 24400 43231 24452 43240
rect 24400 43197 24409 43231
rect 24409 43197 24443 43231
rect 24443 43197 24452 43231
rect 24400 43188 24452 43197
rect 26332 43256 26384 43308
rect 26424 43231 26476 43240
rect 12624 43120 12676 43172
rect 13268 43120 13320 43172
rect 15384 43120 15436 43172
rect 22468 43120 22520 43172
rect 5632 43052 5684 43104
rect 7472 43052 7524 43104
rect 9496 43052 9548 43104
rect 11796 43052 11848 43104
rect 15108 43052 15160 43104
rect 17408 43052 17460 43104
rect 22560 43052 22612 43104
rect 22652 43052 22704 43104
rect 23940 43052 23992 43104
rect 26424 43197 26433 43231
rect 26433 43197 26467 43231
rect 26467 43197 26476 43231
rect 26424 43188 26476 43197
rect 26240 43120 26292 43172
rect 26884 43188 26936 43240
rect 27620 43231 27672 43240
rect 27620 43197 27629 43231
rect 27629 43197 27663 43231
rect 27663 43197 27672 43231
rect 27620 43188 27672 43197
rect 28632 43188 28684 43240
rect 31116 43231 31168 43240
rect 31116 43197 31125 43231
rect 31125 43197 31159 43231
rect 31159 43197 31168 43231
rect 31116 43188 31168 43197
rect 26148 43052 26200 43104
rect 27712 43120 27764 43172
rect 28264 43120 28316 43172
rect 27160 43052 27212 43104
rect 29184 43052 29236 43104
rect 29552 43095 29604 43104
rect 29552 43061 29561 43095
rect 29561 43061 29595 43095
rect 29595 43061 29604 43095
rect 29552 43052 29604 43061
rect 11253 42950 11305 43002
rect 11317 42950 11369 43002
rect 11381 42950 11433 43002
rect 11445 42950 11497 43002
rect 11509 42950 11561 43002
rect 21557 42950 21609 43002
rect 21621 42950 21673 43002
rect 21685 42950 21737 43002
rect 21749 42950 21801 43002
rect 21813 42950 21865 43002
rect 9220 42848 9272 42900
rect 9404 42848 9456 42900
rect 9956 42848 10008 42900
rect 15384 42891 15436 42900
rect 11796 42823 11848 42832
rect 5724 42755 5776 42764
rect 5724 42721 5733 42755
rect 5733 42721 5767 42755
rect 5767 42721 5776 42755
rect 5724 42712 5776 42721
rect 7012 42712 7064 42764
rect 7564 42712 7616 42764
rect 8024 42712 8076 42764
rect 5172 42644 5224 42696
rect 7840 42644 7892 42696
rect 9128 42712 9180 42764
rect 9772 42755 9824 42764
rect 7196 42576 7248 42628
rect 9772 42721 9781 42755
rect 9781 42721 9815 42755
rect 9815 42721 9824 42755
rect 9772 42712 9824 42721
rect 10508 42712 10560 42764
rect 11796 42789 11830 42823
rect 11830 42789 11848 42823
rect 11796 42780 11848 42789
rect 10968 42755 11020 42764
rect 9588 42687 9640 42696
rect 9588 42653 9597 42687
rect 9597 42653 9631 42687
rect 9631 42653 9640 42687
rect 9588 42644 9640 42653
rect 10968 42721 10977 42755
rect 10977 42721 11011 42755
rect 11011 42721 11020 42755
rect 10968 42712 11020 42721
rect 11612 42712 11664 42764
rect 12992 42712 13044 42764
rect 14924 42780 14976 42832
rect 15384 42857 15393 42891
rect 15393 42857 15427 42891
rect 15427 42857 15436 42891
rect 15384 42848 15436 42857
rect 22560 42848 22612 42900
rect 23480 42848 23532 42900
rect 28264 42891 28316 42900
rect 20904 42780 20956 42832
rect 21364 42780 21416 42832
rect 14832 42755 14884 42764
rect 14832 42721 14841 42755
rect 14841 42721 14875 42755
rect 14875 42721 14884 42755
rect 14832 42712 14884 42721
rect 15200 42755 15252 42764
rect 15200 42721 15209 42755
rect 15209 42721 15243 42755
rect 15243 42721 15252 42755
rect 15200 42712 15252 42721
rect 16948 42755 17000 42764
rect 16948 42721 16957 42755
rect 16957 42721 16991 42755
rect 16991 42721 17000 42755
rect 16948 42712 17000 42721
rect 11152 42644 11204 42696
rect 13452 42644 13504 42696
rect 14464 42644 14516 42696
rect 15016 42687 15068 42696
rect 15016 42653 15025 42687
rect 15025 42653 15059 42687
rect 15059 42653 15068 42687
rect 17224 42687 17276 42696
rect 15016 42644 15068 42653
rect 17224 42653 17233 42687
rect 17233 42653 17267 42687
rect 17267 42653 17276 42687
rect 17224 42644 17276 42653
rect 17500 42755 17552 42764
rect 17500 42721 17509 42755
rect 17509 42721 17543 42755
rect 17543 42721 17552 42755
rect 17500 42712 17552 42721
rect 17684 42712 17736 42764
rect 18512 42712 18564 42764
rect 19248 42712 19300 42764
rect 19340 42712 19392 42764
rect 22468 42712 22520 42764
rect 23112 42755 23164 42764
rect 10784 42576 10836 42628
rect 15568 42576 15620 42628
rect 15844 42576 15896 42628
rect 17960 42644 18012 42696
rect 20996 42644 21048 42696
rect 17408 42576 17460 42628
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 2044 42551 2096 42560
rect 2044 42517 2053 42551
rect 2053 42517 2087 42551
rect 2087 42517 2096 42551
rect 2044 42508 2096 42517
rect 2320 42508 2372 42560
rect 3056 42551 3108 42560
rect 3056 42517 3065 42551
rect 3065 42517 3099 42551
rect 3099 42517 3108 42551
rect 3056 42508 3108 42517
rect 4160 42508 4212 42560
rect 4252 42508 4304 42560
rect 9128 42508 9180 42560
rect 10048 42508 10100 42560
rect 10140 42508 10192 42560
rect 10600 42508 10652 42560
rect 13268 42508 13320 42560
rect 16120 42508 16172 42560
rect 17316 42508 17368 42560
rect 17684 42551 17736 42560
rect 17684 42517 17693 42551
rect 17693 42517 17727 42551
rect 17727 42517 17736 42551
rect 17684 42508 17736 42517
rect 19524 42508 19576 42560
rect 20536 42576 20588 42628
rect 22652 42644 22704 42696
rect 23112 42721 23121 42755
rect 23121 42721 23155 42755
rect 23155 42721 23164 42755
rect 23756 42755 23808 42764
rect 23112 42712 23164 42721
rect 23756 42721 23765 42755
rect 23765 42721 23799 42755
rect 23799 42721 23808 42755
rect 23756 42712 23808 42721
rect 28264 42857 28273 42891
rect 28273 42857 28307 42891
rect 28307 42857 28316 42891
rect 28264 42848 28316 42857
rect 24216 42712 24268 42764
rect 25044 42712 25096 42764
rect 27620 42780 27672 42832
rect 26240 42755 26292 42764
rect 26240 42721 26249 42755
rect 26249 42721 26283 42755
rect 26283 42721 26292 42755
rect 26240 42712 26292 42721
rect 27712 42755 27764 42764
rect 27712 42721 27721 42755
rect 27721 42721 27755 42755
rect 27755 42721 27764 42755
rect 27712 42712 27764 42721
rect 28724 42755 28776 42764
rect 23572 42576 23624 42628
rect 24952 42687 25004 42696
rect 24952 42653 24961 42687
rect 24961 42653 24995 42687
rect 24995 42653 25004 42687
rect 24952 42644 25004 42653
rect 25688 42644 25740 42696
rect 26424 42644 26476 42696
rect 26976 42644 27028 42696
rect 27804 42687 27856 42696
rect 27804 42653 27813 42687
rect 27813 42653 27847 42687
rect 27847 42653 27856 42687
rect 27804 42644 27856 42653
rect 27896 42687 27948 42696
rect 27896 42653 27905 42687
rect 27905 42653 27939 42687
rect 27939 42653 27948 42687
rect 28724 42721 28733 42755
rect 28733 42721 28767 42755
rect 28767 42721 28776 42755
rect 28724 42712 28776 42721
rect 29368 42755 29420 42764
rect 29368 42721 29377 42755
rect 29377 42721 29411 42755
rect 29411 42721 29420 42755
rect 29368 42712 29420 42721
rect 30656 42712 30708 42764
rect 31208 42712 31260 42764
rect 27896 42644 27948 42653
rect 29184 42644 29236 42696
rect 20076 42508 20128 42560
rect 22744 42508 22796 42560
rect 23112 42508 23164 42560
rect 24308 42551 24360 42560
rect 24308 42517 24317 42551
rect 24317 42517 24351 42551
rect 24351 42517 24360 42551
rect 24308 42508 24360 42517
rect 26332 42551 26384 42560
rect 26332 42517 26341 42551
rect 26341 42517 26375 42551
rect 26375 42517 26384 42551
rect 26332 42508 26384 42517
rect 26516 42508 26568 42560
rect 27436 42508 27488 42560
rect 30380 42508 30432 42560
rect 6102 42406 6154 42458
rect 6166 42406 6218 42458
rect 6230 42406 6282 42458
rect 6294 42406 6346 42458
rect 6358 42406 6410 42458
rect 16405 42406 16457 42458
rect 16469 42406 16521 42458
rect 16533 42406 16585 42458
rect 16597 42406 16649 42458
rect 16661 42406 16713 42458
rect 26709 42406 26761 42458
rect 26773 42406 26825 42458
rect 26837 42406 26889 42458
rect 26901 42406 26953 42458
rect 26965 42406 27017 42458
rect 4988 42347 5040 42356
rect 4988 42313 4997 42347
rect 4997 42313 5031 42347
rect 5031 42313 5040 42347
rect 4988 42304 5040 42313
rect 7288 42347 7340 42356
rect 7288 42313 7297 42347
rect 7297 42313 7331 42347
rect 7331 42313 7340 42347
rect 7288 42304 7340 42313
rect 9956 42304 10008 42356
rect 7656 42236 7708 42288
rect 8576 42236 8628 42288
rect 9404 42236 9456 42288
rect 5632 42168 5684 42220
rect 7380 42168 7432 42220
rect 11060 42304 11112 42356
rect 11888 42304 11940 42356
rect 2136 42100 2188 42152
rect 5540 42100 5592 42152
rect 6644 42143 6696 42152
rect 6644 42109 6653 42143
rect 6653 42109 6687 42143
rect 6687 42109 6696 42143
rect 6644 42100 6696 42109
rect 7472 42143 7524 42152
rect 7472 42109 7481 42143
rect 7481 42109 7515 42143
rect 7515 42109 7524 42143
rect 7472 42100 7524 42109
rect 7656 42143 7708 42152
rect 7656 42109 7665 42143
rect 7665 42109 7699 42143
rect 7699 42109 7708 42143
rect 7656 42100 7708 42109
rect 8024 42143 8076 42152
rect 6552 42032 6604 42084
rect 8024 42109 8033 42143
rect 8033 42109 8067 42143
rect 8067 42109 8076 42143
rect 8024 42100 8076 42109
rect 8944 42143 8996 42152
rect 8944 42109 8953 42143
rect 8953 42109 8987 42143
rect 8987 42109 8996 42143
rect 8944 42100 8996 42109
rect 9128 42143 9180 42152
rect 9128 42109 9137 42143
rect 9137 42109 9171 42143
rect 9171 42109 9180 42143
rect 9128 42100 9180 42109
rect 9496 42143 9548 42152
rect 8116 42032 8168 42084
rect 9496 42109 9505 42143
rect 9505 42109 9539 42143
rect 9539 42109 9548 42143
rect 9496 42100 9548 42109
rect 13084 42168 13136 42220
rect 15016 42168 15068 42220
rect 10140 42143 10192 42152
rect 10140 42109 10149 42143
rect 10149 42109 10183 42143
rect 10183 42109 10192 42143
rect 10140 42100 10192 42109
rect 10232 42100 10284 42152
rect 10784 42100 10836 42152
rect 12072 42100 12124 42152
rect 13360 42100 13412 42152
rect 14556 42143 14608 42152
rect 9404 42032 9456 42084
rect 9588 42032 9640 42084
rect 12992 42032 13044 42084
rect 14556 42109 14565 42143
rect 14565 42109 14599 42143
rect 14599 42109 14608 42143
rect 14556 42100 14608 42109
rect 14648 42143 14700 42152
rect 14648 42109 14657 42143
rect 14657 42109 14691 42143
rect 14691 42109 14700 42143
rect 14648 42100 14700 42109
rect 4804 41964 4856 42016
rect 6000 41964 6052 42016
rect 9496 41964 9548 42016
rect 9680 42007 9732 42016
rect 9680 41973 9689 42007
rect 9689 41973 9723 42007
rect 9723 41973 9732 42007
rect 9680 41964 9732 41973
rect 10968 41964 11020 42016
rect 13728 41964 13780 42016
rect 14740 42032 14792 42084
rect 16120 42168 16172 42220
rect 16396 42236 16448 42288
rect 19432 42304 19484 42356
rect 21272 42347 21324 42356
rect 21272 42313 21281 42347
rect 21281 42313 21315 42347
rect 21315 42313 21324 42347
rect 21272 42304 21324 42313
rect 23020 42304 23072 42356
rect 23388 42279 23440 42288
rect 16212 42143 16264 42152
rect 16212 42109 16221 42143
rect 16221 42109 16255 42143
rect 16255 42109 16264 42143
rect 16212 42100 16264 42109
rect 18512 42168 18564 42220
rect 21456 42168 21508 42220
rect 23388 42245 23397 42279
rect 23397 42245 23431 42279
rect 23431 42245 23440 42279
rect 23388 42236 23440 42245
rect 24032 42236 24084 42288
rect 16856 42100 16908 42152
rect 17684 42100 17736 42152
rect 15384 42007 15436 42016
rect 15384 41973 15393 42007
rect 15393 41973 15427 42007
rect 15427 41973 15436 42007
rect 15384 41964 15436 41973
rect 15844 42007 15896 42016
rect 15844 41973 15853 42007
rect 15853 41973 15887 42007
rect 15887 41973 15896 42007
rect 15844 41964 15896 41973
rect 16212 41964 16264 42016
rect 16948 41964 17000 42016
rect 17132 41964 17184 42016
rect 17500 41964 17552 42016
rect 17960 42032 18012 42084
rect 20720 42100 20772 42152
rect 21824 42100 21876 42152
rect 22192 42168 22244 42220
rect 22836 42168 22888 42220
rect 22928 42168 22980 42220
rect 23112 42143 23164 42152
rect 20168 42075 20220 42084
rect 20168 42041 20202 42075
rect 20202 42041 20220 42075
rect 20168 42032 20220 42041
rect 23112 42109 23121 42143
rect 23121 42109 23155 42143
rect 23155 42109 23164 42143
rect 23112 42100 23164 42109
rect 23296 42100 23348 42152
rect 26332 42304 26384 42356
rect 26608 42304 26660 42356
rect 24400 42143 24452 42152
rect 24400 42109 24409 42143
rect 24409 42109 24443 42143
rect 24443 42109 24452 42143
rect 24400 42100 24452 42109
rect 25044 42100 25096 42152
rect 26240 42133 26292 42152
rect 26240 42100 26249 42133
rect 26249 42100 26283 42133
rect 26283 42100 26292 42133
rect 23940 42032 23992 42084
rect 24308 42032 24360 42084
rect 26424 42111 26437 42130
rect 26437 42111 26471 42130
rect 26471 42111 26476 42130
rect 26424 42078 26476 42111
rect 26700 42100 26752 42152
rect 26792 42143 26844 42152
rect 26792 42109 26801 42143
rect 26801 42109 26835 42143
rect 26835 42109 26844 42143
rect 26792 42100 26844 42109
rect 26884 42032 26936 42084
rect 18604 41964 18656 42016
rect 19524 41964 19576 42016
rect 22192 41964 22244 42016
rect 22560 41964 22612 42016
rect 23388 41964 23440 42016
rect 23664 41964 23716 42016
rect 24216 41964 24268 42016
rect 29368 42304 29420 42356
rect 27896 42236 27948 42288
rect 28908 42168 28960 42220
rect 29920 42211 29972 42220
rect 29920 42177 29929 42211
rect 29929 42177 29963 42211
rect 29963 42177 29972 42211
rect 29920 42168 29972 42177
rect 27160 42100 27212 42152
rect 29092 42100 29144 42152
rect 29276 42100 29328 42152
rect 30472 42100 30524 42152
rect 31116 42143 31168 42152
rect 31116 42109 31125 42143
rect 31125 42109 31159 42143
rect 31159 42109 31168 42143
rect 31116 42100 31168 42109
rect 27344 41964 27396 42016
rect 27528 42007 27580 42016
rect 27528 41973 27537 42007
rect 27537 41973 27571 42007
rect 27571 41973 27580 42007
rect 27528 41964 27580 41973
rect 28264 41964 28316 42016
rect 30012 42032 30064 42084
rect 29184 41964 29236 42016
rect 30288 42007 30340 42016
rect 30288 41973 30297 42007
rect 30297 41973 30331 42007
rect 30331 41973 30340 42007
rect 30288 41964 30340 41973
rect 11253 41862 11305 41914
rect 11317 41862 11369 41914
rect 11381 41862 11433 41914
rect 11445 41862 11497 41914
rect 11509 41862 11561 41914
rect 21557 41862 21609 41914
rect 21621 41862 21673 41914
rect 21685 41862 21737 41914
rect 21749 41862 21801 41914
rect 21813 41862 21865 41914
rect 2688 41803 2740 41812
rect 2688 41769 2697 41803
rect 2697 41769 2731 41803
rect 2731 41769 2740 41803
rect 2688 41760 2740 41769
rect 8760 41760 8812 41812
rect 8944 41760 8996 41812
rect 12532 41760 12584 41812
rect 20536 41760 20588 41812
rect 5816 41692 5868 41744
rect 3700 41667 3752 41676
rect 3700 41633 3709 41667
rect 3709 41633 3743 41667
rect 3743 41633 3752 41667
rect 3700 41624 3752 41633
rect 4528 41624 4580 41676
rect 6644 41624 6696 41676
rect 8116 41624 8168 41676
rect 8576 41667 8628 41676
rect 8576 41633 8585 41667
rect 8585 41633 8619 41667
rect 8619 41633 8628 41667
rect 8576 41624 8628 41633
rect 8852 41624 8904 41676
rect 9312 41624 9364 41676
rect 9496 41624 9548 41676
rect 9772 41692 9824 41744
rect 10416 41692 10468 41744
rect 14188 41735 14240 41744
rect 14188 41701 14197 41735
rect 14197 41701 14231 41735
rect 14231 41701 14240 41735
rect 14188 41692 14240 41701
rect 15752 41692 15804 41744
rect 16304 41692 16356 41744
rect 5356 41556 5408 41608
rect 8300 41556 8352 41608
rect 8668 41599 8720 41608
rect 8668 41565 8677 41599
rect 8677 41565 8711 41599
rect 8711 41565 8720 41599
rect 8668 41556 8720 41565
rect 9220 41556 9272 41608
rect 10048 41624 10100 41676
rect 12808 41624 12860 41676
rect 13084 41667 13136 41676
rect 13084 41633 13093 41667
rect 13093 41633 13127 41667
rect 13127 41633 13136 41667
rect 13084 41624 13136 41633
rect 13360 41667 13412 41676
rect 13360 41633 13369 41667
rect 13369 41633 13403 41667
rect 13403 41633 13412 41667
rect 13360 41624 13412 41633
rect 16212 41624 16264 41676
rect 17316 41692 17368 41744
rect 10324 41556 10376 41608
rect 12624 41556 12676 41608
rect 15200 41556 15252 41608
rect 17040 41599 17092 41608
rect 17040 41565 17049 41599
rect 17049 41565 17083 41599
rect 17083 41565 17092 41599
rect 17040 41556 17092 41565
rect 1860 41420 1912 41472
rect 3240 41463 3292 41472
rect 3240 41429 3249 41463
rect 3249 41429 3283 41463
rect 3283 41429 3292 41463
rect 3240 41420 3292 41429
rect 5632 41420 5684 41472
rect 6644 41488 6696 41540
rect 10140 41488 10192 41540
rect 9864 41463 9916 41472
rect 9864 41429 9873 41463
rect 9873 41429 9907 41463
rect 9907 41429 9916 41463
rect 10600 41488 10652 41540
rect 19340 41624 19392 41676
rect 20260 41667 20312 41676
rect 20260 41633 20269 41667
rect 20269 41633 20303 41667
rect 20303 41633 20312 41667
rect 20260 41624 20312 41633
rect 23296 41692 23348 41744
rect 21272 41624 21324 41676
rect 18604 41556 18656 41608
rect 22100 41624 22152 41676
rect 23480 41624 23532 41676
rect 23940 41803 23992 41812
rect 23940 41769 23949 41803
rect 23949 41769 23983 41803
rect 23983 41769 23992 41803
rect 23940 41760 23992 41769
rect 25872 41760 25924 41812
rect 26792 41760 26844 41812
rect 30012 41803 30064 41812
rect 25412 41692 25464 41744
rect 29000 41692 29052 41744
rect 30012 41769 30021 41803
rect 30021 41769 30055 41803
rect 30055 41769 30064 41803
rect 30012 41760 30064 41769
rect 30932 41760 30984 41812
rect 31116 41692 31168 41744
rect 24860 41624 24912 41676
rect 25044 41667 25096 41676
rect 25044 41633 25053 41667
rect 25053 41633 25087 41667
rect 25087 41633 25096 41667
rect 25044 41624 25096 41633
rect 25780 41624 25832 41676
rect 26792 41624 26844 41676
rect 30472 41624 30524 41676
rect 22284 41556 22336 41608
rect 26148 41556 26200 41608
rect 26700 41556 26752 41608
rect 28632 41599 28684 41608
rect 28632 41565 28641 41599
rect 28641 41565 28675 41599
rect 28675 41565 28684 41599
rect 28632 41556 28684 41565
rect 22008 41488 22060 41540
rect 23388 41488 23440 41540
rect 26240 41488 26292 41540
rect 26884 41488 26936 41540
rect 27804 41488 27856 41540
rect 10416 41463 10468 41472
rect 9864 41420 9916 41429
rect 10416 41429 10425 41463
rect 10425 41429 10459 41463
rect 10459 41429 10468 41463
rect 10416 41420 10468 41429
rect 10784 41463 10836 41472
rect 10784 41429 10793 41463
rect 10793 41429 10827 41463
rect 10827 41429 10836 41463
rect 10784 41420 10836 41429
rect 15476 41463 15528 41472
rect 15476 41429 15485 41463
rect 15485 41429 15519 41463
rect 15519 41429 15528 41463
rect 15476 41420 15528 41429
rect 15752 41420 15804 41472
rect 19340 41420 19392 41472
rect 22744 41420 22796 41472
rect 24952 41420 25004 41472
rect 25044 41420 25096 41472
rect 25320 41420 25372 41472
rect 26424 41463 26476 41472
rect 26424 41429 26433 41463
rect 26433 41429 26467 41463
rect 26467 41429 26476 41463
rect 26424 41420 26476 41429
rect 26608 41420 26660 41472
rect 27160 41463 27212 41472
rect 27160 41429 27169 41463
rect 27169 41429 27203 41463
rect 27203 41429 27212 41463
rect 27160 41420 27212 41429
rect 27896 41420 27948 41472
rect 30472 41463 30524 41472
rect 30472 41429 30481 41463
rect 30481 41429 30515 41463
rect 30515 41429 30524 41463
rect 30472 41420 30524 41429
rect 6102 41318 6154 41370
rect 6166 41318 6218 41370
rect 6230 41318 6282 41370
rect 6294 41318 6346 41370
rect 6358 41318 6410 41370
rect 16405 41318 16457 41370
rect 16469 41318 16521 41370
rect 16533 41318 16585 41370
rect 16597 41318 16649 41370
rect 16661 41318 16713 41370
rect 26709 41318 26761 41370
rect 26773 41318 26825 41370
rect 26837 41318 26889 41370
rect 26901 41318 26953 41370
rect 26965 41318 27017 41370
rect 3240 41216 3292 41268
rect 4344 41216 4396 41268
rect 4436 41216 4488 41268
rect 3976 41080 4028 41132
rect 3516 40944 3568 40996
rect 3792 40944 3844 40996
rect 4436 41012 4488 41064
rect 5080 41012 5132 41064
rect 5448 41012 5500 41064
rect 9220 41216 9272 41268
rect 13820 41216 13872 41268
rect 14832 41216 14884 41268
rect 16856 41216 16908 41268
rect 17040 41216 17092 41268
rect 17224 41216 17276 41268
rect 18604 41259 18656 41268
rect 9680 41148 9732 41200
rect 12808 41148 12860 41200
rect 14280 41148 14332 41200
rect 17776 41191 17828 41200
rect 17776 41157 17785 41191
rect 17785 41157 17819 41191
rect 17819 41157 17828 41191
rect 17776 41148 17828 41157
rect 18604 41225 18613 41259
rect 18613 41225 18647 41259
rect 18647 41225 18656 41259
rect 18604 41216 18656 41225
rect 19248 41259 19300 41268
rect 19248 41225 19257 41259
rect 19257 41225 19291 41259
rect 19291 41225 19300 41259
rect 19248 41216 19300 41225
rect 19524 41148 19576 41200
rect 8300 41080 8352 41132
rect 11060 41080 11112 41132
rect 11612 41080 11664 41132
rect 16120 41080 16172 41132
rect 16856 41080 16908 41132
rect 8484 41012 8536 41064
rect 8852 41012 8904 41064
rect 2504 40919 2556 40928
rect 2504 40885 2513 40919
rect 2513 40885 2547 40919
rect 2547 40885 2556 40919
rect 2504 40876 2556 40885
rect 3608 40876 3660 40928
rect 5908 40944 5960 40996
rect 7840 40944 7892 40996
rect 8576 40944 8628 40996
rect 9312 41012 9364 41064
rect 10232 41055 10284 41064
rect 10232 41021 10241 41055
rect 10241 41021 10275 41055
rect 10275 41021 10284 41055
rect 10232 41012 10284 41021
rect 10416 41055 10468 41064
rect 10416 41021 10425 41055
rect 10425 41021 10459 41055
rect 10459 41021 10468 41055
rect 10416 41012 10468 41021
rect 10600 41055 10652 41064
rect 10600 41021 10609 41055
rect 10609 41021 10643 41055
rect 10643 41021 10652 41055
rect 10600 41012 10652 41021
rect 10692 41055 10744 41064
rect 10692 41021 10701 41055
rect 10701 41021 10735 41055
rect 10735 41021 10744 41055
rect 10692 41012 10744 41021
rect 13084 41012 13136 41064
rect 15476 41055 15528 41064
rect 15476 41021 15485 41055
rect 15485 41021 15519 41055
rect 15519 41021 15528 41055
rect 15476 41012 15528 41021
rect 10140 40944 10192 40996
rect 12256 40944 12308 40996
rect 14372 40944 14424 40996
rect 5724 40919 5776 40928
rect 5724 40885 5733 40919
rect 5733 40885 5767 40919
rect 5767 40885 5776 40919
rect 5724 40876 5776 40885
rect 6828 40876 6880 40928
rect 7104 40919 7156 40928
rect 7104 40885 7113 40919
rect 7113 40885 7147 40919
rect 7147 40885 7156 40919
rect 7104 40876 7156 40885
rect 10876 40919 10928 40928
rect 10876 40885 10885 40919
rect 10885 40885 10919 40919
rect 10919 40885 10928 40919
rect 10876 40876 10928 40885
rect 14740 40876 14792 40928
rect 16948 41012 17000 41064
rect 17224 41012 17276 41064
rect 17316 40987 17368 40996
rect 17316 40953 17325 40987
rect 17325 40953 17359 40987
rect 17359 40953 17368 40987
rect 17316 40944 17368 40953
rect 17684 40944 17736 40996
rect 17960 40987 18012 40996
rect 17960 40953 17969 40987
rect 17969 40953 18003 40987
rect 18003 40953 18012 40987
rect 17960 40944 18012 40953
rect 19248 41080 19300 41132
rect 19432 41055 19484 41064
rect 19432 41021 19441 41055
rect 19441 41021 19475 41055
rect 19475 41021 19484 41055
rect 19432 41012 19484 41021
rect 19340 40944 19392 40996
rect 20996 41216 21048 41268
rect 21272 41216 21324 41268
rect 20444 41148 20496 41200
rect 20076 41080 20128 41132
rect 21088 41148 21140 41200
rect 23480 41216 23532 41268
rect 24308 41216 24360 41268
rect 25780 41259 25832 41268
rect 25780 41225 25789 41259
rect 25789 41225 25823 41259
rect 25823 41225 25832 41259
rect 25780 41216 25832 41225
rect 24584 41148 24636 41200
rect 26332 41148 26384 41200
rect 23020 41080 23072 41132
rect 20352 41012 20404 41064
rect 20444 41012 20496 41064
rect 22284 41012 22336 41064
rect 22468 41012 22520 41064
rect 23112 41055 23164 41064
rect 23112 41021 23121 41055
rect 23121 41021 23155 41055
rect 23155 41021 23164 41055
rect 23112 41012 23164 41021
rect 23480 41012 23532 41064
rect 25136 41080 25188 41132
rect 26148 41123 26200 41132
rect 26148 41089 26157 41123
rect 26157 41089 26191 41123
rect 26191 41089 26200 41123
rect 26148 41080 26200 41089
rect 26240 41055 26292 41064
rect 24216 40944 24268 40996
rect 26240 41021 26249 41055
rect 26249 41021 26283 41055
rect 26283 41021 26292 41055
rect 26240 41012 26292 41021
rect 26332 41055 26384 41064
rect 26332 41021 26341 41055
rect 26341 41021 26375 41055
rect 26375 41021 26384 41055
rect 28632 41123 28684 41132
rect 28632 41089 28641 41123
rect 28641 41089 28675 41123
rect 28675 41089 28684 41123
rect 28632 41080 28684 41089
rect 26332 41012 26384 41021
rect 27068 41012 27120 41064
rect 30288 41012 30340 41064
rect 26608 40944 26660 40996
rect 16212 40876 16264 40928
rect 16948 40876 17000 40928
rect 18604 40876 18656 40928
rect 19708 40876 19760 40928
rect 21916 40876 21968 40928
rect 22284 40876 22336 40928
rect 30564 40876 30616 40928
rect 31024 40919 31076 40928
rect 31024 40885 31033 40919
rect 31033 40885 31067 40919
rect 31067 40885 31076 40919
rect 31024 40876 31076 40885
rect 11253 40774 11305 40826
rect 11317 40774 11369 40826
rect 11381 40774 11433 40826
rect 11445 40774 11497 40826
rect 11509 40774 11561 40826
rect 21557 40774 21609 40826
rect 21621 40774 21673 40826
rect 21685 40774 21737 40826
rect 21749 40774 21801 40826
rect 21813 40774 21865 40826
rect 1400 40536 1452 40588
rect 2872 40672 2924 40724
rect 3976 40672 4028 40724
rect 8484 40672 8536 40724
rect 10232 40672 10284 40724
rect 12256 40715 12308 40724
rect 12256 40681 12265 40715
rect 12265 40681 12299 40715
rect 12299 40681 12308 40715
rect 12256 40672 12308 40681
rect 2780 40604 2832 40656
rect 3700 40604 3752 40656
rect 3240 40536 3292 40588
rect 3332 40536 3384 40588
rect 3792 40536 3844 40588
rect 5448 40604 5500 40656
rect 4068 40468 4120 40520
rect 4804 40579 4856 40588
rect 4804 40545 4813 40579
rect 4813 40545 4847 40579
rect 4847 40545 4856 40579
rect 4804 40536 4856 40545
rect 5080 40536 5132 40588
rect 5632 40536 5684 40588
rect 8300 40604 8352 40656
rect 8668 40604 8720 40656
rect 8484 40579 8536 40588
rect 8484 40545 8493 40579
rect 8493 40545 8527 40579
rect 8527 40545 8536 40579
rect 8484 40536 8536 40545
rect 10324 40604 10376 40656
rect 8944 40536 8996 40588
rect 9312 40536 9364 40588
rect 10140 40579 10192 40588
rect 10140 40545 10149 40579
rect 10149 40545 10183 40579
rect 10183 40545 10192 40579
rect 10140 40536 10192 40545
rect 13820 40672 13872 40724
rect 14740 40672 14792 40724
rect 13728 40647 13780 40656
rect 13728 40613 13762 40647
rect 13762 40613 13780 40647
rect 13728 40604 13780 40613
rect 17224 40672 17276 40724
rect 17408 40672 17460 40724
rect 19248 40672 19300 40724
rect 21180 40672 21232 40724
rect 16120 40647 16172 40656
rect 16120 40613 16129 40647
rect 16129 40613 16163 40647
rect 16163 40613 16172 40647
rect 16120 40604 16172 40613
rect 17132 40604 17184 40656
rect 9864 40468 9916 40520
rect 10324 40511 10376 40520
rect 10324 40477 10333 40511
rect 10333 40477 10367 40511
rect 10367 40477 10376 40511
rect 10324 40468 10376 40477
rect 10968 40468 11020 40520
rect 12808 40579 12860 40588
rect 12808 40545 12817 40579
rect 12817 40545 12851 40579
rect 12851 40545 12860 40579
rect 12808 40536 12860 40545
rect 12992 40579 13044 40588
rect 12992 40545 13001 40579
rect 13001 40545 13035 40579
rect 13035 40545 13044 40579
rect 12992 40536 13044 40545
rect 13544 40536 13596 40588
rect 16856 40579 16908 40588
rect 16856 40545 16865 40579
rect 16865 40545 16899 40579
rect 16899 40545 16908 40579
rect 16856 40536 16908 40545
rect 18052 40604 18104 40656
rect 22100 40604 22152 40656
rect 22468 40672 22520 40724
rect 22652 40672 22704 40724
rect 27252 40672 27304 40724
rect 23480 40604 23532 40656
rect 24216 40604 24268 40656
rect 17316 40536 17368 40588
rect 18512 40536 18564 40588
rect 19432 40536 19484 40588
rect 22008 40579 22060 40588
rect 22008 40545 22017 40579
rect 22017 40545 22051 40579
rect 22051 40545 22060 40579
rect 22008 40536 22060 40545
rect 22192 40579 22244 40588
rect 22192 40545 22201 40579
rect 22201 40545 22235 40579
rect 22235 40545 22244 40579
rect 22192 40536 22244 40545
rect 22284 40579 22336 40588
rect 22284 40545 22293 40579
rect 22293 40545 22327 40579
rect 22327 40545 22336 40579
rect 22284 40536 22336 40545
rect 22468 40579 22520 40588
rect 22468 40545 22477 40579
rect 22477 40545 22511 40579
rect 22511 40545 22520 40579
rect 22468 40536 22520 40545
rect 23112 40536 23164 40588
rect 26056 40604 26108 40656
rect 12624 40511 12676 40520
rect 12624 40477 12633 40511
rect 12633 40477 12667 40511
rect 12667 40477 12676 40511
rect 12624 40468 12676 40477
rect 8852 40400 8904 40452
rect 1952 40375 2004 40384
rect 1952 40341 1961 40375
rect 1961 40341 1995 40375
rect 1995 40341 2004 40375
rect 1952 40332 2004 40341
rect 5264 40332 5316 40384
rect 5540 40332 5592 40384
rect 10232 40332 10284 40384
rect 10692 40400 10744 40452
rect 12072 40400 12124 40452
rect 12532 40400 12584 40452
rect 10600 40332 10652 40384
rect 11428 40332 11480 40384
rect 13084 40468 13136 40520
rect 17776 40468 17828 40520
rect 14556 40332 14608 40384
rect 16028 40332 16080 40384
rect 16212 40332 16264 40384
rect 17960 40332 18012 40384
rect 23204 40468 23256 40520
rect 24860 40468 24912 40520
rect 24952 40468 25004 40520
rect 25504 40536 25556 40588
rect 27344 40604 27396 40656
rect 25320 40511 25372 40520
rect 25320 40477 25329 40511
rect 25329 40477 25363 40511
rect 25363 40477 25372 40511
rect 25320 40468 25372 40477
rect 26056 40468 26108 40520
rect 27252 40579 27304 40588
rect 27252 40545 27261 40579
rect 27261 40545 27295 40579
rect 27295 40545 27304 40579
rect 27252 40536 27304 40545
rect 27436 40536 27488 40588
rect 28632 40536 28684 40588
rect 30288 40536 30340 40588
rect 26332 40468 26384 40520
rect 28172 40511 28224 40520
rect 28172 40477 28181 40511
rect 28181 40477 28215 40511
rect 28215 40477 28224 40511
rect 28172 40468 28224 40477
rect 28540 40468 28592 40520
rect 28908 40468 28960 40520
rect 27620 40400 27672 40452
rect 20076 40332 20128 40384
rect 21180 40375 21232 40384
rect 21180 40341 21189 40375
rect 21189 40341 21223 40375
rect 21223 40341 21232 40375
rect 21180 40332 21232 40341
rect 22008 40332 22060 40384
rect 22284 40332 22336 40384
rect 23296 40332 23348 40384
rect 25780 40375 25832 40384
rect 25780 40341 25789 40375
rect 25789 40341 25823 40375
rect 25823 40341 25832 40375
rect 25780 40332 25832 40341
rect 27344 40332 27396 40384
rect 30564 40332 30616 40384
rect 6102 40230 6154 40282
rect 6166 40230 6218 40282
rect 6230 40230 6282 40282
rect 6294 40230 6346 40282
rect 6358 40230 6410 40282
rect 16405 40230 16457 40282
rect 16469 40230 16521 40282
rect 16533 40230 16585 40282
rect 16597 40230 16649 40282
rect 16661 40230 16713 40282
rect 26709 40230 26761 40282
rect 26773 40230 26825 40282
rect 26837 40230 26889 40282
rect 26901 40230 26953 40282
rect 26965 40230 27017 40282
rect 4068 40128 4120 40180
rect 4344 40060 4396 40112
rect 4988 40060 5040 40112
rect 2504 39992 2556 40044
rect 4068 40035 4120 40044
rect 2228 39967 2280 39976
rect 1400 39788 1452 39840
rect 1676 39831 1728 39840
rect 1676 39797 1685 39831
rect 1685 39797 1719 39831
rect 1719 39797 1728 39831
rect 1676 39788 1728 39797
rect 2228 39933 2237 39967
rect 2237 39933 2271 39967
rect 2271 39933 2280 39967
rect 2228 39924 2280 39933
rect 2412 39967 2464 39976
rect 2412 39933 2421 39967
rect 2421 39933 2455 39967
rect 2455 39933 2464 39967
rect 2412 39924 2464 39933
rect 3424 39924 3476 39976
rect 3700 39924 3752 39976
rect 4068 40001 4077 40035
rect 4077 40001 4111 40035
rect 4111 40001 4120 40035
rect 4068 39992 4120 40001
rect 4528 40035 4580 40044
rect 4528 40001 4537 40035
rect 4537 40001 4571 40035
rect 4571 40001 4580 40035
rect 4528 39992 4580 40001
rect 5632 39992 5684 40044
rect 6644 39992 6696 40044
rect 3884 39924 3936 39976
rect 3976 39967 4028 39976
rect 3976 39933 3985 39967
rect 3985 39933 4019 39967
rect 4019 39933 4028 39967
rect 3976 39924 4028 39933
rect 4344 39967 4396 39976
rect 4344 39933 4353 39967
rect 4353 39933 4387 39967
rect 4387 39933 4396 39967
rect 4344 39924 4396 39933
rect 4988 39924 5040 39976
rect 2596 39788 2648 39840
rect 2688 39788 2740 39840
rect 5632 39831 5684 39840
rect 5632 39797 5641 39831
rect 5641 39797 5675 39831
rect 5675 39797 5684 39831
rect 7840 39924 7892 39976
rect 9404 40060 9456 40112
rect 10324 40128 10376 40180
rect 16304 40128 16356 40180
rect 17316 40128 17368 40180
rect 23112 40171 23164 40180
rect 23112 40137 23121 40171
rect 23121 40137 23155 40171
rect 23155 40137 23164 40171
rect 23112 40128 23164 40137
rect 10140 40060 10192 40112
rect 9680 39992 9732 40044
rect 12440 40035 12492 40044
rect 12440 40001 12449 40035
rect 12449 40001 12483 40035
rect 12483 40001 12492 40035
rect 12440 39992 12492 40001
rect 12624 39992 12676 40044
rect 14372 39992 14424 40044
rect 9496 39933 9499 39954
rect 9499 39933 9533 39954
rect 9533 39933 9548 39954
rect 6644 39899 6696 39908
rect 6644 39865 6653 39899
rect 6653 39865 6687 39899
rect 6687 39865 6696 39899
rect 6644 39856 6696 39865
rect 9496 39902 9548 39933
rect 9588 39933 9597 39954
rect 9597 39933 9631 39954
rect 9631 39933 9640 39954
rect 9588 39902 9640 39933
rect 10784 39967 10836 39976
rect 10784 39933 10793 39967
rect 10793 39933 10827 39967
rect 10827 39933 10836 39967
rect 10784 39924 10836 39933
rect 11428 39967 11480 39976
rect 11428 39933 11437 39967
rect 11437 39933 11471 39967
rect 11471 39933 11480 39967
rect 11428 39924 11480 39933
rect 11980 39924 12032 39976
rect 12992 39924 13044 39976
rect 14004 39924 14056 39976
rect 14280 39967 14332 39976
rect 14280 39933 14289 39967
rect 14289 39933 14323 39967
rect 14323 39933 14332 39967
rect 14280 39924 14332 39933
rect 14556 40060 14608 40112
rect 21456 40060 21508 40112
rect 24768 40128 24820 40180
rect 30288 40171 30340 40180
rect 30288 40137 30297 40171
rect 30297 40137 30331 40171
rect 30331 40137 30340 40171
rect 30288 40128 30340 40137
rect 30380 40128 30432 40180
rect 30656 40128 30708 40180
rect 23572 40060 23624 40112
rect 14740 39924 14792 39976
rect 5632 39788 5684 39797
rect 6368 39788 6420 39840
rect 7012 39788 7064 39840
rect 10692 39856 10744 39908
rect 13544 39856 13596 39908
rect 16948 39924 17000 39976
rect 17592 39924 17644 39976
rect 17960 39967 18012 39976
rect 17960 39933 17978 39967
rect 17978 39933 18012 39967
rect 17960 39924 18012 39933
rect 19524 39924 19576 39976
rect 17684 39856 17736 39908
rect 19340 39856 19392 39908
rect 19616 39899 19668 39908
rect 19616 39865 19625 39899
rect 19625 39865 19659 39899
rect 19659 39865 19668 39899
rect 19616 39856 19668 39865
rect 13452 39788 13504 39840
rect 13728 39788 13780 39840
rect 14004 39788 14056 39840
rect 21180 39924 21232 39976
rect 21916 39924 21968 39976
rect 20720 39856 20772 39908
rect 20628 39788 20680 39840
rect 22008 39788 22060 39840
rect 22560 39992 22612 40044
rect 23940 39992 23992 40044
rect 22192 39967 22244 39976
rect 22192 39933 22201 39967
rect 22201 39933 22235 39967
rect 22235 39933 22244 39967
rect 22192 39924 22244 39933
rect 23112 39924 23164 39976
rect 23296 39967 23348 39976
rect 23296 39933 23305 39967
rect 23305 39933 23339 39967
rect 23339 39933 23348 39967
rect 23296 39924 23348 39933
rect 22928 39856 22980 39908
rect 23664 39967 23716 39976
rect 23664 39933 23673 39967
rect 23673 39933 23707 39967
rect 23707 39933 23716 39967
rect 23664 39924 23716 39933
rect 24216 39924 24268 39976
rect 26240 39992 26292 40044
rect 28172 39992 28224 40044
rect 24584 39967 24636 39976
rect 24584 39933 24593 39967
rect 24593 39933 24627 39967
rect 24627 39933 24636 39967
rect 24584 39924 24636 39933
rect 24860 39924 24912 39976
rect 25780 39924 25832 39976
rect 26516 39924 26568 39976
rect 29460 39992 29512 40044
rect 28448 39924 28500 39976
rect 29276 39924 29328 39976
rect 31024 39992 31076 40044
rect 28632 39856 28684 39908
rect 29920 39967 29972 39976
rect 29920 39933 29929 39967
rect 29929 39933 29963 39967
rect 29963 39933 29972 39967
rect 29920 39924 29972 39933
rect 30472 39924 30524 39976
rect 31300 39924 31352 39976
rect 22560 39831 22612 39840
rect 22560 39797 22569 39831
rect 22569 39797 22603 39831
rect 22603 39797 22612 39831
rect 22560 39788 22612 39797
rect 22836 39788 22888 39840
rect 25320 39788 25372 39840
rect 26332 39788 26384 39840
rect 27436 39788 27488 39840
rect 29644 39788 29696 39840
rect 11253 39686 11305 39738
rect 11317 39686 11369 39738
rect 11381 39686 11433 39738
rect 11445 39686 11497 39738
rect 11509 39686 11561 39738
rect 21557 39686 21609 39738
rect 21621 39686 21673 39738
rect 21685 39686 21737 39738
rect 21749 39686 21801 39738
rect 21813 39686 21865 39738
rect 3240 39627 3292 39636
rect 3240 39593 3249 39627
rect 3249 39593 3283 39627
rect 3283 39593 3292 39627
rect 3240 39584 3292 39593
rect 4252 39584 4304 39636
rect 4528 39584 4580 39636
rect 9588 39584 9640 39636
rect 15200 39584 15252 39636
rect 22468 39584 22520 39636
rect 22652 39584 22704 39636
rect 23940 39584 23992 39636
rect 24308 39627 24360 39636
rect 24308 39593 24317 39627
rect 24317 39593 24351 39627
rect 24351 39593 24360 39627
rect 24308 39584 24360 39593
rect 2780 39516 2832 39568
rect 3148 39516 3200 39568
rect 3332 39516 3384 39568
rect 1400 39491 1452 39500
rect 1400 39457 1409 39491
rect 1409 39457 1443 39491
rect 1443 39457 1452 39491
rect 1400 39448 1452 39457
rect 1676 39491 1728 39500
rect 1676 39457 1710 39491
rect 1710 39457 1728 39491
rect 1676 39448 1728 39457
rect 2136 39448 2188 39500
rect 2688 39448 2740 39500
rect 3424 39491 3476 39500
rect 3424 39457 3433 39491
rect 3433 39457 3467 39491
rect 3467 39457 3476 39491
rect 3424 39448 3476 39457
rect 4344 39516 4396 39568
rect 5080 39516 5132 39568
rect 3884 39448 3936 39500
rect 4988 39491 5040 39500
rect 4988 39457 4997 39491
rect 4997 39457 5031 39491
rect 5031 39457 5040 39491
rect 4988 39448 5040 39457
rect 6368 39516 6420 39568
rect 12440 39516 12492 39568
rect 17132 39516 17184 39568
rect 18328 39516 18380 39568
rect 19708 39516 19760 39568
rect 23388 39559 23440 39568
rect 7012 39491 7064 39500
rect 7012 39457 7021 39491
rect 7021 39457 7055 39491
rect 7055 39457 7064 39491
rect 7012 39448 7064 39457
rect 7472 39491 7524 39500
rect 7472 39457 7481 39491
rect 7481 39457 7515 39491
rect 7515 39457 7524 39491
rect 7472 39448 7524 39457
rect 8300 39491 8352 39500
rect 8300 39457 8309 39491
rect 8309 39457 8343 39491
rect 8343 39457 8352 39491
rect 8300 39448 8352 39457
rect 8392 39448 8444 39500
rect 10416 39448 10468 39500
rect 11152 39448 11204 39500
rect 13820 39448 13872 39500
rect 15108 39448 15160 39500
rect 15936 39448 15988 39500
rect 18236 39491 18288 39500
rect 18236 39457 18254 39491
rect 18254 39457 18288 39491
rect 18236 39448 18288 39457
rect 20536 39491 20588 39500
rect 20536 39457 20554 39491
rect 20554 39457 20588 39491
rect 20536 39448 20588 39457
rect 4252 39380 4304 39432
rect 4988 39312 5040 39364
rect 6460 39380 6512 39432
rect 7196 39423 7248 39432
rect 7196 39389 7205 39423
rect 7205 39389 7239 39423
rect 7239 39389 7248 39423
rect 7196 39380 7248 39389
rect 12440 39380 12492 39432
rect 13452 39380 13504 39432
rect 13728 39380 13780 39432
rect 15568 39380 15620 39432
rect 19616 39380 19668 39432
rect 8208 39312 8260 39364
rect 14832 39312 14884 39364
rect 15384 39312 15436 39364
rect 2688 39244 2740 39296
rect 3792 39244 3844 39296
rect 4068 39244 4120 39296
rect 8944 39244 8996 39296
rect 15200 39244 15252 39296
rect 15660 39287 15712 39296
rect 15660 39253 15669 39287
rect 15669 39253 15703 39287
rect 15703 39253 15712 39287
rect 15660 39244 15712 39253
rect 18144 39244 18196 39296
rect 18512 39244 18564 39296
rect 19616 39244 19668 39296
rect 20628 39244 20680 39296
rect 22376 39448 22428 39500
rect 22560 39491 22612 39500
rect 22560 39457 22569 39491
rect 22569 39457 22603 39491
rect 22603 39457 22612 39491
rect 22560 39448 22612 39457
rect 22744 39491 22796 39500
rect 22744 39457 22753 39491
rect 22753 39457 22787 39491
rect 22787 39457 22796 39491
rect 22744 39448 22796 39457
rect 23388 39525 23397 39559
rect 23397 39525 23431 39559
rect 23431 39525 23440 39559
rect 23388 39516 23440 39525
rect 23480 39516 23532 39568
rect 24952 39516 25004 39568
rect 26148 39559 26200 39568
rect 26148 39525 26157 39559
rect 26157 39525 26191 39559
rect 26191 39525 26200 39559
rect 26148 39516 26200 39525
rect 23664 39448 23716 39500
rect 23204 39380 23256 39432
rect 25320 39448 25372 39500
rect 28172 39584 28224 39636
rect 28356 39584 28408 39636
rect 29000 39627 29052 39636
rect 29000 39593 29009 39627
rect 29009 39593 29043 39627
rect 29043 39593 29052 39627
rect 29000 39584 29052 39593
rect 29460 39584 29512 39636
rect 27252 39516 27304 39568
rect 26424 39448 26476 39500
rect 27160 39491 27212 39500
rect 27160 39457 27169 39491
rect 27169 39457 27203 39491
rect 27203 39457 27212 39491
rect 27160 39448 27212 39457
rect 27528 39491 27580 39500
rect 27528 39457 27537 39491
rect 27537 39457 27571 39491
rect 27571 39457 27580 39491
rect 27528 39448 27580 39457
rect 27712 39491 27764 39500
rect 27712 39457 27721 39491
rect 27721 39457 27755 39491
rect 27755 39457 27764 39491
rect 27712 39448 27764 39457
rect 22560 39312 22612 39364
rect 23112 39312 23164 39364
rect 24400 39312 24452 39364
rect 27988 39380 28040 39432
rect 27804 39312 27856 39364
rect 22468 39244 22520 39296
rect 23020 39244 23072 39296
rect 27436 39244 27488 39296
rect 29184 39516 29236 39568
rect 29644 39559 29696 39568
rect 29644 39525 29653 39559
rect 29653 39525 29687 39559
rect 29687 39525 29696 39559
rect 29644 39516 29696 39525
rect 30564 39516 30616 39568
rect 28172 39312 28224 39364
rect 28540 39491 28592 39500
rect 28540 39457 28549 39491
rect 28549 39457 28583 39491
rect 28583 39457 28592 39491
rect 28540 39448 28592 39457
rect 29092 39448 29144 39500
rect 28632 39423 28684 39432
rect 28632 39389 28641 39423
rect 28641 39389 28675 39423
rect 28675 39389 28684 39423
rect 28632 39380 28684 39389
rect 29920 39380 29972 39432
rect 29276 39312 29328 39364
rect 29092 39244 29144 39296
rect 30380 39287 30432 39296
rect 30380 39253 30389 39287
rect 30389 39253 30423 39287
rect 30423 39253 30432 39287
rect 30380 39244 30432 39253
rect 6102 39142 6154 39194
rect 6166 39142 6218 39194
rect 6230 39142 6282 39194
rect 6294 39142 6346 39194
rect 6358 39142 6410 39194
rect 16405 39142 16457 39194
rect 16469 39142 16521 39194
rect 16533 39142 16585 39194
rect 16597 39142 16649 39194
rect 16661 39142 16713 39194
rect 26709 39142 26761 39194
rect 26773 39142 26825 39194
rect 26837 39142 26889 39194
rect 26901 39142 26953 39194
rect 26965 39142 27017 39194
rect 5816 39083 5868 39092
rect 5816 39049 5825 39083
rect 5825 39049 5859 39083
rect 5859 39049 5868 39083
rect 5816 39040 5868 39049
rect 6460 39040 6512 39092
rect 6828 39040 6880 39092
rect 7380 39040 7432 39092
rect 8392 39083 8444 39092
rect 8392 39049 8401 39083
rect 8401 39049 8435 39083
rect 8435 39049 8444 39083
rect 8392 39040 8444 39049
rect 9772 39040 9824 39092
rect 15660 39040 15712 39092
rect 18052 39040 18104 39092
rect 5356 38972 5408 39024
rect 6276 38972 6328 39024
rect 9864 39015 9916 39024
rect 9864 38981 9873 39015
rect 9873 38981 9907 39015
rect 9907 38981 9916 39015
rect 9864 38972 9916 38981
rect 1400 38947 1452 38956
rect 1400 38913 1409 38947
rect 1409 38913 1443 38947
rect 1443 38913 1452 38947
rect 1400 38904 1452 38913
rect 8668 38904 8720 38956
rect 13084 38972 13136 39024
rect 15292 39015 15344 39024
rect 15292 38981 15301 39015
rect 15301 38981 15335 39015
rect 15335 38981 15344 39015
rect 15292 38972 15344 38981
rect 12440 38904 12492 38956
rect 3792 38879 3844 38888
rect 1768 38768 1820 38820
rect 2504 38768 2556 38820
rect 3792 38845 3801 38879
rect 3801 38845 3835 38879
rect 3835 38845 3844 38879
rect 3792 38836 3844 38845
rect 4160 38836 4212 38888
rect 7840 38879 7892 38888
rect 3516 38768 3568 38820
rect 4620 38768 4672 38820
rect 5632 38768 5684 38820
rect 7012 38768 7064 38820
rect 7840 38845 7849 38879
rect 7849 38845 7883 38879
rect 7883 38845 7892 38879
rect 7840 38836 7892 38845
rect 8116 38836 8168 38888
rect 8944 38836 8996 38888
rect 10048 38879 10100 38888
rect 10048 38845 10057 38879
rect 10057 38845 10091 38879
rect 10091 38845 10100 38879
rect 10048 38836 10100 38845
rect 13176 38879 13228 38888
rect 9312 38768 9364 38820
rect 9956 38768 10008 38820
rect 11152 38768 11204 38820
rect 2228 38700 2280 38752
rect 11796 38700 11848 38752
rect 13176 38845 13185 38879
rect 13185 38845 13219 38879
rect 13219 38845 13228 38879
rect 13176 38836 13228 38845
rect 13360 38879 13412 38888
rect 13360 38845 13369 38879
rect 13369 38845 13403 38879
rect 13403 38845 13412 38879
rect 15568 38904 15620 38956
rect 16856 38904 16908 38956
rect 17500 38904 17552 38956
rect 19248 39040 19300 39092
rect 20536 39083 20588 39092
rect 20536 39049 20545 39083
rect 20545 39049 20579 39083
rect 20579 39049 20588 39083
rect 20536 39040 20588 39049
rect 22284 39083 22336 39092
rect 22284 39049 22293 39083
rect 22293 39049 22327 39083
rect 22327 39049 22336 39083
rect 22284 39040 22336 39049
rect 23388 39040 23440 39092
rect 25320 39040 25372 39092
rect 25780 39040 25832 39092
rect 26516 39040 26568 39092
rect 27712 39040 27764 39092
rect 29920 39040 29972 39092
rect 31300 39083 31352 39092
rect 31300 39049 31309 39083
rect 31309 39049 31343 39083
rect 31343 39049 31352 39083
rect 31300 39040 31352 39049
rect 19800 38972 19852 39024
rect 20444 38972 20496 39024
rect 13360 38836 13412 38845
rect 15200 38879 15252 38888
rect 13452 38768 13504 38820
rect 15200 38845 15209 38879
rect 15209 38845 15243 38879
rect 15243 38845 15252 38879
rect 15200 38836 15252 38845
rect 15384 38879 15436 38888
rect 15384 38845 15393 38879
rect 15393 38845 15427 38879
rect 15427 38845 15436 38879
rect 15384 38836 15436 38845
rect 15476 38879 15528 38888
rect 15476 38845 15485 38879
rect 15485 38845 15519 38879
rect 15519 38845 15528 38879
rect 20904 38947 20956 38956
rect 15476 38836 15528 38845
rect 15292 38768 15344 38820
rect 16212 38768 16264 38820
rect 17868 38768 17920 38820
rect 16856 38700 16908 38752
rect 18512 38879 18564 38888
rect 18512 38845 18521 38879
rect 18521 38845 18555 38879
rect 18555 38845 18564 38879
rect 18512 38836 18564 38845
rect 19432 38836 19484 38888
rect 19984 38836 20036 38888
rect 20536 38836 20588 38888
rect 20904 38913 20913 38947
rect 20913 38913 20947 38947
rect 20947 38913 20956 38947
rect 20904 38904 20956 38913
rect 21364 38972 21416 39024
rect 24584 38972 24636 39024
rect 25412 38972 25464 39024
rect 23204 38904 23256 38956
rect 23388 38947 23440 38956
rect 23388 38913 23397 38947
rect 23397 38913 23431 38947
rect 23431 38913 23440 38947
rect 23388 38904 23440 38913
rect 23480 38947 23532 38956
rect 23480 38913 23489 38947
rect 23489 38913 23523 38947
rect 23523 38913 23532 38947
rect 23480 38904 23532 38913
rect 24768 38904 24820 38956
rect 28448 38972 28500 39024
rect 30380 38972 30432 39024
rect 31116 38972 31168 39024
rect 27804 38904 27856 38956
rect 21180 38836 21232 38888
rect 22376 38879 22428 38888
rect 20352 38768 20404 38820
rect 22376 38845 22385 38879
rect 22385 38845 22419 38879
rect 22419 38845 22428 38879
rect 22376 38836 22428 38845
rect 23112 38879 23164 38888
rect 23112 38845 23121 38879
rect 23121 38845 23155 38879
rect 23155 38845 23164 38879
rect 23112 38836 23164 38845
rect 23296 38879 23348 38888
rect 23296 38845 23305 38879
rect 23305 38845 23339 38879
rect 23339 38845 23348 38879
rect 23296 38836 23348 38845
rect 23572 38836 23624 38888
rect 26240 38836 26292 38888
rect 26608 38879 26660 38888
rect 26608 38845 26617 38879
rect 26617 38845 26651 38879
rect 26651 38845 26660 38879
rect 26608 38836 26660 38845
rect 27528 38836 27580 38888
rect 27620 38836 27672 38888
rect 27896 38879 27948 38888
rect 27896 38845 27905 38879
rect 27905 38845 27939 38879
rect 27939 38845 27948 38879
rect 27896 38836 27948 38845
rect 27988 38879 28040 38888
rect 27988 38845 27997 38879
rect 27997 38845 28031 38879
rect 28031 38845 28040 38879
rect 28264 38879 28316 38888
rect 27988 38836 28040 38845
rect 28264 38845 28273 38879
rect 28273 38845 28307 38879
rect 28307 38845 28316 38879
rect 28264 38836 28316 38845
rect 30472 38879 30524 38888
rect 30472 38845 30481 38879
rect 30481 38845 30515 38879
rect 30515 38845 30524 38879
rect 30472 38836 30524 38845
rect 31024 38836 31076 38888
rect 19708 38700 19760 38752
rect 20904 38700 20956 38752
rect 22008 38700 22060 38752
rect 22284 38700 22336 38752
rect 23664 38700 23716 38752
rect 23848 38743 23900 38752
rect 23848 38709 23857 38743
rect 23857 38709 23891 38743
rect 23891 38709 23900 38743
rect 23848 38700 23900 38709
rect 24308 38700 24360 38752
rect 25044 38700 25096 38752
rect 25780 38811 25832 38820
rect 25780 38777 25789 38811
rect 25789 38777 25823 38811
rect 25823 38777 25832 38811
rect 25780 38768 25832 38777
rect 26424 38700 26476 38752
rect 28448 38743 28500 38752
rect 28448 38709 28457 38743
rect 28457 38709 28491 38743
rect 28491 38709 28500 38743
rect 28448 38700 28500 38709
rect 30380 38743 30432 38752
rect 30380 38709 30389 38743
rect 30389 38709 30423 38743
rect 30423 38709 30432 38743
rect 30380 38700 30432 38709
rect 11253 38598 11305 38650
rect 11317 38598 11369 38650
rect 11381 38598 11433 38650
rect 11445 38598 11497 38650
rect 11509 38598 11561 38650
rect 21557 38598 21609 38650
rect 21621 38598 21673 38650
rect 21685 38598 21737 38650
rect 21749 38598 21801 38650
rect 21813 38598 21865 38650
rect 1768 38539 1820 38548
rect 1768 38505 1777 38539
rect 1777 38505 1811 38539
rect 1811 38505 1820 38539
rect 1768 38496 1820 38505
rect 1768 38360 1820 38412
rect 2228 38496 2280 38548
rect 2504 38496 2556 38548
rect 2136 38335 2188 38344
rect 2136 38301 2145 38335
rect 2145 38301 2179 38335
rect 2179 38301 2188 38335
rect 2136 38292 2188 38301
rect 2412 38360 2464 38412
rect 3148 38360 3200 38412
rect 3884 38403 3936 38412
rect 3884 38369 3893 38403
rect 3893 38369 3927 38403
rect 3927 38369 3936 38403
rect 3884 38360 3936 38369
rect 4344 38496 4396 38548
rect 7196 38496 7248 38548
rect 7840 38496 7892 38548
rect 4252 38428 4304 38480
rect 6920 38428 6972 38480
rect 8668 38496 8720 38548
rect 9680 38496 9732 38548
rect 11152 38496 11204 38548
rect 5540 38403 5592 38412
rect 2596 38292 2648 38344
rect 5264 38335 5316 38344
rect 4436 38224 4488 38276
rect 4160 38156 4212 38208
rect 5264 38301 5273 38335
rect 5273 38301 5307 38335
rect 5307 38301 5316 38335
rect 5264 38292 5316 38301
rect 5540 38369 5549 38403
rect 5549 38369 5583 38403
rect 5583 38369 5592 38403
rect 5540 38360 5592 38369
rect 5816 38360 5868 38412
rect 6644 38360 6696 38412
rect 9220 38428 9272 38480
rect 12532 38496 12584 38548
rect 13452 38496 13504 38548
rect 14648 38496 14700 38548
rect 17408 38496 17460 38548
rect 9128 38403 9180 38412
rect 9128 38369 9137 38403
rect 9137 38369 9171 38403
rect 9171 38369 9180 38403
rect 9128 38360 9180 38369
rect 5724 38292 5776 38344
rect 8116 38292 8168 38344
rect 8852 38292 8904 38344
rect 9312 38403 9364 38412
rect 9312 38369 9321 38403
rect 9321 38369 9355 38403
rect 9355 38369 9364 38403
rect 10048 38403 10100 38412
rect 9312 38360 9364 38369
rect 10048 38369 10057 38403
rect 10057 38369 10091 38403
rect 10091 38369 10100 38403
rect 10048 38360 10100 38369
rect 10416 38360 10468 38412
rect 10968 38403 11020 38412
rect 10968 38369 10977 38403
rect 10977 38369 11011 38403
rect 11011 38369 11020 38403
rect 10968 38360 11020 38369
rect 4896 38224 4948 38276
rect 5356 38224 5408 38276
rect 4712 38156 4764 38208
rect 9588 38224 9640 38276
rect 11704 38360 11756 38412
rect 7656 38156 7708 38208
rect 10048 38199 10100 38208
rect 10048 38165 10057 38199
rect 10057 38165 10091 38199
rect 10091 38165 10100 38199
rect 10048 38156 10100 38165
rect 12624 38360 12676 38412
rect 16948 38428 17000 38480
rect 17316 38428 17368 38480
rect 16672 38360 16724 38412
rect 17224 38360 17276 38412
rect 17500 38403 17552 38412
rect 17500 38369 17509 38403
rect 17509 38369 17543 38403
rect 17543 38369 17552 38403
rect 17500 38360 17552 38369
rect 17868 38496 17920 38548
rect 18236 38539 18288 38548
rect 18236 38505 18245 38539
rect 18245 38505 18279 38539
rect 18279 38505 18288 38539
rect 18236 38496 18288 38505
rect 19064 38496 19116 38548
rect 20352 38496 20404 38548
rect 22008 38496 22060 38548
rect 18144 38360 18196 38412
rect 18696 38403 18748 38412
rect 18696 38369 18705 38403
rect 18705 38369 18739 38403
rect 18739 38369 18748 38403
rect 18696 38360 18748 38369
rect 12440 38335 12492 38344
rect 12440 38301 12449 38335
rect 12449 38301 12483 38335
rect 12483 38301 12492 38335
rect 12440 38292 12492 38301
rect 13084 38292 13136 38344
rect 17776 38335 17828 38344
rect 16672 38267 16724 38276
rect 16672 38233 16681 38267
rect 16681 38233 16715 38267
rect 16715 38233 16724 38267
rect 16672 38224 16724 38233
rect 17776 38301 17785 38335
rect 17785 38301 17819 38335
rect 17819 38301 17828 38335
rect 17776 38292 17828 38301
rect 16304 38156 16356 38208
rect 16948 38156 17000 38208
rect 22744 38428 22796 38480
rect 23112 38496 23164 38548
rect 24216 38496 24268 38548
rect 24492 38496 24544 38548
rect 23664 38428 23716 38480
rect 23848 38428 23900 38480
rect 20076 38403 20128 38412
rect 20076 38369 20110 38403
rect 20110 38369 20128 38403
rect 20076 38360 20128 38369
rect 22100 38403 22152 38412
rect 22100 38369 22109 38403
rect 22109 38369 22143 38403
rect 22143 38369 22152 38403
rect 27344 38496 27396 38548
rect 25320 38428 25372 38480
rect 26240 38471 26292 38480
rect 26240 38437 26249 38471
rect 26249 38437 26283 38471
rect 26283 38437 26292 38471
rect 26240 38428 26292 38437
rect 27528 38471 27580 38480
rect 27528 38437 27537 38471
rect 27537 38437 27571 38471
rect 27571 38437 27580 38471
rect 27528 38428 27580 38437
rect 22100 38360 22152 38369
rect 25228 38403 25280 38412
rect 25228 38369 25237 38403
rect 25237 38369 25271 38403
rect 25271 38369 25280 38403
rect 25228 38360 25280 38369
rect 26608 38360 26660 38412
rect 19616 38292 19668 38344
rect 24860 38224 24912 38276
rect 21180 38199 21232 38208
rect 21180 38165 21189 38199
rect 21189 38165 21223 38199
rect 21223 38165 21232 38199
rect 21180 38156 21232 38165
rect 22100 38156 22152 38208
rect 23572 38156 23624 38208
rect 23848 38156 23900 38208
rect 24400 38156 24452 38208
rect 24768 38156 24820 38208
rect 27712 38292 27764 38344
rect 28264 38428 28316 38480
rect 28172 38403 28224 38412
rect 28172 38369 28181 38403
rect 28181 38369 28215 38403
rect 28215 38369 28224 38403
rect 28172 38360 28224 38369
rect 30472 38496 30524 38548
rect 31116 38496 31168 38548
rect 28540 38428 28592 38480
rect 27896 38292 27948 38344
rect 28724 38403 28776 38412
rect 28724 38369 28733 38403
rect 28733 38369 28767 38403
rect 28767 38369 28776 38403
rect 28724 38360 28776 38369
rect 28632 38292 28684 38344
rect 29368 38335 29420 38344
rect 25136 38224 25188 38276
rect 25320 38224 25372 38276
rect 26240 38224 26292 38276
rect 29368 38301 29377 38335
rect 29377 38301 29411 38335
rect 29411 38301 29420 38335
rect 29368 38292 29420 38301
rect 25412 38199 25464 38208
rect 25412 38165 25421 38199
rect 25421 38165 25455 38199
rect 25455 38165 25464 38199
rect 25412 38156 25464 38165
rect 27804 38156 27856 38208
rect 28080 38156 28132 38208
rect 28908 38156 28960 38208
rect 30748 38199 30800 38208
rect 30748 38165 30757 38199
rect 30757 38165 30791 38199
rect 30791 38165 30800 38199
rect 30748 38156 30800 38165
rect 6102 38054 6154 38106
rect 6166 38054 6218 38106
rect 6230 38054 6282 38106
rect 6294 38054 6346 38106
rect 6358 38054 6410 38106
rect 16405 38054 16457 38106
rect 16469 38054 16521 38106
rect 16533 38054 16585 38106
rect 16597 38054 16649 38106
rect 16661 38054 16713 38106
rect 26709 38054 26761 38106
rect 26773 38054 26825 38106
rect 26837 38054 26889 38106
rect 26901 38054 26953 38106
rect 26965 38054 27017 38106
rect 5356 37952 5408 38004
rect 7472 37952 7524 38004
rect 9404 37952 9456 38004
rect 9496 37952 9548 38004
rect 15292 37995 15344 38004
rect 3884 37884 3936 37936
rect 15292 37961 15301 37995
rect 15301 37961 15335 37995
rect 15335 37961 15344 37995
rect 15292 37952 15344 37961
rect 4252 37859 4304 37868
rect 4252 37825 4261 37859
rect 4261 37825 4295 37859
rect 4295 37825 4304 37859
rect 4252 37816 4304 37825
rect 5908 37816 5960 37868
rect 11152 37884 11204 37936
rect 11796 37884 11848 37936
rect 11888 37884 11940 37936
rect 12072 37884 12124 37936
rect 12808 37884 12860 37936
rect 13176 37884 13228 37936
rect 15476 37884 15528 37936
rect 12440 37816 12492 37868
rect 12716 37816 12768 37868
rect 15752 37859 15804 37868
rect 15752 37825 15761 37859
rect 15761 37825 15795 37859
rect 15795 37825 15804 37859
rect 15752 37816 15804 37825
rect 2044 37748 2096 37800
rect 3148 37748 3200 37800
rect 4160 37791 4212 37800
rect 4160 37757 4169 37791
rect 4169 37757 4203 37791
rect 4203 37757 4212 37791
rect 4160 37748 4212 37757
rect 4344 37791 4396 37800
rect 4344 37757 4353 37791
rect 4353 37757 4387 37791
rect 4387 37757 4396 37791
rect 4344 37748 4396 37757
rect 4436 37748 4488 37800
rect 6828 37791 6880 37800
rect 6828 37757 6837 37791
rect 6837 37757 6871 37791
rect 6871 37757 6880 37791
rect 6828 37748 6880 37757
rect 7288 37748 7340 37800
rect 7564 37791 7616 37800
rect 7564 37757 7573 37791
rect 7573 37757 7607 37791
rect 7607 37757 7616 37791
rect 7564 37748 7616 37757
rect 8944 37791 8996 37800
rect 8944 37757 8953 37791
rect 8953 37757 8987 37791
rect 8987 37757 8996 37791
rect 8944 37748 8996 37757
rect 10416 37748 10468 37800
rect 2596 37612 2648 37664
rect 7380 37680 7432 37732
rect 10048 37723 10100 37732
rect 10048 37689 10057 37723
rect 10057 37689 10091 37723
rect 10091 37689 10100 37723
rect 10048 37680 10100 37689
rect 11152 37748 11204 37800
rect 11704 37791 11756 37800
rect 11704 37757 11713 37791
rect 11713 37757 11747 37791
rect 11747 37757 11756 37791
rect 11704 37748 11756 37757
rect 11888 37791 11940 37800
rect 11888 37757 11897 37791
rect 11897 37757 11931 37791
rect 11931 37757 11940 37791
rect 11888 37748 11940 37757
rect 12072 37791 12124 37800
rect 12072 37757 12081 37791
rect 12081 37757 12115 37791
rect 12115 37757 12124 37791
rect 12072 37748 12124 37757
rect 12624 37748 12676 37800
rect 12992 37791 13044 37800
rect 12992 37757 13001 37791
rect 13001 37757 13035 37791
rect 13035 37757 13044 37791
rect 12992 37748 13044 37757
rect 13176 37748 13228 37800
rect 14556 37748 14608 37800
rect 15108 37748 15160 37800
rect 15384 37680 15436 37732
rect 15844 37748 15896 37800
rect 15936 37791 15988 37800
rect 15936 37757 15945 37791
rect 15945 37757 15979 37791
rect 15979 37757 15988 37791
rect 18696 37952 18748 38004
rect 20076 37995 20128 38004
rect 20076 37961 20085 37995
rect 20085 37961 20119 37995
rect 20119 37961 20128 37995
rect 20076 37952 20128 37961
rect 20536 37952 20588 38004
rect 22468 37995 22520 38004
rect 17408 37884 17460 37936
rect 17500 37884 17552 37936
rect 15936 37748 15988 37757
rect 16948 37748 17000 37800
rect 17776 37816 17828 37868
rect 20720 37884 20772 37936
rect 22468 37961 22477 37995
rect 22477 37961 22511 37995
rect 22511 37961 22520 37995
rect 22468 37952 22520 37961
rect 23020 37952 23072 38004
rect 25228 37952 25280 38004
rect 26608 37952 26660 38004
rect 27344 37995 27396 38004
rect 27344 37961 27353 37995
rect 27353 37961 27387 37995
rect 27387 37961 27396 37995
rect 27344 37952 27396 37961
rect 27528 37952 27580 38004
rect 31116 37952 31168 38004
rect 19800 37816 19852 37868
rect 18512 37791 18564 37800
rect 3516 37612 3568 37664
rect 3792 37655 3844 37664
rect 3792 37621 3801 37655
rect 3801 37621 3835 37655
rect 3835 37621 3844 37655
rect 3792 37612 3844 37621
rect 4988 37612 5040 37664
rect 5816 37612 5868 37664
rect 6828 37612 6880 37664
rect 7196 37612 7248 37664
rect 10784 37612 10836 37664
rect 10968 37612 11020 37664
rect 11704 37612 11756 37664
rect 12348 37612 12400 37664
rect 12992 37612 13044 37664
rect 14004 37612 14056 37664
rect 15844 37612 15896 37664
rect 16948 37655 17000 37664
rect 16948 37621 16957 37655
rect 16957 37621 16991 37655
rect 16991 37621 17000 37655
rect 16948 37612 17000 37621
rect 18512 37757 18521 37791
rect 18521 37757 18555 37791
rect 18555 37757 18564 37791
rect 18512 37748 18564 37757
rect 19432 37748 19484 37800
rect 19708 37791 19760 37800
rect 17960 37680 18012 37732
rect 19064 37680 19116 37732
rect 19708 37757 19717 37791
rect 19717 37757 19751 37791
rect 19751 37757 19760 37791
rect 19708 37748 19760 37757
rect 21180 37816 21232 37868
rect 25136 37884 25188 37936
rect 27252 37884 27304 37936
rect 21916 37816 21968 37868
rect 22192 37816 22244 37868
rect 23204 37816 23256 37868
rect 24400 37816 24452 37868
rect 21088 37791 21140 37800
rect 21088 37757 21097 37791
rect 21097 37757 21131 37791
rect 21131 37757 21140 37791
rect 21088 37748 21140 37757
rect 22100 37791 22152 37800
rect 22100 37757 22109 37791
rect 22109 37757 22143 37791
rect 22143 37757 22152 37791
rect 23112 37791 23164 37800
rect 22100 37748 22152 37757
rect 23112 37757 23121 37791
rect 23121 37757 23155 37791
rect 23155 37757 23164 37791
rect 23112 37748 23164 37757
rect 23480 37791 23532 37800
rect 19800 37680 19852 37732
rect 21364 37680 21416 37732
rect 23480 37757 23489 37791
rect 23489 37757 23523 37791
rect 23523 37757 23532 37791
rect 23480 37748 23532 37757
rect 23664 37791 23716 37800
rect 23664 37757 23673 37791
rect 23673 37757 23707 37791
rect 23707 37757 23716 37791
rect 23664 37748 23716 37757
rect 24492 37748 24544 37800
rect 25412 37748 25464 37800
rect 26240 37748 26292 37800
rect 27896 37816 27948 37868
rect 17868 37612 17920 37664
rect 20996 37612 21048 37664
rect 23572 37680 23624 37732
rect 23756 37680 23808 37732
rect 25780 37680 25832 37732
rect 26424 37680 26476 37732
rect 27620 37791 27672 37800
rect 27620 37757 27629 37791
rect 27629 37757 27663 37791
rect 27663 37757 27672 37791
rect 27620 37748 27672 37757
rect 28172 37748 28224 37800
rect 29000 37884 29052 37936
rect 29184 37816 29236 37868
rect 29368 37816 29420 37868
rect 28080 37680 28132 37732
rect 28908 37748 28960 37800
rect 30380 37748 30432 37800
rect 27896 37612 27948 37664
rect 28724 37612 28776 37664
rect 29184 37612 29236 37664
rect 11253 37510 11305 37562
rect 11317 37510 11369 37562
rect 11381 37510 11433 37562
rect 11445 37510 11497 37562
rect 11509 37510 11561 37562
rect 21557 37510 21609 37562
rect 21621 37510 21673 37562
rect 21685 37510 21737 37562
rect 21749 37510 21801 37562
rect 21813 37510 21865 37562
rect 3148 37408 3200 37460
rect 5724 37408 5776 37460
rect 7288 37408 7340 37460
rect 8392 37408 8444 37460
rect 9128 37408 9180 37460
rect 9404 37408 9456 37460
rect 3792 37340 3844 37392
rect 2136 37272 2188 37324
rect 2504 37272 2556 37324
rect 3884 37315 3936 37324
rect 3884 37281 3893 37315
rect 3893 37281 3927 37315
rect 3927 37281 3936 37315
rect 6460 37340 6512 37392
rect 9956 37408 10008 37460
rect 12624 37408 12676 37460
rect 3884 37272 3936 37281
rect 4712 37315 4764 37324
rect 4712 37281 4746 37315
rect 4746 37281 4764 37315
rect 4712 37272 4764 37281
rect 5264 37272 5316 37324
rect 6644 37315 6696 37324
rect 6644 37281 6653 37315
rect 6653 37281 6687 37315
rect 6687 37281 6696 37315
rect 6644 37272 6696 37281
rect 6920 37315 6972 37324
rect 6920 37281 6954 37315
rect 6954 37281 6972 37315
rect 6920 37272 6972 37281
rect 9772 37272 9824 37324
rect 11060 37340 11112 37392
rect 10876 37272 10928 37324
rect 11152 37272 11204 37324
rect 13084 37340 13136 37392
rect 15476 37340 15528 37392
rect 15936 37408 15988 37460
rect 16304 37408 16356 37460
rect 20996 37451 21048 37460
rect 12348 37315 12400 37324
rect 12348 37281 12382 37315
rect 12382 37281 12400 37315
rect 12348 37272 12400 37281
rect 15660 37272 15712 37324
rect 17040 37340 17092 37392
rect 16856 37315 16908 37324
rect 16856 37281 16865 37315
rect 16865 37281 16899 37315
rect 16899 37281 16908 37315
rect 16856 37272 16908 37281
rect 2228 37068 2280 37120
rect 10600 37068 10652 37120
rect 14096 37111 14148 37120
rect 14096 37077 14105 37111
rect 14105 37077 14139 37111
rect 14139 37077 14148 37111
rect 14096 37068 14148 37077
rect 18236 37272 18288 37324
rect 19616 37315 19668 37324
rect 19616 37281 19625 37315
rect 19625 37281 19659 37315
rect 19659 37281 19668 37315
rect 19616 37272 19668 37281
rect 19892 37315 19944 37324
rect 19892 37281 19926 37315
rect 19926 37281 19944 37315
rect 20996 37417 21005 37451
rect 21005 37417 21039 37451
rect 21039 37417 21048 37451
rect 20996 37408 21048 37417
rect 21088 37408 21140 37460
rect 21916 37408 21968 37460
rect 22192 37451 22244 37460
rect 22192 37417 22201 37451
rect 22201 37417 22235 37451
rect 22235 37417 22244 37451
rect 22192 37408 22244 37417
rect 22468 37408 22520 37460
rect 24492 37408 24544 37460
rect 26424 37451 26476 37460
rect 26424 37417 26433 37451
rect 26433 37417 26467 37451
rect 26467 37417 26476 37451
rect 26424 37408 26476 37417
rect 27620 37408 27672 37460
rect 30564 37408 30616 37460
rect 21180 37340 21232 37392
rect 19892 37272 19944 37281
rect 22100 37315 22152 37324
rect 22100 37281 22109 37315
rect 22109 37281 22143 37315
rect 22143 37281 22152 37315
rect 23296 37340 23348 37392
rect 23848 37383 23900 37392
rect 23848 37349 23857 37383
rect 23857 37349 23891 37383
rect 23891 37349 23900 37383
rect 23848 37340 23900 37349
rect 24860 37340 24912 37392
rect 26240 37340 26292 37392
rect 27252 37340 27304 37392
rect 27344 37340 27396 37392
rect 22100 37272 22152 37281
rect 24492 37272 24544 37324
rect 27620 37315 27672 37324
rect 23020 37204 23072 37256
rect 27068 37204 27120 37256
rect 27620 37281 27629 37315
rect 27629 37281 27663 37315
rect 27663 37281 27672 37315
rect 27620 37272 27672 37281
rect 28080 37272 28132 37324
rect 28172 37272 28224 37324
rect 30748 37272 30800 37324
rect 31116 37315 31168 37324
rect 31116 37281 31125 37315
rect 31125 37281 31159 37315
rect 31159 37281 31168 37315
rect 31116 37272 31168 37281
rect 19064 37179 19116 37188
rect 19064 37145 19073 37179
rect 19073 37145 19107 37179
rect 19107 37145 19116 37179
rect 19064 37136 19116 37145
rect 22376 37179 22428 37188
rect 22376 37145 22385 37179
rect 22385 37145 22419 37179
rect 22419 37145 22428 37179
rect 22376 37136 22428 37145
rect 22928 37136 22980 37188
rect 18328 37068 18380 37120
rect 22744 37068 22796 37120
rect 23204 37111 23256 37120
rect 23204 37077 23213 37111
rect 23213 37077 23247 37111
rect 23247 37077 23256 37111
rect 23204 37068 23256 37077
rect 23388 37068 23440 37120
rect 27528 37136 27580 37188
rect 26424 37068 26476 37120
rect 6102 36966 6154 37018
rect 6166 36966 6218 37018
rect 6230 36966 6282 37018
rect 6294 36966 6346 37018
rect 6358 36966 6410 37018
rect 16405 36966 16457 37018
rect 16469 36966 16521 37018
rect 16533 36966 16585 37018
rect 16597 36966 16649 37018
rect 16661 36966 16713 37018
rect 26709 36966 26761 37018
rect 26773 36966 26825 37018
rect 26837 36966 26889 37018
rect 26901 36966 26953 37018
rect 26965 36966 27017 37018
rect 7196 36907 7248 36916
rect 7196 36873 7205 36907
rect 7205 36873 7239 36907
rect 7239 36873 7248 36907
rect 7196 36864 7248 36873
rect 7656 36907 7708 36916
rect 7656 36873 7665 36907
rect 7665 36873 7699 36907
rect 7699 36873 7708 36907
rect 7656 36864 7708 36873
rect 1768 36728 1820 36780
rect 3240 36796 3292 36848
rect 4344 36796 4396 36848
rect 7748 36796 7800 36848
rect 2044 36771 2096 36780
rect 2044 36737 2053 36771
rect 2053 36737 2087 36771
rect 2087 36737 2096 36771
rect 2044 36728 2096 36737
rect 5264 36771 5316 36780
rect 5264 36737 5273 36771
rect 5273 36737 5307 36771
rect 5307 36737 5316 36771
rect 5264 36728 5316 36737
rect 2136 36703 2188 36712
rect 2136 36669 2145 36703
rect 2145 36669 2179 36703
rect 2179 36669 2188 36703
rect 2136 36660 2188 36669
rect 2412 36703 2464 36712
rect 2044 36592 2096 36644
rect 2412 36669 2421 36703
rect 2421 36669 2455 36703
rect 2455 36669 2464 36703
rect 2412 36660 2464 36669
rect 3976 36660 4028 36712
rect 9312 36864 9364 36916
rect 9772 36864 9824 36916
rect 11888 36907 11940 36916
rect 11888 36873 11897 36907
rect 11897 36873 11931 36907
rect 11931 36873 11940 36907
rect 11888 36864 11940 36873
rect 9220 36796 9272 36848
rect 9404 36796 9456 36848
rect 12900 36796 12952 36848
rect 19524 36864 19576 36916
rect 19892 36864 19944 36916
rect 21916 36864 21968 36916
rect 22100 36907 22152 36916
rect 22100 36873 22109 36907
rect 22109 36873 22143 36907
rect 22143 36873 22152 36907
rect 23296 36907 23348 36916
rect 22100 36864 22152 36873
rect 23296 36873 23305 36907
rect 23305 36873 23339 36907
rect 23339 36873 23348 36907
rect 23296 36864 23348 36873
rect 23664 36864 23716 36916
rect 25320 36864 25372 36916
rect 17776 36796 17828 36848
rect 2872 36592 2924 36644
rect 5080 36592 5132 36644
rect 8208 36592 8260 36644
rect 9404 36660 9456 36712
rect 11060 36660 11112 36712
rect 12532 36728 12584 36780
rect 12808 36771 12860 36780
rect 12808 36737 12817 36771
rect 12817 36737 12851 36771
rect 12851 36737 12860 36771
rect 12808 36728 12860 36737
rect 12624 36703 12676 36712
rect 12624 36669 12633 36703
rect 12633 36669 12667 36703
rect 12667 36669 12676 36703
rect 12624 36660 12676 36669
rect 12716 36703 12768 36712
rect 12716 36669 12725 36703
rect 12725 36669 12759 36703
rect 12759 36669 12768 36703
rect 14096 36728 14148 36780
rect 12716 36660 12768 36669
rect 13084 36660 13136 36712
rect 16948 36660 17000 36712
rect 17500 36660 17552 36712
rect 19708 36796 19760 36848
rect 21088 36796 21140 36848
rect 21364 36796 21416 36848
rect 24860 36796 24912 36848
rect 28448 36796 28500 36848
rect 19800 36703 19852 36712
rect 1676 36567 1728 36576
rect 1676 36533 1685 36567
rect 1685 36533 1719 36567
rect 1719 36533 1728 36567
rect 1676 36524 1728 36533
rect 3148 36524 3200 36576
rect 7012 36524 7064 36576
rect 8392 36567 8444 36576
rect 8392 36533 8401 36567
rect 8401 36533 8435 36567
rect 8435 36533 8444 36567
rect 8392 36524 8444 36533
rect 10416 36592 10468 36644
rect 10784 36635 10836 36644
rect 10784 36601 10818 36635
rect 10818 36601 10836 36635
rect 10784 36592 10836 36601
rect 14740 36592 14792 36644
rect 13268 36524 13320 36576
rect 14096 36567 14148 36576
rect 14096 36533 14105 36567
rect 14105 36533 14139 36567
rect 14139 36533 14148 36567
rect 14096 36524 14148 36533
rect 15568 36567 15620 36576
rect 15568 36533 15577 36567
rect 15577 36533 15611 36567
rect 15611 36533 15620 36567
rect 15568 36524 15620 36533
rect 17316 36524 17368 36576
rect 17868 36524 17920 36576
rect 18144 36567 18196 36576
rect 18144 36533 18153 36567
rect 18153 36533 18187 36567
rect 18187 36533 18196 36567
rect 18144 36524 18196 36533
rect 19800 36669 19809 36703
rect 19809 36669 19843 36703
rect 19843 36669 19852 36703
rect 19800 36660 19852 36669
rect 22192 36728 22244 36780
rect 22560 36728 22612 36780
rect 23112 36728 23164 36780
rect 23756 36728 23808 36780
rect 27988 36728 28040 36780
rect 21364 36660 21416 36712
rect 21272 36635 21324 36644
rect 21272 36601 21281 36635
rect 21281 36601 21315 36635
rect 21315 36601 21324 36635
rect 21272 36592 21324 36601
rect 21456 36592 21508 36644
rect 22652 36660 22704 36712
rect 23020 36660 23072 36712
rect 23848 36660 23900 36712
rect 21824 36592 21876 36644
rect 22560 36592 22612 36644
rect 23204 36592 23256 36644
rect 26608 36660 26660 36712
rect 26792 36703 26844 36712
rect 26792 36669 26801 36703
rect 26801 36669 26835 36703
rect 26835 36669 26844 36703
rect 26792 36660 26844 36669
rect 27068 36660 27120 36712
rect 27160 36703 27212 36712
rect 27160 36669 27169 36703
rect 27169 36669 27203 36703
rect 27203 36669 27212 36703
rect 27896 36703 27948 36712
rect 27160 36660 27212 36669
rect 27896 36669 27905 36703
rect 27905 36669 27939 36703
rect 27939 36669 27948 36703
rect 27896 36660 27948 36669
rect 28080 36703 28132 36712
rect 28080 36669 28089 36703
rect 28089 36669 28123 36703
rect 28123 36669 28132 36703
rect 28080 36660 28132 36669
rect 27804 36592 27856 36644
rect 29184 36592 29236 36644
rect 22192 36524 22244 36576
rect 24952 36524 25004 36576
rect 26056 36524 26108 36576
rect 27528 36524 27580 36576
rect 30840 36567 30892 36576
rect 30840 36533 30849 36567
rect 30849 36533 30883 36567
rect 30883 36533 30892 36567
rect 30840 36524 30892 36533
rect 11253 36422 11305 36474
rect 11317 36422 11369 36474
rect 11381 36422 11433 36474
rect 11445 36422 11497 36474
rect 11509 36422 11561 36474
rect 21557 36422 21609 36474
rect 21621 36422 21673 36474
rect 21685 36422 21737 36474
rect 21749 36422 21801 36474
rect 21813 36422 21865 36474
rect 5080 36363 5132 36372
rect 5080 36329 5089 36363
rect 5089 36329 5123 36363
rect 5123 36329 5132 36363
rect 5080 36320 5132 36329
rect 6920 36320 6972 36372
rect 8392 36320 8444 36372
rect 10324 36320 10376 36372
rect 10600 36363 10652 36372
rect 10600 36329 10609 36363
rect 10609 36329 10643 36363
rect 10643 36329 10652 36363
rect 10600 36320 10652 36329
rect 3332 36252 3384 36304
rect 3884 36252 3936 36304
rect 4712 36252 4764 36304
rect 7472 36252 7524 36304
rect 1676 36227 1728 36236
rect 1676 36193 1710 36227
rect 1710 36193 1728 36227
rect 1676 36184 1728 36193
rect 3976 36184 4028 36236
rect 4436 36184 4488 36236
rect 6920 36184 6972 36236
rect 7288 36227 7340 36236
rect 7288 36193 7297 36227
rect 7297 36193 7331 36227
rect 7331 36193 7340 36227
rect 7288 36184 7340 36193
rect 7656 36227 7708 36236
rect 7656 36193 7665 36227
rect 7665 36193 7699 36227
rect 7699 36193 7708 36227
rect 7656 36184 7708 36193
rect 10416 36252 10468 36304
rect 11796 36252 11848 36304
rect 17684 36320 17736 36372
rect 18236 36363 18288 36372
rect 18236 36329 18245 36363
rect 18245 36329 18279 36363
rect 18279 36329 18288 36363
rect 18236 36320 18288 36329
rect 21456 36320 21508 36372
rect 26056 36363 26108 36372
rect 26056 36329 26065 36363
rect 26065 36329 26099 36363
rect 26099 36329 26108 36363
rect 26056 36320 26108 36329
rect 26332 36320 26384 36372
rect 27160 36320 27212 36372
rect 17408 36252 17460 36304
rect 17868 36252 17920 36304
rect 22100 36252 22152 36304
rect 22284 36252 22336 36304
rect 23572 36295 23624 36304
rect 23572 36261 23581 36295
rect 23581 36261 23615 36295
rect 23615 36261 23624 36295
rect 23572 36252 23624 36261
rect 26516 36252 26568 36304
rect 27344 36252 27396 36304
rect 9220 36227 9272 36236
rect 9220 36193 9229 36227
rect 9229 36193 9263 36227
rect 9263 36193 9272 36227
rect 9220 36184 9272 36193
rect 13084 36184 13136 36236
rect 13268 36227 13320 36236
rect 13268 36193 13302 36227
rect 13302 36193 13320 36227
rect 13268 36184 13320 36193
rect 15016 36184 15068 36236
rect 4252 36116 4304 36168
rect 2136 35980 2188 36032
rect 3424 36048 3476 36100
rect 5540 36116 5592 36168
rect 7380 36116 7432 36168
rect 7288 36048 7340 36100
rect 10232 36116 10284 36168
rect 15476 36159 15528 36168
rect 15476 36125 15485 36159
rect 15485 36125 15519 36159
rect 15519 36125 15528 36159
rect 15476 36116 15528 36125
rect 17224 36184 17276 36236
rect 17500 36227 17552 36236
rect 17500 36193 17509 36227
rect 17509 36193 17543 36227
rect 17543 36193 17552 36227
rect 17500 36184 17552 36193
rect 9220 36048 9272 36100
rect 2780 36023 2832 36032
rect 2780 35989 2789 36023
rect 2789 35989 2823 36023
rect 2823 35989 2832 36023
rect 2780 35980 2832 35989
rect 3792 35980 3844 36032
rect 4160 35980 4212 36032
rect 5172 35980 5224 36032
rect 12900 36048 12952 36100
rect 11980 35980 12032 36032
rect 13728 35980 13780 36032
rect 14096 35980 14148 36032
rect 16856 35980 16908 36032
rect 17776 36227 17828 36236
rect 17776 36193 17785 36227
rect 17785 36193 17819 36227
rect 17819 36193 17828 36227
rect 17776 36184 17828 36193
rect 17960 36184 18012 36236
rect 21364 36184 21416 36236
rect 21456 36184 21508 36236
rect 23296 36184 23348 36236
rect 23940 36184 23992 36236
rect 26056 36184 26108 36236
rect 27436 36227 27488 36236
rect 27436 36193 27445 36227
rect 27445 36193 27479 36227
rect 27479 36193 27488 36227
rect 27436 36184 27488 36193
rect 27620 36227 27672 36236
rect 27620 36193 27629 36227
rect 27629 36193 27663 36227
rect 27663 36193 27672 36227
rect 27620 36184 27672 36193
rect 17868 36159 17920 36168
rect 17868 36125 17877 36159
rect 17877 36125 17911 36159
rect 17911 36125 17920 36159
rect 17868 36116 17920 36125
rect 18052 36048 18104 36100
rect 20168 36116 20220 36168
rect 21180 36116 21232 36168
rect 26424 36116 26476 36168
rect 27344 36159 27396 36168
rect 27344 36125 27353 36159
rect 27353 36125 27387 36159
rect 27387 36125 27396 36159
rect 27344 36116 27396 36125
rect 18880 36048 18932 36100
rect 22008 36048 22060 36100
rect 24492 36048 24544 36100
rect 26792 36048 26844 36100
rect 29092 36252 29144 36304
rect 30104 36184 30156 36236
rect 30748 36184 30800 36236
rect 29920 36116 29972 36168
rect 19156 35980 19208 36032
rect 20812 35980 20864 36032
rect 22744 36023 22796 36032
rect 22744 35989 22753 36023
rect 22753 35989 22787 36023
rect 22787 35989 22796 36023
rect 22744 35980 22796 35989
rect 23020 35980 23072 36032
rect 23664 35980 23716 36032
rect 25136 36023 25188 36032
rect 25136 35989 25145 36023
rect 25145 35989 25179 36023
rect 25179 35989 25188 36023
rect 25136 35980 25188 35989
rect 25504 35980 25556 36032
rect 28264 35980 28316 36032
rect 29736 36023 29788 36032
rect 29736 35989 29745 36023
rect 29745 35989 29779 36023
rect 29779 35989 29788 36023
rect 29736 35980 29788 35989
rect 30380 36023 30432 36032
rect 30380 35989 30389 36023
rect 30389 35989 30423 36023
rect 30423 35989 30432 36023
rect 30380 35980 30432 35989
rect 30656 35980 30708 36032
rect 6102 35878 6154 35930
rect 6166 35878 6218 35930
rect 6230 35878 6282 35930
rect 6294 35878 6346 35930
rect 6358 35878 6410 35930
rect 16405 35878 16457 35930
rect 16469 35878 16521 35930
rect 16533 35878 16585 35930
rect 16597 35878 16649 35930
rect 16661 35878 16713 35930
rect 26709 35878 26761 35930
rect 26773 35878 26825 35930
rect 26837 35878 26889 35930
rect 26901 35878 26953 35930
rect 26965 35878 27017 35930
rect 5448 35776 5500 35828
rect 3056 35708 3108 35760
rect 3976 35708 4028 35760
rect 6736 35708 6788 35760
rect 9496 35708 9548 35760
rect 2412 35640 2464 35692
rect 4252 35683 4304 35692
rect 4252 35649 4261 35683
rect 4261 35649 4295 35683
rect 4295 35649 4304 35683
rect 4252 35640 4304 35649
rect 3148 35572 3200 35624
rect 3608 35436 3660 35488
rect 4160 35615 4212 35624
rect 4160 35581 4169 35615
rect 4169 35581 4203 35615
rect 4203 35581 4212 35615
rect 4160 35572 4212 35581
rect 5724 35640 5776 35692
rect 5908 35640 5960 35692
rect 7380 35640 7432 35692
rect 4436 35572 4488 35624
rect 5080 35572 5132 35624
rect 6460 35572 6512 35624
rect 7932 35572 7984 35624
rect 10324 35640 10376 35692
rect 11888 35640 11940 35692
rect 13452 35640 13504 35692
rect 4712 35504 4764 35556
rect 5172 35547 5224 35556
rect 4160 35436 4212 35488
rect 5172 35513 5181 35547
rect 5181 35513 5215 35547
rect 5215 35513 5224 35547
rect 5172 35504 5224 35513
rect 6920 35504 6972 35556
rect 10140 35572 10192 35624
rect 10232 35615 10284 35624
rect 10232 35581 10241 35615
rect 10241 35581 10275 35615
rect 10275 35581 10284 35615
rect 10232 35572 10284 35581
rect 10416 35572 10468 35624
rect 11980 35615 12032 35624
rect 11980 35581 11989 35615
rect 11989 35581 12023 35615
rect 12023 35581 12032 35615
rect 11980 35572 12032 35581
rect 14372 35615 14424 35624
rect 14372 35581 14381 35615
rect 14381 35581 14415 35615
rect 14415 35581 14424 35615
rect 14372 35572 14424 35581
rect 10600 35504 10652 35556
rect 11152 35504 11204 35556
rect 12624 35504 12676 35556
rect 13544 35547 13596 35556
rect 5080 35479 5132 35488
rect 5080 35445 5089 35479
rect 5089 35445 5123 35479
rect 5123 35445 5132 35479
rect 5080 35436 5132 35445
rect 7196 35436 7248 35488
rect 7288 35436 7340 35488
rect 9220 35479 9272 35488
rect 9220 35445 9229 35479
rect 9229 35445 9263 35479
rect 9263 35445 9272 35479
rect 9220 35436 9272 35445
rect 9404 35436 9456 35488
rect 10140 35436 10192 35488
rect 10416 35479 10468 35488
rect 10416 35445 10425 35479
rect 10425 35445 10459 35479
rect 10459 35445 10468 35479
rect 10416 35436 10468 35445
rect 10876 35479 10928 35488
rect 10876 35445 10885 35479
rect 10885 35445 10919 35479
rect 10919 35445 10928 35479
rect 10876 35436 10928 35445
rect 12164 35479 12216 35488
rect 12164 35445 12173 35479
rect 12173 35445 12207 35479
rect 12207 35445 12216 35479
rect 12164 35436 12216 35445
rect 13544 35513 13553 35547
rect 13553 35513 13587 35547
rect 13587 35513 13596 35547
rect 13544 35504 13596 35513
rect 14924 35504 14976 35556
rect 14096 35436 14148 35488
rect 14372 35436 14424 35488
rect 15108 35572 15160 35624
rect 16856 35572 16908 35624
rect 17960 35776 18012 35828
rect 17868 35708 17920 35760
rect 19248 35776 19300 35828
rect 19524 35776 19576 35828
rect 18328 35708 18380 35760
rect 21272 35776 21324 35828
rect 21548 35776 21600 35828
rect 27160 35776 27212 35828
rect 27344 35776 27396 35828
rect 28080 35776 28132 35828
rect 17500 35640 17552 35692
rect 23204 35708 23256 35760
rect 24952 35708 25004 35760
rect 27620 35708 27672 35760
rect 27712 35708 27764 35760
rect 27896 35708 27948 35760
rect 29000 35708 29052 35760
rect 17316 35572 17368 35624
rect 18052 35615 18104 35624
rect 18052 35581 18061 35615
rect 18061 35581 18095 35615
rect 18095 35581 18104 35615
rect 18052 35572 18104 35581
rect 19248 35615 19300 35624
rect 19248 35581 19257 35615
rect 19257 35581 19291 35615
rect 19291 35581 19300 35615
rect 19248 35572 19300 35581
rect 23848 35683 23900 35692
rect 23848 35649 23857 35683
rect 23857 35649 23891 35683
rect 23891 35649 23900 35683
rect 23848 35640 23900 35649
rect 27988 35683 28040 35692
rect 15384 35504 15436 35556
rect 18972 35504 19024 35556
rect 19524 35547 19576 35556
rect 19524 35513 19558 35547
rect 19558 35513 19576 35547
rect 19524 35504 19576 35513
rect 16948 35479 17000 35488
rect 16948 35445 16957 35479
rect 16957 35445 16991 35479
rect 16991 35445 17000 35479
rect 16948 35436 17000 35445
rect 17224 35436 17276 35488
rect 19800 35436 19852 35488
rect 21180 35572 21232 35624
rect 21456 35615 21508 35624
rect 21456 35581 21465 35615
rect 21465 35581 21499 35615
rect 21499 35581 21508 35615
rect 21456 35572 21508 35581
rect 22192 35615 22244 35624
rect 22192 35581 22201 35615
rect 22201 35581 22235 35615
rect 22235 35581 22244 35615
rect 22192 35572 22244 35581
rect 23664 35615 23716 35624
rect 23664 35581 23673 35615
rect 23673 35581 23707 35615
rect 23707 35581 23716 35615
rect 23664 35572 23716 35581
rect 25136 35572 25188 35624
rect 27988 35649 27997 35683
rect 27997 35649 28031 35683
rect 28031 35649 28040 35683
rect 27988 35640 28040 35649
rect 28816 35640 28868 35692
rect 27252 35572 27304 35624
rect 27712 35615 27764 35624
rect 27712 35581 27721 35615
rect 27721 35581 27755 35615
rect 27755 35581 27764 35615
rect 27712 35572 27764 35581
rect 27804 35572 27856 35624
rect 28264 35615 28316 35624
rect 20996 35504 21048 35556
rect 21548 35504 21600 35556
rect 22836 35547 22888 35556
rect 22836 35513 22845 35547
rect 22845 35513 22879 35547
rect 22879 35513 22888 35547
rect 22836 35504 22888 35513
rect 23848 35504 23900 35556
rect 25320 35504 25372 35556
rect 26608 35504 26660 35556
rect 27528 35504 27580 35556
rect 28264 35581 28273 35615
rect 28273 35581 28307 35615
rect 28307 35581 28316 35615
rect 28264 35572 28316 35581
rect 29644 35572 29696 35624
rect 29828 35615 29880 35624
rect 29828 35581 29837 35615
rect 29837 35581 29871 35615
rect 29871 35581 29880 35615
rect 30104 35615 30156 35624
rect 29828 35572 29880 35581
rect 30104 35581 30113 35615
rect 30113 35581 30147 35615
rect 30147 35581 30156 35615
rect 30104 35572 30156 35581
rect 22192 35436 22244 35488
rect 22376 35479 22428 35488
rect 22376 35445 22385 35479
rect 22385 35445 22419 35479
rect 22419 35445 22428 35479
rect 22376 35436 22428 35445
rect 25228 35436 25280 35488
rect 27160 35436 27212 35488
rect 30380 35504 30432 35556
rect 30288 35479 30340 35488
rect 30288 35445 30297 35479
rect 30297 35445 30331 35479
rect 30331 35445 30340 35479
rect 30288 35436 30340 35445
rect 30564 35436 30616 35488
rect 11253 35334 11305 35386
rect 11317 35334 11369 35386
rect 11381 35334 11433 35386
rect 11445 35334 11497 35386
rect 11509 35334 11561 35386
rect 21557 35334 21609 35386
rect 21621 35334 21673 35386
rect 21685 35334 21737 35386
rect 21749 35334 21801 35386
rect 21813 35334 21865 35386
rect 2228 35232 2280 35284
rect 5816 35232 5868 35284
rect 10232 35232 10284 35284
rect 3056 35164 3108 35216
rect 2780 35096 2832 35148
rect 3332 35139 3384 35148
rect 3332 35105 3341 35139
rect 3341 35105 3375 35139
rect 3375 35105 3384 35139
rect 3332 35096 3384 35105
rect 3608 35139 3660 35148
rect 3608 35105 3642 35139
rect 3642 35105 3660 35139
rect 3608 35096 3660 35105
rect 5264 35096 5316 35148
rect 5724 35096 5776 35148
rect 7012 35096 7064 35148
rect 7472 35096 7524 35148
rect 8484 35164 8536 35216
rect 9404 35164 9456 35216
rect 12992 35232 13044 35284
rect 10416 35164 10468 35216
rect 11704 35164 11756 35216
rect 12072 35164 12124 35216
rect 14740 35232 14792 35284
rect 7840 35139 7892 35148
rect 7840 35105 7874 35139
rect 7874 35105 7892 35139
rect 7840 35096 7892 35105
rect 10232 35096 10284 35148
rect 11060 35096 11112 35148
rect 12164 35096 12216 35148
rect 2044 35028 2096 35080
rect 2872 35028 2924 35080
rect 4712 35003 4764 35012
rect 4712 34969 4721 35003
rect 4721 34969 4755 35003
rect 4755 34969 4764 35003
rect 14464 35096 14516 35148
rect 14924 35139 14976 35148
rect 14924 35105 14933 35139
rect 14933 35105 14967 35139
rect 14967 35105 14976 35139
rect 14924 35096 14976 35105
rect 15292 35232 15344 35284
rect 15476 35275 15528 35284
rect 15476 35241 15485 35275
rect 15485 35241 15519 35275
rect 15519 35241 15528 35275
rect 15476 35232 15528 35241
rect 17132 35232 17184 35284
rect 22468 35232 22520 35284
rect 23572 35232 23624 35284
rect 24860 35275 24912 35284
rect 24860 35241 24869 35275
rect 24869 35241 24903 35275
rect 24903 35241 24912 35275
rect 24860 35232 24912 35241
rect 25412 35232 25464 35284
rect 27068 35232 27120 35284
rect 28540 35232 28592 35284
rect 29736 35232 29788 35284
rect 14648 35028 14700 35080
rect 16856 35164 16908 35216
rect 16948 35139 17000 35148
rect 16948 35105 16982 35139
rect 16982 35105 17000 35139
rect 16948 35096 17000 35105
rect 15476 35028 15528 35080
rect 4712 34960 4764 34969
rect 15292 34960 15344 35012
rect 19340 35164 19392 35216
rect 19064 35139 19116 35148
rect 19064 35105 19073 35139
rect 19073 35105 19107 35139
rect 19107 35105 19116 35139
rect 19064 35096 19116 35105
rect 19800 35139 19852 35148
rect 18696 35028 18748 35080
rect 19800 35105 19809 35139
rect 19809 35105 19843 35139
rect 19843 35105 19852 35139
rect 19800 35096 19852 35105
rect 20628 35096 20680 35148
rect 21824 35096 21876 35148
rect 22008 35139 22060 35148
rect 22008 35105 22017 35139
rect 22017 35105 22051 35139
rect 22051 35105 22060 35139
rect 22008 35096 22060 35105
rect 19708 35028 19760 35080
rect 19984 35071 20036 35080
rect 19984 35037 19993 35071
rect 19993 35037 20027 35071
rect 20027 35037 20036 35071
rect 19984 35028 20036 35037
rect 29552 35164 29604 35216
rect 22376 35096 22428 35148
rect 25596 35096 25648 35148
rect 27436 35096 27488 35148
rect 27896 35096 27948 35148
rect 29736 35096 29788 35148
rect 22468 35071 22520 35080
rect 22468 35037 22477 35071
rect 22477 35037 22511 35071
rect 22511 35037 22520 35071
rect 22468 35028 22520 35037
rect 26240 35071 26292 35080
rect 26240 35037 26249 35071
rect 26249 35037 26283 35071
rect 26283 35037 26292 35071
rect 26240 35028 26292 35037
rect 2872 34892 2924 34944
rect 3516 34892 3568 34944
rect 3700 34892 3752 34944
rect 5356 34892 5408 34944
rect 5816 34892 5868 34944
rect 8944 34935 8996 34944
rect 8944 34901 8953 34935
rect 8953 34901 8987 34935
rect 8987 34901 8996 34935
rect 8944 34892 8996 34901
rect 9220 34892 9272 34944
rect 10692 34892 10744 34944
rect 13360 34892 13412 34944
rect 14648 34892 14700 34944
rect 15568 34892 15620 34944
rect 17040 34892 17092 34944
rect 17316 34892 17368 34944
rect 18512 34935 18564 34944
rect 18512 34901 18521 34935
rect 18521 34901 18555 34935
rect 18555 34901 18564 34935
rect 18512 34892 18564 34901
rect 18788 34892 18840 34944
rect 20444 34892 20496 34944
rect 22376 34960 22428 35012
rect 23940 34892 23992 34944
rect 24952 34892 25004 34944
rect 26056 34892 26108 34944
rect 29276 35028 29328 35080
rect 29828 35028 29880 35080
rect 30932 35071 30984 35080
rect 30932 35037 30941 35071
rect 30941 35037 30975 35071
rect 30975 35037 30984 35071
rect 30932 35028 30984 35037
rect 27252 34935 27304 34944
rect 27252 34901 27261 34935
rect 27261 34901 27295 34935
rect 27295 34901 27304 34935
rect 27252 34892 27304 34901
rect 29552 34935 29604 34944
rect 29552 34901 29561 34935
rect 29561 34901 29595 34935
rect 29595 34901 29604 34935
rect 29552 34892 29604 34901
rect 6102 34790 6154 34842
rect 6166 34790 6218 34842
rect 6230 34790 6282 34842
rect 6294 34790 6346 34842
rect 6358 34790 6410 34842
rect 16405 34790 16457 34842
rect 16469 34790 16521 34842
rect 16533 34790 16585 34842
rect 16597 34790 16649 34842
rect 16661 34790 16713 34842
rect 26709 34790 26761 34842
rect 26773 34790 26825 34842
rect 26837 34790 26889 34842
rect 26901 34790 26953 34842
rect 26965 34790 27017 34842
rect 2412 34620 2464 34672
rect 3240 34620 3292 34672
rect 1676 34484 1728 34536
rect 2044 34527 2096 34536
rect 2044 34493 2053 34527
rect 2053 34493 2087 34527
rect 2087 34493 2096 34527
rect 2044 34484 2096 34493
rect 2228 34527 2280 34536
rect 2228 34493 2237 34527
rect 2237 34493 2271 34527
rect 2271 34493 2280 34527
rect 2228 34484 2280 34493
rect 4252 34484 4304 34536
rect 4712 34484 4764 34536
rect 5264 34527 5316 34536
rect 5264 34493 5273 34527
rect 5273 34493 5307 34527
rect 5307 34493 5316 34527
rect 5264 34484 5316 34493
rect 2780 34459 2832 34468
rect 2780 34425 2789 34459
rect 2789 34425 2823 34459
rect 2823 34425 2832 34459
rect 2780 34416 2832 34425
rect 5172 34416 5224 34468
rect 5724 34484 5776 34536
rect 6368 34484 6420 34536
rect 7380 34620 7432 34672
rect 7840 34688 7892 34740
rect 10140 34688 10192 34740
rect 10692 34688 10744 34740
rect 13544 34731 13596 34740
rect 7656 34620 7708 34672
rect 7012 34484 7064 34536
rect 7380 34527 7432 34536
rect 7380 34493 7389 34527
rect 7389 34493 7423 34527
rect 7423 34493 7432 34527
rect 7380 34484 7432 34493
rect 7932 34552 7984 34604
rect 9680 34620 9732 34672
rect 12624 34620 12676 34672
rect 13544 34697 13553 34731
rect 13553 34697 13587 34731
rect 13587 34697 13596 34731
rect 13544 34688 13596 34697
rect 14372 34688 14424 34740
rect 13728 34620 13780 34672
rect 8944 34595 8996 34604
rect 8944 34561 8953 34595
rect 8953 34561 8987 34595
rect 8987 34561 8996 34595
rect 8944 34552 8996 34561
rect 8116 34484 8168 34536
rect 9312 34484 9364 34536
rect 12164 34552 12216 34604
rect 14648 34552 14700 34604
rect 14464 34484 14516 34536
rect 15016 34688 15068 34740
rect 15384 34731 15436 34740
rect 15384 34697 15393 34731
rect 15393 34697 15427 34731
rect 15427 34697 15436 34731
rect 15384 34688 15436 34697
rect 17040 34688 17092 34740
rect 17500 34688 17552 34740
rect 15476 34620 15528 34672
rect 15384 34552 15436 34604
rect 15568 34527 15620 34536
rect 15568 34493 15577 34527
rect 15577 34493 15611 34527
rect 15611 34493 15620 34527
rect 15568 34484 15620 34493
rect 15660 34484 15712 34536
rect 16212 34620 16264 34672
rect 7656 34416 7708 34468
rect 10876 34416 10928 34468
rect 2504 34348 2556 34400
rect 5724 34348 5776 34400
rect 6552 34348 6604 34400
rect 6736 34391 6788 34400
rect 6736 34357 6745 34391
rect 6745 34357 6779 34391
rect 6779 34357 6788 34391
rect 6736 34348 6788 34357
rect 6828 34348 6880 34400
rect 9220 34348 9272 34400
rect 12992 34416 13044 34468
rect 13360 34459 13412 34468
rect 13360 34425 13369 34459
rect 13369 34425 13403 34459
rect 13403 34425 13412 34459
rect 13360 34416 13412 34425
rect 13452 34416 13504 34468
rect 14188 34416 14240 34468
rect 18512 34552 18564 34604
rect 18052 34527 18104 34536
rect 12072 34348 12124 34400
rect 14740 34391 14792 34400
rect 14740 34357 14749 34391
rect 14749 34357 14783 34391
rect 14783 34357 14792 34391
rect 14740 34348 14792 34357
rect 15016 34348 15068 34400
rect 15844 34348 15896 34400
rect 18052 34493 18061 34527
rect 18061 34493 18095 34527
rect 18095 34493 18104 34527
rect 18052 34484 18104 34493
rect 18328 34484 18380 34536
rect 18972 34620 19024 34672
rect 19984 34620 20036 34672
rect 23940 34620 23992 34672
rect 24308 34620 24360 34672
rect 25228 34620 25280 34672
rect 19616 34552 19668 34604
rect 19248 34484 19300 34536
rect 26608 34688 26660 34740
rect 29644 34688 29696 34740
rect 30012 34688 30064 34740
rect 25596 34663 25648 34672
rect 25596 34629 25605 34663
rect 25605 34629 25639 34663
rect 25639 34629 25648 34663
rect 25596 34620 25648 34629
rect 29000 34620 29052 34672
rect 26608 34552 26660 34604
rect 30932 34595 30984 34604
rect 30932 34561 30941 34595
rect 30941 34561 30975 34595
rect 30975 34561 30984 34595
rect 30932 34552 30984 34561
rect 16764 34416 16816 34468
rect 17040 34416 17092 34468
rect 17960 34416 18012 34468
rect 20444 34459 20496 34468
rect 20444 34425 20478 34459
rect 20478 34425 20496 34459
rect 20444 34416 20496 34425
rect 20720 34416 20772 34468
rect 24860 34527 24912 34536
rect 24860 34493 24869 34527
rect 24869 34493 24903 34527
rect 24903 34493 24912 34527
rect 24860 34484 24912 34493
rect 25320 34484 25372 34536
rect 25412 34527 25464 34536
rect 25412 34493 25421 34527
rect 25421 34493 25455 34527
rect 25455 34493 25464 34527
rect 26056 34527 26108 34536
rect 25412 34484 25464 34493
rect 26056 34493 26065 34527
rect 26065 34493 26099 34527
rect 26099 34493 26108 34527
rect 26056 34484 26108 34493
rect 26516 34484 26568 34536
rect 26148 34416 26200 34468
rect 30288 34484 30340 34536
rect 16304 34348 16356 34400
rect 20536 34348 20588 34400
rect 20628 34348 20680 34400
rect 22008 34348 22060 34400
rect 22652 34348 22704 34400
rect 25320 34348 25372 34400
rect 28080 34348 28132 34400
rect 11253 34246 11305 34298
rect 11317 34246 11369 34298
rect 11381 34246 11433 34298
rect 11445 34246 11497 34298
rect 11509 34246 11561 34298
rect 21557 34246 21609 34298
rect 21621 34246 21673 34298
rect 21685 34246 21737 34298
rect 21749 34246 21801 34298
rect 21813 34246 21865 34298
rect 2504 34076 2556 34128
rect 1400 34051 1452 34060
rect 1400 34017 1409 34051
rect 1409 34017 1443 34051
rect 1443 34017 1452 34051
rect 1400 34008 1452 34017
rect 3332 34008 3384 34060
rect 5356 34144 5408 34196
rect 6184 34144 6236 34196
rect 6460 34144 6512 34196
rect 6828 34187 6880 34196
rect 6828 34153 6837 34187
rect 6837 34153 6871 34187
rect 6871 34153 6880 34187
rect 6828 34144 6880 34153
rect 9312 34144 9364 34196
rect 8944 34076 8996 34128
rect 9128 34076 9180 34128
rect 14096 34144 14148 34196
rect 19524 34144 19576 34196
rect 20720 34187 20772 34196
rect 20720 34153 20729 34187
rect 20729 34153 20763 34187
rect 20763 34153 20772 34187
rect 20720 34144 20772 34153
rect 2780 33872 2832 33924
rect 1400 33804 1452 33856
rect 3056 33847 3108 33856
rect 3056 33813 3065 33847
rect 3065 33813 3099 33847
rect 3099 33813 3108 33847
rect 3056 33804 3108 33813
rect 3424 33804 3476 33856
rect 4068 33804 4120 33856
rect 5172 34051 5224 34060
rect 5172 34017 5181 34051
rect 5181 34017 5215 34051
rect 5215 34017 5224 34051
rect 5172 34008 5224 34017
rect 5356 34051 5408 34060
rect 5356 34017 5365 34051
rect 5365 34017 5399 34051
rect 5399 34017 5408 34051
rect 5356 34008 5408 34017
rect 5448 34051 5500 34060
rect 5448 34017 5457 34051
rect 5457 34017 5491 34051
rect 5491 34017 5500 34051
rect 5448 34008 5500 34017
rect 5816 33940 5868 33992
rect 6460 34008 6512 34060
rect 8300 34008 8352 34060
rect 6920 33983 6972 33992
rect 6920 33949 6929 33983
rect 6929 33949 6963 33983
rect 6963 33949 6972 33983
rect 6920 33940 6972 33949
rect 8852 33983 8904 33992
rect 8852 33949 8861 33983
rect 8861 33949 8895 33983
rect 8895 33949 8904 33983
rect 8852 33940 8904 33949
rect 9128 33940 9180 33992
rect 12808 34076 12860 34128
rect 13452 34119 13504 34128
rect 13452 34085 13461 34119
rect 13461 34085 13495 34119
rect 13495 34085 13504 34119
rect 13452 34076 13504 34085
rect 14832 34076 14884 34128
rect 16304 34076 16356 34128
rect 18512 34076 18564 34128
rect 13360 34008 13412 34060
rect 13728 34008 13780 34060
rect 16212 34008 16264 34060
rect 19892 34076 19944 34128
rect 10232 33940 10284 33992
rect 7288 33872 7340 33924
rect 10324 33872 10376 33924
rect 4712 33804 4764 33856
rect 5632 33804 5684 33856
rect 9588 33804 9640 33856
rect 9772 33804 9824 33856
rect 11980 33940 12032 33992
rect 14832 33940 14884 33992
rect 15108 33983 15160 33992
rect 15108 33949 15117 33983
rect 15117 33949 15151 33983
rect 15151 33949 15160 33983
rect 15108 33940 15160 33949
rect 15292 33940 15344 33992
rect 17776 33983 17828 33992
rect 17776 33949 17785 33983
rect 17785 33949 17819 33983
rect 17819 33949 17828 33983
rect 17776 33940 17828 33949
rect 14740 33872 14792 33924
rect 18604 33872 18656 33924
rect 11520 33804 11572 33856
rect 12072 33847 12124 33856
rect 12072 33813 12081 33847
rect 12081 33813 12115 33847
rect 12115 33813 12124 33847
rect 12072 33804 12124 33813
rect 12992 33847 13044 33856
rect 12992 33813 13001 33847
rect 13001 33813 13035 33847
rect 13035 33813 13044 33847
rect 12992 33804 13044 33813
rect 13636 33804 13688 33856
rect 14924 33804 14976 33856
rect 17224 33804 17276 33856
rect 19156 34008 19208 34060
rect 19800 34008 19852 34060
rect 20076 34008 20128 34060
rect 20628 34076 20680 34128
rect 23664 34119 23716 34128
rect 23664 34085 23673 34119
rect 23673 34085 23707 34119
rect 23707 34085 23716 34119
rect 23664 34076 23716 34085
rect 22376 34051 22428 34060
rect 19064 33872 19116 33924
rect 19340 33940 19392 33992
rect 22376 34017 22385 34051
rect 22385 34017 22419 34051
rect 22419 34017 22428 34051
rect 22376 34008 22428 34017
rect 22652 34008 22704 34060
rect 25596 34144 25648 34196
rect 27528 34187 27580 34196
rect 24584 34076 24636 34128
rect 25412 34076 25464 34128
rect 26056 34076 26108 34128
rect 19892 33872 19944 33924
rect 21916 33940 21968 33992
rect 20536 33872 20588 33924
rect 22284 33983 22336 33992
rect 22284 33949 22293 33983
rect 22293 33949 22327 33983
rect 22327 33949 22336 33983
rect 22284 33940 22336 33949
rect 23388 33940 23440 33992
rect 24768 33940 24820 33992
rect 26516 34008 26568 34060
rect 27528 34153 27537 34187
rect 27537 34153 27571 34187
rect 27571 34153 27580 34187
rect 27528 34144 27580 34153
rect 27712 34144 27764 34196
rect 29736 34187 29788 34196
rect 29736 34153 29745 34187
rect 29745 34153 29779 34187
rect 29779 34153 29788 34187
rect 29736 34144 29788 34153
rect 29920 34144 29972 34196
rect 27988 34008 28040 34060
rect 28356 34008 28408 34060
rect 28816 34008 28868 34060
rect 29184 34051 29236 34060
rect 29184 34017 29193 34051
rect 29193 34017 29227 34051
rect 29227 34017 29236 34051
rect 29184 34008 29236 34017
rect 29276 34051 29328 34060
rect 29276 34017 29285 34051
rect 29285 34017 29319 34051
rect 29319 34017 29328 34051
rect 29552 34051 29604 34060
rect 29276 34008 29328 34017
rect 29552 34017 29561 34051
rect 29561 34017 29595 34051
rect 29595 34017 29604 34051
rect 29552 34008 29604 34017
rect 30012 34008 30064 34060
rect 31668 34008 31720 34060
rect 23020 33872 23072 33924
rect 19708 33804 19760 33856
rect 20168 33804 20220 33856
rect 21916 33804 21968 33856
rect 22376 33804 22428 33856
rect 22836 33804 22888 33856
rect 25228 33872 25280 33924
rect 25872 33872 25924 33924
rect 29092 33940 29144 33992
rect 23388 33804 23440 33856
rect 25412 33804 25464 33856
rect 26148 33847 26200 33856
rect 26148 33813 26157 33847
rect 26157 33813 26191 33847
rect 26191 33813 26200 33847
rect 26148 33804 26200 33813
rect 6102 33702 6154 33754
rect 6166 33702 6218 33754
rect 6230 33702 6282 33754
rect 6294 33702 6346 33754
rect 6358 33702 6410 33754
rect 16405 33702 16457 33754
rect 16469 33702 16521 33754
rect 16533 33702 16585 33754
rect 16597 33702 16649 33754
rect 16661 33702 16713 33754
rect 26709 33702 26761 33754
rect 26773 33702 26825 33754
rect 26837 33702 26889 33754
rect 26901 33702 26953 33754
rect 26965 33702 27017 33754
rect 4528 33643 4580 33652
rect 4528 33609 4537 33643
rect 4537 33609 4571 33643
rect 4571 33609 4580 33643
rect 4528 33600 4580 33609
rect 5448 33600 5500 33652
rect 6000 33600 6052 33652
rect 11796 33600 11848 33652
rect 13176 33600 13228 33652
rect 13360 33600 13412 33652
rect 18788 33600 18840 33652
rect 19800 33600 19852 33652
rect 2412 33532 2464 33584
rect 4252 33532 4304 33584
rect 5264 33532 5316 33584
rect 2044 33439 2096 33448
rect 2044 33405 2053 33439
rect 2053 33405 2087 33439
rect 2087 33405 2096 33439
rect 2044 33396 2096 33405
rect 3148 33464 3200 33516
rect 3056 33396 3108 33448
rect 5724 33532 5776 33584
rect 5816 33439 5868 33448
rect 2596 33328 2648 33380
rect 2872 33371 2924 33380
rect 2872 33337 2881 33371
rect 2881 33337 2915 33371
rect 2915 33337 2924 33371
rect 2872 33328 2924 33337
rect 1952 33260 2004 33312
rect 2136 33260 2188 33312
rect 3332 33328 3384 33380
rect 3240 33303 3292 33312
rect 3240 33269 3249 33303
rect 3249 33269 3283 33303
rect 3283 33269 3292 33303
rect 3240 33260 3292 33269
rect 3884 33303 3936 33312
rect 3884 33269 3893 33303
rect 3893 33269 3927 33303
rect 3927 33269 3936 33303
rect 3884 33260 3936 33269
rect 4896 33260 4948 33312
rect 5816 33405 5825 33439
rect 5825 33405 5859 33439
rect 5859 33405 5868 33439
rect 5816 33396 5868 33405
rect 5724 33328 5776 33380
rect 7564 33464 7616 33516
rect 7288 33396 7340 33448
rect 10048 33532 10100 33584
rect 6460 33371 6512 33380
rect 6460 33337 6485 33371
rect 6485 33337 6512 33371
rect 7840 33439 7892 33448
rect 7840 33405 7849 33439
rect 7849 33405 7883 33439
rect 7883 33405 7892 33439
rect 7840 33396 7892 33405
rect 8668 33396 8720 33448
rect 9772 33507 9824 33516
rect 9772 33473 9781 33507
rect 9781 33473 9815 33507
rect 9815 33473 9824 33507
rect 9772 33464 9824 33473
rect 11152 33464 11204 33516
rect 11980 33507 12032 33516
rect 8944 33439 8996 33448
rect 8944 33405 8953 33439
rect 8953 33405 8987 33439
rect 8987 33405 8996 33439
rect 8944 33396 8996 33405
rect 9220 33439 9272 33448
rect 9220 33405 9229 33439
rect 9229 33405 9263 33439
rect 9263 33405 9272 33439
rect 9220 33396 9272 33405
rect 9680 33396 9732 33448
rect 10692 33439 10744 33448
rect 10692 33405 10701 33439
rect 10701 33405 10735 33439
rect 10735 33405 10744 33439
rect 10692 33396 10744 33405
rect 11980 33473 11989 33507
rect 11989 33473 12023 33507
rect 12023 33473 12032 33507
rect 11980 33464 12032 33473
rect 11796 33396 11848 33448
rect 12256 33439 12308 33448
rect 12256 33405 12265 33439
rect 12265 33405 12299 33439
rect 12299 33405 12308 33439
rect 12256 33396 12308 33405
rect 6460 33328 6512 33337
rect 9312 33328 9364 33380
rect 17224 33532 17276 33584
rect 20536 33600 20588 33652
rect 21456 33643 21508 33652
rect 21456 33609 21465 33643
rect 21465 33609 21499 33643
rect 21499 33609 21508 33643
rect 21456 33600 21508 33609
rect 15108 33464 15160 33516
rect 19248 33464 19300 33516
rect 14096 33439 14148 33448
rect 14096 33405 14105 33439
rect 14105 33405 14139 33439
rect 14139 33405 14148 33439
rect 14096 33396 14148 33405
rect 7104 33260 7156 33312
rect 7288 33303 7340 33312
rect 7288 33269 7297 33303
rect 7297 33269 7331 33303
rect 7331 33269 7340 33303
rect 7288 33260 7340 33269
rect 7564 33260 7616 33312
rect 8024 33260 8076 33312
rect 13820 33328 13872 33380
rect 15752 33328 15804 33380
rect 16304 33328 16356 33380
rect 18512 33439 18564 33448
rect 18512 33405 18521 33439
rect 18521 33405 18555 33439
rect 18555 33405 18564 33439
rect 18512 33396 18564 33405
rect 19156 33396 19208 33448
rect 19432 33439 19484 33448
rect 19432 33405 19441 33439
rect 19441 33405 19475 33439
rect 19475 33405 19484 33439
rect 19984 33464 20036 33516
rect 20628 33464 20680 33516
rect 21916 33507 21968 33516
rect 21916 33473 21925 33507
rect 21925 33473 21959 33507
rect 21959 33473 21968 33507
rect 21916 33464 21968 33473
rect 23204 33507 23256 33516
rect 23204 33473 23213 33507
rect 23213 33473 23247 33507
rect 23247 33473 23256 33507
rect 23204 33464 23256 33473
rect 19432 33396 19484 33405
rect 19800 33439 19852 33448
rect 19800 33405 19809 33439
rect 19809 33405 19843 33439
rect 19843 33405 19852 33439
rect 19800 33396 19852 33405
rect 20076 33396 20128 33448
rect 20904 33396 20956 33448
rect 21824 33439 21876 33448
rect 21824 33405 21833 33439
rect 21833 33405 21867 33439
rect 21867 33405 21876 33439
rect 21824 33396 21876 33405
rect 22744 33396 22796 33448
rect 24492 33396 24544 33448
rect 24860 33396 24912 33448
rect 25596 33532 25648 33584
rect 25228 33464 25280 33516
rect 29092 33532 29144 33584
rect 29736 33532 29788 33584
rect 28080 33464 28132 33516
rect 29276 33464 29328 33516
rect 29828 33507 29880 33516
rect 29828 33473 29837 33507
rect 29837 33473 29871 33507
rect 29871 33473 29880 33507
rect 29828 33464 29880 33473
rect 16764 33328 16816 33380
rect 14924 33260 14976 33312
rect 15200 33260 15252 33312
rect 17316 33303 17368 33312
rect 17316 33269 17325 33303
rect 17325 33269 17359 33303
rect 17359 33269 17368 33303
rect 17316 33260 17368 33269
rect 17776 33260 17828 33312
rect 18788 33260 18840 33312
rect 19524 33260 19576 33312
rect 19708 33260 19760 33312
rect 20536 33328 20588 33380
rect 23204 33328 23256 33380
rect 23388 33328 23440 33380
rect 25596 33396 25648 33448
rect 25228 33328 25280 33380
rect 25780 33328 25832 33380
rect 20628 33260 20680 33312
rect 20812 33303 20864 33312
rect 20812 33269 20821 33303
rect 20821 33269 20855 33303
rect 20855 33269 20864 33303
rect 20812 33260 20864 33269
rect 20904 33260 20956 33312
rect 21180 33260 21232 33312
rect 21456 33260 21508 33312
rect 21916 33260 21968 33312
rect 23756 33260 23808 33312
rect 24584 33260 24636 33312
rect 25044 33260 25096 33312
rect 25412 33260 25464 33312
rect 26240 33396 26292 33448
rect 27988 33439 28040 33448
rect 27988 33405 27997 33439
rect 27997 33405 28031 33439
rect 28031 33405 28040 33439
rect 27988 33396 28040 33405
rect 28356 33439 28408 33448
rect 28356 33405 28365 33439
rect 28365 33405 28399 33439
rect 28399 33405 28408 33439
rect 28356 33396 28408 33405
rect 28632 33396 28684 33448
rect 28816 33396 28868 33448
rect 29644 33396 29696 33448
rect 30012 33396 30064 33448
rect 28448 33260 28500 33312
rect 30656 33260 30708 33312
rect 11253 33158 11305 33210
rect 11317 33158 11369 33210
rect 11381 33158 11433 33210
rect 11445 33158 11497 33210
rect 11509 33158 11561 33210
rect 21557 33158 21609 33210
rect 21621 33158 21673 33210
rect 21685 33158 21737 33210
rect 21749 33158 21801 33210
rect 21813 33158 21865 33210
rect 2044 33056 2096 33108
rect 1676 32988 1728 33040
rect 1676 32716 1728 32768
rect 2228 32920 2280 32972
rect 2872 32963 2924 32972
rect 2872 32929 2881 32963
rect 2881 32929 2915 32963
rect 2915 32929 2924 32963
rect 2872 32920 2924 32929
rect 2044 32852 2096 32904
rect 2136 32784 2188 32836
rect 6736 32988 6788 33040
rect 3516 32963 3568 32972
rect 3516 32929 3525 32963
rect 3525 32929 3559 32963
rect 3559 32929 3568 32963
rect 3516 32920 3568 32929
rect 3884 32963 3936 32972
rect 3884 32929 3893 32963
rect 3893 32929 3927 32963
rect 3927 32929 3936 32963
rect 3884 32920 3936 32929
rect 5540 32920 5592 32972
rect 4896 32895 4948 32904
rect 4896 32861 4905 32895
rect 4905 32861 4939 32895
rect 4939 32861 4948 32895
rect 4896 32852 4948 32861
rect 5448 32895 5500 32904
rect 5448 32861 5457 32895
rect 5457 32861 5491 32895
rect 5491 32861 5500 32895
rect 5448 32852 5500 32861
rect 5632 32895 5684 32904
rect 5632 32861 5641 32895
rect 5641 32861 5675 32895
rect 5675 32861 5684 32895
rect 5632 32852 5684 32861
rect 3056 32716 3108 32768
rect 3608 32784 3660 32836
rect 3884 32784 3936 32836
rect 3976 32716 4028 32768
rect 4344 32716 4396 32768
rect 4988 32784 5040 32836
rect 6828 32920 6880 32972
rect 6644 32895 6696 32904
rect 6644 32861 6653 32895
rect 6653 32861 6687 32895
rect 6687 32861 6696 32895
rect 6644 32852 6696 32861
rect 7104 32988 7156 33040
rect 10692 33056 10744 33108
rect 11612 33099 11664 33108
rect 11612 33065 11621 33099
rect 11621 33065 11655 33099
rect 11655 33065 11664 33099
rect 11612 33056 11664 33065
rect 11704 33056 11756 33108
rect 12072 33056 12124 33108
rect 13820 33099 13872 33108
rect 8300 32988 8352 33040
rect 9864 32988 9916 33040
rect 9956 32988 10008 33040
rect 12532 32988 12584 33040
rect 13820 33065 13829 33099
rect 13829 33065 13863 33099
rect 13863 33065 13872 33099
rect 13820 33056 13872 33065
rect 15752 33099 15804 33108
rect 15752 33065 15761 33099
rect 15761 33065 15795 33099
rect 15795 33065 15804 33099
rect 15752 33056 15804 33065
rect 18512 33056 18564 33108
rect 9312 32963 9364 32972
rect 9312 32929 9321 32963
rect 9321 32929 9355 32963
rect 9355 32929 9364 32963
rect 9312 32920 9364 32929
rect 10416 32920 10468 32972
rect 11612 32920 11664 32972
rect 12256 32920 12308 32972
rect 8760 32895 8812 32904
rect 8760 32861 8769 32895
rect 8769 32861 8803 32895
rect 8803 32861 8812 32895
rect 8760 32852 8812 32861
rect 9680 32852 9732 32904
rect 6828 32784 6880 32836
rect 12532 32784 12584 32836
rect 12716 32920 12768 32972
rect 13820 32920 13872 32972
rect 16028 32988 16080 33040
rect 17592 32988 17644 33040
rect 18328 32988 18380 33040
rect 22284 33056 22336 33108
rect 22560 33056 22612 33108
rect 22744 33056 22796 33108
rect 23664 33056 23716 33108
rect 24584 33056 24636 33108
rect 24768 33056 24820 33108
rect 25504 33056 25556 33108
rect 25872 33056 25924 33108
rect 26332 33056 26384 33108
rect 26608 33056 26660 33108
rect 30472 33056 30524 33108
rect 19616 32988 19668 33040
rect 21272 33031 21324 33040
rect 21272 32997 21281 33031
rect 21281 32997 21315 33031
rect 21315 32997 21324 33031
rect 21272 32988 21324 32997
rect 14372 32963 14424 32972
rect 12900 32784 12952 32836
rect 13268 32852 13320 32904
rect 14372 32929 14381 32963
rect 14381 32929 14415 32963
rect 14415 32929 14424 32963
rect 14372 32920 14424 32929
rect 15016 32963 15068 32972
rect 15016 32929 15025 32963
rect 15025 32929 15059 32963
rect 15059 32929 15068 32963
rect 15016 32920 15068 32929
rect 15108 32920 15160 32972
rect 15384 32963 15436 32972
rect 15384 32929 15393 32963
rect 15393 32929 15427 32963
rect 15427 32929 15436 32963
rect 15384 32920 15436 32929
rect 15476 32920 15528 32972
rect 15752 32920 15804 32972
rect 17224 32963 17276 32972
rect 17224 32929 17233 32963
rect 17233 32929 17267 32963
rect 17267 32929 17276 32963
rect 17224 32920 17276 32929
rect 18512 32920 18564 32972
rect 19340 32920 19392 32972
rect 19708 32963 19760 32972
rect 19708 32929 19717 32963
rect 19717 32929 19751 32963
rect 19751 32929 19760 32963
rect 19708 32920 19760 32929
rect 19800 32920 19852 32972
rect 15660 32852 15712 32904
rect 16212 32852 16264 32904
rect 5356 32716 5408 32768
rect 6000 32716 6052 32768
rect 6644 32716 6696 32768
rect 8116 32716 8168 32768
rect 8300 32716 8352 32768
rect 9404 32716 9456 32768
rect 10784 32716 10836 32768
rect 11152 32716 11204 32768
rect 12992 32716 13044 32768
rect 13360 32759 13412 32768
rect 13360 32725 13369 32759
rect 13369 32725 13403 32759
rect 13403 32725 13412 32759
rect 13360 32716 13412 32725
rect 14464 32784 14516 32836
rect 15200 32784 15252 32836
rect 19156 32852 19208 32904
rect 19432 32852 19484 32904
rect 17408 32716 17460 32768
rect 17960 32716 18012 32768
rect 19248 32784 19300 32836
rect 19156 32716 19208 32768
rect 19616 32716 19668 32768
rect 19984 32716 20036 32768
rect 20168 32920 20220 32972
rect 20536 32920 20588 32972
rect 20720 32963 20772 32972
rect 20720 32929 20729 32963
rect 20729 32929 20763 32963
rect 20763 32929 20772 32963
rect 20720 32920 20772 32929
rect 20904 32963 20956 32972
rect 20904 32929 20913 32963
rect 20913 32929 20947 32963
rect 20947 32929 20956 32963
rect 20904 32920 20956 32929
rect 22192 32963 22244 32972
rect 22192 32929 22201 32963
rect 22201 32929 22235 32963
rect 22235 32929 22244 32963
rect 22192 32920 22244 32929
rect 20444 32784 20496 32836
rect 20168 32716 20220 32768
rect 20812 32716 20864 32768
rect 24952 32988 25004 33040
rect 25044 32988 25096 33040
rect 26056 32988 26108 33040
rect 22468 32920 22520 32972
rect 23572 32920 23624 32972
rect 24860 32920 24912 32972
rect 25596 32963 25648 32972
rect 25596 32929 25605 32963
rect 25605 32929 25639 32963
rect 25639 32929 25648 32963
rect 25596 32920 25648 32929
rect 25780 32963 25832 32972
rect 25780 32929 25789 32963
rect 25789 32929 25823 32963
rect 25823 32929 25832 32963
rect 25780 32920 25832 32929
rect 26148 32963 26200 32972
rect 24952 32852 25004 32904
rect 25872 32852 25924 32904
rect 26148 32929 26157 32963
rect 26157 32929 26191 32963
rect 26191 32929 26200 32963
rect 26148 32920 26200 32929
rect 28356 32988 28408 33040
rect 28632 32988 28684 33040
rect 28172 32920 28224 32972
rect 28816 32920 28868 32972
rect 29736 32963 29788 32972
rect 29736 32929 29745 32963
rect 29745 32929 29779 32963
rect 29779 32929 29788 32963
rect 29736 32920 29788 32929
rect 29920 32963 29972 32972
rect 29920 32929 29929 32963
rect 29929 32929 29963 32963
rect 29963 32929 29972 32963
rect 29920 32920 29972 32929
rect 26056 32852 26108 32904
rect 28632 32852 28684 32904
rect 29828 32895 29880 32904
rect 29828 32861 29837 32895
rect 29837 32861 29871 32895
rect 29871 32861 29880 32895
rect 29828 32852 29880 32861
rect 23940 32784 23992 32836
rect 29000 32784 29052 32836
rect 21916 32716 21968 32768
rect 22100 32716 22152 32768
rect 27620 32716 27672 32768
rect 29368 32759 29420 32768
rect 29368 32725 29377 32759
rect 29377 32725 29411 32759
rect 29411 32725 29420 32759
rect 29368 32716 29420 32725
rect 29828 32716 29880 32768
rect 6102 32614 6154 32666
rect 6166 32614 6218 32666
rect 6230 32614 6282 32666
rect 6294 32614 6346 32666
rect 6358 32614 6410 32666
rect 16405 32614 16457 32666
rect 16469 32614 16521 32666
rect 16533 32614 16585 32666
rect 16597 32614 16649 32666
rect 16661 32614 16713 32666
rect 26709 32614 26761 32666
rect 26773 32614 26825 32666
rect 26837 32614 26889 32666
rect 26901 32614 26953 32666
rect 26965 32614 27017 32666
rect 2044 32512 2096 32564
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 2228 32444 2280 32496
rect 2044 32376 2096 32428
rect 2504 32512 2556 32564
rect 3332 32512 3384 32564
rect 4896 32512 4948 32564
rect 5172 32512 5224 32564
rect 2412 32444 2464 32496
rect 3516 32444 3568 32496
rect 5264 32444 5316 32496
rect 3240 32419 3292 32428
rect 3240 32385 3249 32419
rect 3249 32385 3283 32419
rect 3283 32385 3292 32419
rect 3240 32376 3292 32385
rect 3332 32376 3384 32428
rect 6736 32512 6788 32564
rect 7656 32512 7708 32564
rect 9128 32555 9180 32564
rect 9128 32521 9137 32555
rect 9137 32521 9171 32555
rect 9171 32521 9180 32555
rect 9128 32512 9180 32521
rect 9680 32555 9732 32564
rect 9680 32521 9689 32555
rect 9689 32521 9723 32555
rect 9723 32521 9732 32555
rect 9680 32512 9732 32521
rect 6460 32444 6512 32496
rect 7380 32444 7432 32496
rect 8116 32444 8168 32496
rect 6000 32376 6052 32428
rect 1676 32240 1728 32292
rect 2596 32308 2648 32360
rect 2228 32172 2280 32224
rect 2780 32172 2832 32224
rect 3148 32308 3200 32360
rect 3976 32351 4028 32360
rect 3976 32317 3985 32351
rect 3985 32317 4019 32351
rect 4019 32317 4028 32351
rect 3976 32308 4028 32317
rect 3608 32240 3660 32292
rect 4528 32308 4580 32360
rect 5356 32308 5408 32360
rect 6828 32351 6880 32360
rect 6828 32317 6837 32351
rect 6837 32317 6871 32351
rect 6871 32317 6880 32351
rect 6828 32308 6880 32317
rect 7196 32351 7248 32360
rect 7196 32317 7205 32351
rect 7205 32317 7239 32351
rect 7239 32317 7248 32351
rect 7196 32308 7248 32317
rect 8024 32351 8076 32360
rect 8024 32317 8033 32351
rect 8033 32317 8067 32351
rect 8067 32317 8076 32351
rect 8024 32308 8076 32317
rect 8668 32444 8720 32496
rect 10508 32444 10560 32496
rect 11060 32444 11112 32496
rect 10968 32419 11020 32428
rect 10968 32385 10977 32419
rect 10977 32385 11011 32419
rect 11011 32385 11020 32419
rect 10968 32376 11020 32385
rect 14096 32512 14148 32564
rect 14556 32555 14608 32564
rect 14556 32521 14565 32555
rect 14565 32521 14599 32555
rect 14599 32521 14608 32555
rect 14556 32512 14608 32521
rect 14924 32512 14976 32564
rect 15108 32512 15160 32564
rect 12900 32444 12952 32496
rect 15476 32444 15528 32496
rect 15752 32487 15804 32496
rect 15752 32453 15761 32487
rect 15761 32453 15795 32487
rect 15795 32453 15804 32487
rect 16028 32512 16080 32564
rect 17224 32512 17276 32564
rect 17408 32512 17460 32564
rect 18972 32512 19024 32564
rect 19708 32512 19760 32564
rect 15752 32444 15804 32453
rect 16304 32444 16356 32496
rect 16580 32444 16632 32496
rect 13360 32376 13412 32428
rect 5540 32240 5592 32292
rect 6000 32240 6052 32292
rect 6920 32240 6972 32292
rect 4344 32172 4396 32224
rect 5172 32215 5224 32224
rect 5172 32181 5181 32215
rect 5181 32181 5215 32215
rect 5215 32181 5224 32215
rect 5172 32172 5224 32181
rect 7196 32172 7248 32224
rect 7380 32240 7432 32292
rect 9220 32308 9272 32360
rect 9588 32351 9640 32360
rect 9588 32317 9597 32351
rect 9597 32317 9631 32351
rect 9631 32317 9640 32351
rect 9588 32308 9640 32317
rect 10784 32351 10836 32360
rect 10784 32317 10793 32351
rect 10793 32317 10827 32351
rect 10827 32317 10836 32351
rect 10784 32308 10836 32317
rect 10876 32308 10928 32360
rect 11152 32351 11204 32360
rect 11152 32317 11161 32351
rect 11161 32317 11195 32351
rect 11195 32317 11204 32351
rect 11152 32308 11204 32317
rect 12624 32308 12676 32360
rect 14280 32351 14332 32360
rect 14280 32317 14289 32351
rect 14289 32317 14323 32351
rect 14323 32317 14332 32351
rect 14280 32308 14332 32317
rect 14832 32308 14884 32360
rect 16028 32308 16080 32360
rect 16212 32351 16264 32360
rect 16212 32317 16221 32351
rect 16221 32317 16255 32351
rect 16255 32317 16264 32351
rect 16212 32308 16264 32317
rect 16304 32308 16356 32360
rect 16580 32351 16632 32360
rect 16580 32317 16589 32351
rect 16589 32317 16623 32351
rect 16623 32317 16632 32351
rect 16580 32308 16632 32317
rect 8024 32172 8076 32224
rect 9864 32240 9916 32292
rect 8208 32172 8260 32224
rect 8300 32172 8352 32224
rect 10600 32215 10652 32224
rect 10600 32181 10609 32215
rect 10609 32181 10643 32215
rect 10643 32181 10652 32215
rect 10600 32172 10652 32181
rect 11888 32240 11940 32292
rect 15292 32240 15344 32292
rect 16488 32240 16540 32292
rect 16764 32351 16816 32360
rect 16764 32317 16773 32351
rect 16773 32317 16807 32351
rect 16807 32317 16816 32351
rect 17316 32376 17368 32428
rect 18052 32444 18104 32496
rect 20168 32444 20220 32496
rect 16764 32308 16816 32317
rect 17224 32308 17276 32360
rect 20076 32376 20128 32428
rect 19708 32351 19760 32360
rect 19708 32317 19717 32351
rect 19717 32317 19751 32351
rect 19751 32317 19760 32351
rect 19708 32308 19760 32317
rect 20628 32444 20680 32496
rect 20444 32419 20496 32428
rect 20444 32385 20453 32419
rect 20453 32385 20487 32419
rect 20487 32385 20496 32419
rect 20444 32376 20496 32385
rect 22100 32512 22152 32564
rect 22192 32512 22244 32564
rect 23572 32555 23624 32564
rect 23572 32521 23581 32555
rect 23581 32521 23615 32555
rect 23615 32521 23624 32555
rect 23572 32512 23624 32521
rect 26608 32512 26660 32564
rect 27988 32512 28040 32564
rect 29920 32512 29972 32564
rect 21272 32444 21324 32496
rect 25044 32487 25096 32496
rect 23480 32376 23532 32428
rect 25044 32453 25053 32487
rect 25053 32453 25087 32487
rect 25087 32453 25096 32487
rect 25044 32444 25096 32453
rect 30932 32419 30984 32428
rect 17868 32240 17920 32292
rect 17960 32240 18012 32292
rect 19156 32240 19208 32292
rect 20444 32240 20496 32292
rect 20996 32308 21048 32360
rect 21272 32308 21324 32360
rect 20628 32240 20680 32292
rect 21916 32308 21968 32360
rect 23388 32308 23440 32360
rect 23940 32308 23992 32360
rect 24768 32308 24820 32360
rect 25228 32308 25280 32360
rect 25504 32351 25556 32360
rect 25504 32317 25513 32351
rect 25513 32317 25547 32351
rect 25547 32317 25556 32351
rect 25504 32308 25556 32317
rect 16948 32172 17000 32224
rect 17316 32172 17368 32224
rect 18328 32172 18380 32224
rect 18788 32172 18840 32224
rect 18972 32172 19024 32224
rect 22008 32172 22060 32224
rect 22284 32172 22336 32224
rect 23020 32172 23072 32224
rect 23756 32172 23808 32224
rect 24860 32283 24912 32292
rect 24860 32249 24885 32283
rect 24885 32249 24912 32283
rect 30932 32385 30941 32419
rect 30941 32385 30975 32419
rect 30975 32385 30984 32419
rect 30932 32376 30984 32385
rect 26148 32308 26200 32360
rect 28448 32351 28500 32360
rect 28448 32317 28466 32351
rect 28466 32317 28500 32351
rect 28448 32308 28500 32317
rect 30380 32308 30432 32360
rect 24860 32240 24912 32249
rect 27528 32240 27580 32292
rect 27988 32240 28040 32292
rect 29092 32240 29144 32292
rect 30656 32283 30708 32292
rect 30656 32249 30674 32283
rect 30674 32249 30708 32283
rect 30656 32240 30708 32249
rect 25412 32172 25464 32224
rect 25780 32172 25832 32224
rect 25964 32172 26016 32224
rect 26056 32172 26108 32224
rect 11253 32070 11305 32122
rect 11317 32070 11369 32122
rect 11381 32070 11433 32122
rect 11445 32070 11497 32122
rect 11509 32070 11561 32122
rect 21557 32070 21609 32122
rect 21621 32070 21673 32122
rect 21685 32070 21737 32122
rect 21749 32070 21801 32122
rect 21813 32070 21865 32122
rect 2872 31968 2924 32020
rect 3516 31968 3568 32020
rect 2596 31900 2648 31952
rect 3148 31900 3200 31952
rect 4436 31900 4488 31952
rect 5172 31968 5224 32020
rect 5816 31968 5868 32020
rect 6920 31968 6972 32020
rect 8760 31968 8812 32020
rect 10784 31968 10836 32020
rect 11060 31968 11112 32020
rect 11888 32011 11940 32020
rect 11888 31977 11897 32011
rect 11897 31977 11931 32011
rect 11931 31977 11940 32011
rect 11888 31968 11940 31977
rect 13176 31968 13228 32020
rect 14280 31968 14332 32020
rect 5540 31900 5592 31952
rect 5724 31900 5776 31952
rect 6736 31900 6788 31952
rect 7840 31900 7892 31952
rect 1676 31832 1728 31884
rect 2228 31875 2280 31884
rect 1952 31807 2004 31816
rect 1952 31773 1961 31807
rect 1961 31773 1995 31807
rect 1995 31773 2004 31807
rect 1952 31764 2004 31773
rect 2228 31841 2237 31875
rect 2237 31841 2271 31875
rect 2271 31841 2280 31875
rect 2228 31832 2280 31841
rect 1308 31696 1360 31748
rect 3332 31764 3384 31816
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 5356 31875 5408 31884
rect 5356 31841 5365 31875
rect 5365 31841 5399 31875
rect 5399 31841 5408 31875
rect 5356 31832 5408 31841
rect 6644 31832 6696 31884
rect 8208 31875 8260 31884
rect 8208 31841 8217 31875
rect 8217 31841 8251 31875
rect 8251 31841 8260 31875
rect 8208 31832 8260 31841
rect 8944 31900 8996 31952
rect 10600 31900 10652 31952
rect 4252 31764 4304 31816
rect 4712 31764 4764 31816
rect 5448 31764 5500 31816
rect 7564 31807 7616 31816
rect 7564 31773 7573 31807
rect 7573 31773 7607 31807
rect 7607 31773 7616 31807
rect 7564 31764 7616 31773
rect 7656 31764 7708 31816
rect 8300 31764 8352 31816
rect 10324 31832 10376 31884
rect 11152 31832 11204 31884
rect 13820 31900 13872 31952
rect 9496 31764 9548 31816
rect 10692 31764 10744 31816
rect 10968 31764 11020 31816
rect 11704 31764 11756 31816
rect 6460 31696 6512 31748
rect 9220 31696 9272 31748
rect 1584 31628 1636 31680
rect 2320 31628 2372 31680
rect 2964 31628 3016 31680
rect 4160 31628 4212 31680
rect 4712 31671 4764 31680
rect 4712 31637 4721 31671
rect 4721 31637 4755 31671
rect 4755 31637 4764 31671
rect 4712 31628 4764 31637
rect 4988 31628 5040 31680
rect 5448 31671 5500 31680
rect 5448 31637 5457 31671
rect 5457 31637 5491 31671
rect 5491 31637 5500 31671
rect 5448 31628 5500 31637
rect 6644 31628 6696 31680
rect 8116 31628 8168 31680
rect 8484 31628 8536 31680
rect 12164 31628 12216 31680
rect 12624 31875 12676 31884
rect 12624 31841 12633 31875
rect 12633 31841 12667 31875
rect 12667 31841 12676 31875
rect 12624 31832 12676 31841
rect 12900 31832 12952 31884
rect 13360 31832 13412 31884
rect 14924 31832 14976 31884
rect 15384 31875 15436 31884
rect 15384 31841 15393 31875
rect 15393 31841 15427 31875
rect 15427 31841 15436 31875
rect 15384 31832 15436 31841
rect 19800 31968 19852 32020
rect 20536 31968 20588 32020
rect 20720 31968 20772 32020
rect 20996 31968 21048 32020
rect 21916 31968 21968 32020
rect 16488 31900 16540 31952
rect 16580 31900 16632 31952
rect 15844 31832 15896 31884
rect 15108 31764 15160 31816
rect 15660 31764 15712 31816
rect 16120 31832 16172 31884
rect 16764 31832 16816 31884
rect 18604 31900 18656 31952
rect 18788 31900 18840 31952
rect 23204 31968 23256 32020
rect 26240 31968 26292 32020
rect 26608 31968 26660 32020
rect 27528 32011 27580 32020
rect 27528 31977 27537 32011
rect 27537 31977 27571 32011
rect 27571 31977 27580 32011
rect 27528 31968 27580 31977
rect 28816 32011 28868 32020
rect 28816 31977 28825 32011
rect 28825 31977 28859 32011
rect 28859 31977 28868 32011
rect 28816 31968 28868 31977
rect 17500 31875 17552 31884
rect 17500 31841 17509 31875
rect 17509 31841 17543 31875
rect 17543 31841 17552 31875
rect 17500 31832 17552 31841
rect 19708 31832 19760 31884
rect 20168 31832 20220 31884
rect 20628 31875 20680 31884
rect 20628 31841 20637 31875
rect 20637 31841 20671 31875
rect 20671 31841 20680 31875
rect 20628 31832 20680 31841
rect 20996 31875 21048 31884
rect 20996 31841 21005 31875
rect 21005 31841 21039 31875
rect 21039 31841 21048 31875
rect 20996 31832 21048 31841
rect 21180 31875 21232 31884
rect 21180 31841 21189 31875
rect 21189 31841 21223 31875
rect 21223 31841 21232 31875
rect 21180 31832 21232 31841
rect 22008 31832 22060 31884
rect 16028 31764 16080 31816
rect 17224 31807 17276 31816
rect 17224 31773 17233 31807
rect 17233 31773 17267 31807
rect 17267 31773 17276 31807
rect 17224 31764 17276 31773
rect 17408 31764 17460 31816
rect 17960 31764 18012 31816
rect 18972 31764 19024 31816
rect 19892 31764 19944 31816
rect 12992 31696 13044 31748
rect 12716 31628 12768 31680
rect 13452 31671 13504 31680
rect 13452 31637 13461 31671
rect 13461 31637 13495 31671
rect 13495 31637 13504 31671
rect 13452 31628 13504 31637
rect 13544 31628 13596 31680
rect 13912 31628 13964 31680
rect 15016 31671 15068 31680
rect 15016 31637 15025 31671
rect 15025 31637 15059 31671
rect 15059 31637 15068 31671
rect 15016 31628 15068 31637
rect 20444 31671 20496 31680
rect 20444 31637 20453 31671
rect 20453 31637 20487 31671
rect 20487 31637 20496 31671
rect 20444 31628 20496 31637
rect 20628 31696 20680 31748
rect 21180 31696 21232 31748
rect 21916 31696 21968 31748
rect 22008 31696 22060 31748
rect 22560 31832 22612 31884
rect 24492 31900 24544 31952
rect 25504 31900 25556 31952
rect 25228 31832 25280 31884
rect 25412 31832 25464 31884
rect 25780 31875 25832 31884
rect 25780 31841 25789 31875
rect 25789 31841 25823 31875
rect 25823 31841 25832 31875
rect 25780 31832 25832 31841
rect 25964 31875 26016 31884
rect 25964 31841 25973 31875
rect 25973 31841 26007 31875
rect 26007 31841 26016 31875
rect 25964 31832 26016 31841
rect 29368 31900 29420 31952
rect 25504 31764 25556 31816
rect 26332 31764 26384 31816
rect 26516 31764 26568 31816
rect 25228 31696 25280 31748
rect 25596 31696 25648 31748
rect 29644 31832 29696 31884
rect 30380 31832 30432 31884
rect 31484 31832 31536 31884
rect 23940 31628 23992 31680
rect 24492 31628 24544 31680
rect 26332 31671 26384 31680
rect 26332 31637 26341 31671
rect 26341 31637 26375 31671
rect 26375 31637 26384 31671
rect 26332 31628 26384 31637
rect 6102 31526 6154 31578
rect 6166 31526 6218 31578
rect 6230 31526 6282 31578
rect 6294 31526 6346 31578
rect 6358 31526 6410 31578
rect 16405 31526 16457 31578
rect 16469 31526 16521 31578
rect 16533 31526 16585 31578
rect 16597 31526 16649 31578
rect 16661 31526 16713 31578
rect 26709 31526 26761 31578
rect 26773 31526 26825 31578
rect 26837 31526 26889 31578
rect 26901 31526 26953 31578
rect 26965 31526 27017 31578
rect 2780 31424 2832 31476
rect 3608 31424 3660 31476
rect 4160 31424 4212 31476
rect 2320 31356 2372 31408
rect 3424 31356 3476 31408
rect 4068 31356 4120 31408
rect 5908 31424 5960 31476
rect 6552 31424 6604 31476
rect 7012 31467 7064 31476
rect 7012 31433 7021 31467
rect 7021 31433 7055 31467
rect 7055 31433 7064 31467
rect 7012 31424 7064 31433
rect 7656 31467 7708 31476
rect 7656 31433 7665 31467
rect 7665 31433 7699 31467
rect 7699 31433 7708 31467
rect 7656 31424 7708 31433
rect 8024 31424 8076 31476
rect 8944 31424 8996 31476
rect 13176 31467 13228 31476
rect 3240 31331 3292 31340
rect 3240 31297 3249 31331
rect 3249 31297 3283 31331
rect 3283 31297 3292 31331
rect 3240 31288 3292 31297
rect 4436 31288 4488 31340
rect 5448 31288 5500 31340
rect 1584 31220 1636 31272
rect 2964 31263 3016 31272
rect 2964 31229 2973 31263
rect 2973 31229 3007 31263
rect 3007 31229 3016 31263
rect 2964 31220 3016 31229
rect 3056 31263 3108 31272
rect 3056 31229 3065 31263
rect 3065 31229 3099 31263
rect 3099 31229 3108 31263
rect 3056 31220 3108 31229
rect 5080 31220 5132 31272
rect 4252 31152 4304 31204
rect 5448 31152 5500 31204
rect 6552 31220 6604 31272
rect 10968 31356 11020 31408
rect 7840 31288 7892 31340
rect 9128 31288 9180 31340
rect 8668 31220 8720 31272
rect 9404 31220 9456 31272
rect 11060 31220 11112 31272
rect 11612 31356 11664 31408
rect 12532 31399 12584 31408
rect 12532 31365 12541 31399
rect 12541 31365 12575 31399
rect 12575 31365 12584 31399
rect 12532 31356 12584 31365
rect 12164 31288 12216 31340
rect 7012 31152 7064 31204
rect 8484 31152 8536 31204
rect 11704 31263 11756 31272
rect 11704 31229 11713 31263
rect 11713 31229 11747 31263
rect 11747 31229 11756 31263
rect 11704 31220 11756 31229
rect 12440 31220 12492 31272
rect 12624 31220 12676 31272
rect 13176 31433 13185 31467
rect 13185 31433 13219 31467
rect 13219 31433 13228 31467
rect 13176 31424 13228 31433
rect 16764 31356 16816 31408
rect 14280 31220 14332 31272
rect 15108 31263 15160 31272
rect 12992 31152 13044 31204
rect 14740 31152 14792 31204
rect 15108 31229 15117 31263
rect 15117 31229 15151 31263
rect 15151 31229 15160 31263
rect 15108 31220 15160 31229
rect 20168 31424 20220 31476
rect 21640 31424 21692 31476
rect 24860 31424 24912 31476
rect 24952 31424 25004 31476
rect 27620 31424 27672 31476
rect 30840 31424 30892 31476
rect 23388 31399 23440 31408
rect 23388 31365 23397 31399
rect 23397 31365 23431 31399
rect 23431 31365 23440 31399
rect 23388 31356 23440 31365
rect 23940 31356 23992 31408
rect 17500 31220 17552 31272
rect 17684 31220 17736 31272
rect 17868 31220 17920 31272
rect 18880 31288 18932 31340
rect 19248 31288 19300 31340
rect 18144 31220 18196 31272
rect 18512 31220 18564 31272
rect 19708 31263 19760 31272
rect 18972 31152 19024 31204
rect 3608 31084 3660 31136
rect 6460 31084 6512 31136
rect 6736 31084 6788 31136
rect 8300 31084 8352 31136
rect 11612 31084 11664 31136
rect 12348 31084 12400 31136
rect 13176 31084 13228 31136
rect 13544 31084 13596 31136
rect 14372 31127 14424 31136
rect 14372 31093 14381 31127
rect 14381 31093 14415 31127
rect 14415 31093 14424 31127
rect 16948 31127 17000 31136
rect 14372 31084 14424 31093
rect 16948 31093 16957 31127
rect 16957 31093 16991 31127
rect 16991 31093 17000 31127
rect 16948 31084 17000 31093
rect 17316 31084 17368 31136
rect 17500 31084 17552 31136
rect 19708 31229 19717 31263
rect 19717 31229 19751 31263
rect 19751 31229 19760 31263
rect 19708 31220 19760 31229
rect 20444 31263 20496 31272
rect 20444 31229 20478 31263
rect 20478 31229 20496 31263
rect 20444 31220 20496 31229
rect 22008 31263 22060 31272
rect 21640 31152 21692 31204
rect 22008 31229 22017 31263
rect 22017 31229 22051 31263
rect 22051 31229 22060 31263
rect 22008 31220 22060 31229
rect 22284 31263 22336 31272
rect 22284 31229 22318 31263
rect 22318 31229 22336 31263
rect 22284 31220 22336 31229
rect 22744 31220 22796 31272
rect 24952 31331 25004 31340
rect 24952 31297 24961 31331
rect 24961 31297 24995 31331
rect 24995 31297 25004 31331
rect 24952 31288 25004 31297
rect 25596 31288 25648 31340
rect 23388 31152 23440 31204
rect 25044 31152 25096 31204
rect 25412 31220 25464 31272
rect 25504 31220 25556 31272
rect 26332 31288 26384 31340
rect 27344 31288 27396 31340
rect 27528 31288 27580 31340
rect 28264 31288 28316 31340
rect 26148 31220 26200 31272
rect 26608 31263 26660 31272
rect 26608 31229 26617 31263
rect 26617 31229 26651 31263
rect 26651 31229 26660 31263
rect 26608 31220 26660 31229
rect 25596 31152 25648 31204
rect 26240 31152 26292 31204
rect 27252 31220 27304 31272
rect 28080 31220 28132 31272
rect 27436 31152 27488 31204
rect 22284 31084 22336 31136
rect 22652 31084 22704 31136
rect 24584 31127 24636 31136
rect 24584 31093 24593 31127
rect 24593 31093 24627 31127
rect 24627 31093 24636 31127
rect 24584 31084 24636 31093
rect 25504 31084 25556 31136
rect 27068 31084 27120 31136
rect 27620 31127 27672 31136
rect 27620 31093 27629 31127
rect 27629 31093 27663 31127
rect 27663 31093 27672 31127
rect 27620 31084 27672 31093
rect 30196 31127 30248 31136
rect 30196 31093 30205 31127
rect 30205 31093 30239 31127
rect 30239 31093 30248 31127
rect 30196 31084 30248 31093
rect 31024 31084 31076 31136
rect 11253 30982 11305 31034
rect 11317 30982 11369 31034
rect 11381 30982 11433 31034
rect 11445 30982 11497 31034
rect 11509 30982 11561 31034
rect 21557 30982 21609 31034
rect 21621 30982 21673 31034
rect 21685 30982 21737 31034
rect 21749 30982 21801 31034
rect 21813 30982 21865 31034
rect 2136 30880 2188 30932
rect 3792 30923 3844 30932
rect 3792 30889 3801 30923
rect 3801 30889 3835 30923
rect 3835 30889 3844 30923
rect 3792 30880 3844 30889
rect 5080 30923 5132 30932
rect 5080 30889 5089 30923
rect 5089 30889 5123 30923
rect 5123 30889 5132 30923
rect 5080 30880 5132 30889
rect 7288 30880 7340 30932
rect 7748 30880 7800 30932
rect 8208 30880 8260 30932
rect 8944 30880 8996 30932
rect 14372 30880 14424 30932
rect 16304 30880 16356 30932
rect 2044 30855 2096 30864
rect 2044 30821 2053 30855
rect 2053 30821 2087 30855
rect 2087 30821 2096 30855
rect 2044 30812 2096 30821
rect 1768 30744 1820 30796
rect 2412 30744 2464 30796
rect 4436 30812 4488 30864
rect 3332 30787 3384 30796
rect 3332 30753 3341 30787
rect 3341 30753 3375 30787
rect 3375 30753 3384 30787
rect 3332 30744 3384 30753
rect 2320 30676 2372 30728
rect 3516 30787 3568 30796
rect 3516 30753 3525 30787
rect 3525 30753 3559 30787
rect 3559 30753 3568 30787
rect 3516 30744 3568 30753
rect 4068 30744 4120 30796
rect 4160 30744 4212 30796
rect 4344 30744 4396 30796
rect 4988 30787 5040 30796
rect 4988 30753 4997 30787
rect 4997 30753 5031 30787
rect 5031 30753 5040 30787
rect 4988 30744 5040 30753
rect 7380 30812 7432 30864
rect 13820 30812 13872 30864
rect 14464 30812 14516 30864
rect 15016 30855 15068 30864
rect 15016 30821 15050 30855
rect 15050 30821 15068 30855
rect 15016 30812 15068 30821
rect 5724 30787 5776 30796
rect 5724 30753 5733 30787
rect 5733 30753 5767 30787
rect 5767 30753 5776 30787
rect 5724 30744 5776 30753
rect 6552 30744 6604 30796
rect 8024 30744 8076 30796
rect 11704 30744 11756 30796
rect 12348 30744 12400 30796
rect 14096 30744 14148 30796
rect 14740 30787 14792 30796
rect 14740 30753 14749 30787
rect 14749 30753 14783 30787
rect 14783 30753 14792 30787
rect 14740 30744 14792 30753
rect 18052 30880 18104 30932
rect 22560 30923 22612 30932
rect 22560 30889 22569 30923
rect 22569 30889 22603 30923
rect 22603 30889 22612 30923
rect 22560 30880 22612 30889
rect 16764 30812 16816 30864
rect 18144 30812 18196 30864
rect 19156 30812 19208 30864
rect 21180 30812 21232 30864
rect 21364 30812 21416 30864
rect 4252 30719 4304 30728
rect 4252 30685 4261 30719
rect 4261 30685 4295 30719
rect 4295 30685 4304 30719
rect 4252 30676 4304 30685
rect 5080 30676 5132 30728
rect 12440 30719 12492 30728
rect 5908 30608 5960 30660
rect 2964 30540 3016 30592
rect 5080 30540 5132 30592
rect 5540 30583 5592 30592
rect 5540 30549 5549 30583
rect 5549 30549 5583 30583
rect 5583 30549 5592 30583
rect 5540 30540 5592 30549
rect 12440 30685 12449 30719
rect 12449 30685 12483 30719
rect 12483 30685 12492 30719
rect 12440 30676 12492 30685
rect 13820 30676 13872 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 13084 30608 13136 30660
rect 13544 30608 13596 30660
rect 8392 30540 8444 30592
rect 12164 30540 12216 30592
rect 13360 30540 13412 30592
rect 18052 30744 18104 30796
rect 20628 30744 20680 30796
rect 21824 30787 21876 30796
rect 21824 30753 21833 30787
rect 21833 30753 21867 30787
rect 21867 30753 21876 30787
rect 21824 30744 21876 30753
rect 22284 30744 22336 30796
rect 23480 30787 23532 30796
rect 17684 30676 17736 30728
rect 22100 30719 22152 30728
rect 22100 30685 22109 30719
rect 22109 30685 22143 30719
rect 22143 30685 22152 30719
rect 22100 30676 22152 30685
rect 22192 30719 22244 30728
rect 22192 30685 22201 30719
rect 22201 30685 22235 30719
rect 22235 30685 22244 30719
rect 22192 30676 22244 30685
rect 18420 30608 18472 30660
rect 19432 30608 19484 30660
rect 20720 30608 20772 30660
rect 21916 30608 21968 30660
rect 23480 30753 23489 30787
rect 23489 30753 23523 30787
rect 23523 30753 23532 30787
rect 23480 30744 23532 30753
rect 24492 30744 24544 30796
rect 27620 30880 27672 30932
rect 29092 30880 29144 30932
rect 24860 30812 24912 30864
rect 25412 30744 25464 30796
rect 25688 30744 25740 30796
rect 26148 30744 26200 30796
rect 27252 30787 27304 30796
rect 27252 30753 27261 30787
rect 27261 30753 27295 30787
rect 27295 30753 27304 30787
rect 27252 30744 27304 30753
rect 23388 30719 23440 30728
rect 23388 30685 23397 30719
rect 23397 30685 23431 30719
rect 23431 30685 23440 30719
rect 23388 30676 23440 30685
rect 23756 30676 23808 30728
rect 23296 30608 23348 30660
rect 24216 30608 24268 30660
rect 25596 30676 25648 30728
rect 27344 30719 27396 30728
rect 27344 30685 27353 30719
rect 27353 30685 27387 30719
rect 27387 30685 27396 30719
rect 27344 30676 27396 30685
rect 27620 30787 27672 30796
rect 27620 30753 27629 30787
rect 27629 30753 27663 30787
rect 27663 30753 27672 30787
rect 28264 30812 28316 30864
rect 27620 30744 27672 30753
rect 27712 30676 27764 30728
rect 31024 30676 31076 30728
rect 17316 30540 17368 30592
rect 17960 30540 18012 30592
rect 19248 30540 19300 30592
rect 23112 30540 23164 30592
rect 25320 30540 25372 30592
rect 27436 30608 27488 30660
rect 30196 30608 30248 30660
rect 27804 30583 27856 30592
rect 27804 30549 27813 30583
rect 27813 30549 27847 30583
rect 27847 30549 27856 30583
rect 27804 30540 27856 30549
rect 30564 30583 30616 30592
rect 30564 30549 30573 30583
rect 30573 30549 30607 30583
rect 30607 30549 30616 30583
rect 30564 30540 30616 30549
rect 6102 30438 6154 30490
rect 6166 30438 6218 30490
rect 6230 30438 6282 30490
rect 6294 30438 6346 30490
rect 6358 30438 6410 30490
rect 16405 30438 16457 30490
rect 16469 30438 16521 30490
rect 16533 30438 16585 30490
rect 16597 30438 16649 30490
rect 16661 30438 16713 30490
rect 26709 30438 26761 30490
rect 26773 30438 26825 30490
rect 26837 30438 26889 30490
rect 26901 30438 26953 30490
rect 26965 30438 27017 30490
rect 2044 30336 2096 30388
rect 4344 30336 4396 30388
rect 6644 30336 6696 30388
rect 4252 30268 4304 30320
rect 1952 30175 2004 30184
rect 1952 30141 1961 30175
rect 1961 30141 1995 30175
rect 1995 30141 2004 30175
rect 1952 30132 2004 30141
rect 2688 30200 2740 30252
rect 2504 30132 2556 30184
rect 3332 30200 3384 30252
rect 4528 30243 4580 30252
rect 4528 30209 4537 30243
rect 4537 30209 4571 30243
rect 4571 30209 4580 30243
rect 4528 30200 4580 30209
rect 5356 30268 5408 30320
rect 6184 30268 6236 30320
rect 7288 30268 7340 30320
rect 7840 30336 7892 30388
rect 8024 30379 8076 30388
rect 8024 30345 8033 30379
rect 8033 30345 8067 30379
rect 8067 30345 8076 30379
rect 8024 30336 8076 30345
rect 8668 30336 8720 30388
rect 12440 30336 12492 30388
rect 12900 30336 12952 30388
rect 13360 30336 13412 30388
rect 17592 30336 17644 30388
rect 23112 30336 23164 30388
rect 7472 30268 7524 30320
rect 19064 30268 19116 30320
rect 19984 30268 20036 30320
rect 20076 30268 20128 30320
rect 3516 30132 3568 30184
rect 3792 30132 3844 30184
rect 7932 30200 7984 30252
rect 12164 30243 12216 30252
rect 1676 30039 1728 30048
rect 1676 30005 1685 30039
rect 1685 30005 1719 30039
rect 1719 30005 1728 30039
rect 1676 29996 1728 30005
rect 4160 29996 4212 30048
rect 5540 30132 5592 30184
rect 7012 30132 7064 30184
rect 7104 30132 7156 30184
rect 4896 30064 4948 30116
rect 6276 30107 6328 30116
rect 6276 30073 6287 30107
rect 6287 30073 6328 30107
rect 6276 30064 6328 30073
rect 6460 30107 6512 30116
rect 6460 30073 6469 30107
rect 6469 30073 6503 30107
rect 6503 30073 6512 30107
rect 6460 30064 6512 30073
rect 5264 29996 5316 30048
rect 5356 29996 5408 30048
rect 5724 29996 5776 30048
rect 6092 30039 6144 30048
rect 6092 30005 6101 30039
rect 6101 30005 6135 30039
rect 6135 30005 6144 30039
rect 6092 29996 6144 30005
rect 8208 30132 8260 30184
rect 12164 30209 12173 30243
rect 12173 30209 12207 30243
rect 12207 30209 12216 30243
rect 12164 30200 12216 30209
rect 16580 30200 16632 30252
rect 18972 30200 19024 30252
rect 22192 30200 22244 30252
rect 23204 30268 23256 30320
rect 23940 30268 23992 30320
rect 27712 30336 27764 30388
rect 24216 30268 24268 30320
rect 24768 30268 24820 30320
rect 25596 30268 25648 30320
rect 11152 30132 11204 30184
rect 8668 30064 8720 30116
rect 9404 30064 9456 30116
rect 9496 30064 9548 30116
rect 10508 30064 10560 30116
rect 12900 30132 12952 30184
rect 14740 30132 14792 30184
rect 16672 30132 16724 30184
rect 19248 30132 19300 30184
rect 20352 30132 20404 30184
rect 20720 30132 20772 30184
rect 21272 30175 21324 30184
rect 21272 30141 21281 30175
rect 21281 30141 21315 30175
rect 21315 30141 21324 30175
rect 21272 30132 21324 30141
rect 21824 30132 21876 30184
rect 22468 30175 22520 30184
rect 22468 30141 22477 30175
rect 22477 30141 22511 30175
rect 22511 30141 22520 30175
rect 22468 30132 22520 30141
rect 12532 30064 12584 30116
rect 15016 30064 15068 30116
rect 18604 30064 18656 30116
rect 23296 30132 23348 30184
rect 25320 30132 25372 30184
rect 25688 30175 25740 30184
rect 25688 30141 25697 30175
rect 25697 30141 25731 30175
rect 25731 30141 25740 30175
rect 25688 30132 25740 30141
rect 26148 30132 26200 30184
rect 27344 30132 27396 30184
rect 28080 30311 28132 30320
rect 28080 30277 28089 30311
rect 28089 30277 28123 30311
rect 28123 30277 28132 30311
rect 28080 30268 28132 30277
rect 30380 30268 30432 30320
rect 30656 30268 30708 30320
rect 28448 30200 28500 30252
rect 30564 30200 30616 30252
rect 7564 29996 7616 30048
rect 8116 29996 8168 30048
rect 8300 29996 8352 30048
rect 11888 29996 11940 30048
rect 12716 29996 12768 30048
rect 13452 29996 13504 30048
rect 14832 29996 14884 30048
rect 16120 29996 16172 30048
rect 19340 29996 19392 30048
rect 23204 29996 23256 30048
rect 25596 30064 25648 30116
rect 26976 30107 27028 30116
rect 26976 30073 27010 30107
rect 27010 30073 27028 30107
rect 26976 30064 27028 30073
rect 27160 30064 27212 30116
rect 23664 29996 23716 30048
rect 11253 29894 11305 29946
rect 11317 29894 11369 29946
rect 11381 29894 11433 29946
rect 11445 29894 11497 29946
rect 11509 29894 11561 29946
rect 21557 29894 21609 29946
rect 21621 29894 21673 29946
rect 21685 29894 21737 29946
rect 21749 29894 21801 29946
rect 21813 29894 21865 29946
rect 3240 29792 3292 29844
rect 1216 29724 1268 29776
rect 1584 29656 1636 29708
rect 1952 29656 2004 29708
rect 2780 29724 2832 29776
rect 3240 29699 3292 29708
rect 1768 29588 1820 29640
rect 1952 29520 2004 29572
rect 3240 29665 3249 29699
rect 3249 29665 3283 29699
rect 3283 29665 3292 29699
rect 3240 29656 3292 29665
rect 4068 29699 4120 29708
rect 4068 29665 4077 29699
rect 4077 29665 4111 29699
rect 4111 29665 4120 29699
rect 4068 29656 4120 29665
rect 4344 29792 4396 29844
rect 5356 29724 5408 29776
rect 6276 29792 6328 29844
rect 9496 29792 9548 29844
rect 10324 29792 10376 29844
rect 10600 29792 10652 29844
rect 11152 29792 11204 29844
rect 5908 29724 5960 29776
rect 7840 29724 7892 29776
rect 9588 29724 9640 29776
rect 14556 29792 14608 29844
rect 16120 29792 16172 29844
rect 16948 29792 17000 29844
rect 11796 29724 11848 29776
rect 14280 29724 14332 29776
rect 4252 29699 4304 29708
rect 4252 29665 4261 29699
rect 4261 29665 4295 29699
rect 4295 29665 4304 29699
rect 4252 29656 4304 29665
rect 4344 29588 4396 29640
rect 4068 29520 4120 29572
rect 6092 29656 6144 29708
rect 6184 29588 6236 29640
rect 6552 29656 6604 29708
rect 7564 29699 7616 29708
rect 7564 29665 7573 29699
rect 7573 29665 7607 29699
rect 7607 29665 7616 29699
rect 7564 29656 7616 29665
rect 7656 29656 7708 29708
rect 8668 29656 8720 29708
rect 7472 29588 7524 29640
rect 7932 29631 7984 29640
rect 7932 29597 7941 29631
rect 7941 29597 7975 29631
rect 7975 29597 7984 29631
rect 7932 29588 7984 29597
rect 6736 29520 6788 29572
rect 10508 29656 10560 29708
rect 10600 29656 10652 29708
rect 11336 29656 11388 29708
rect 11704 29699 11756 29708
rect 11704 29665 11713 29699
rect 11713 29665 11747 29699
rect 11747 29665 11756 29699
rect 11704 29656 11756 29665
rect 13084 29699 13136 29708
rect 9404 29631 9456 29640
rect 9404 29597 9413 29631
rect 9413 29597 9447 29631
rect 9447 29597 9456 29631
rect 9404 29588 9456 29597
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 10600 29520 10652 29572
rect 10876 29520 10928 29572
rect 11428 29520 11480 29572
rect 13084 29665 13093 29699
rect 13093 29665 13127 29699
rect 13127 29665 13136 29699
rect 13084 29656 13136 29665
rect 13259 29699 13311 29708
rect 13259 29665 13265 29699
rect 13265 29665 13299 29699
rect 13299 29665 13311 29699
rect 13259 29656 13311 29665
rect 13452 29699 13504 29708
rect 13452 29665 13461 29699
rect 13461 29665 13495 29699
rect 13495 29665 13504 29699
rect 13452 29656 13504 29665
rect 14464 29656 14516 29708
rect 16580 29724 16632 29776
rect 17500 29724 17552 29776
rect 18144 29792 18196 29844
rect 18880 29792 18932 29844
rect 21180 29792 21232 29844
rect 15844 29656 15896 29708
rect 16672 29699 16724 29708
rect 16672 29665 16681 29699
rect 16681 29665 16715 29699
rect 16715 29665 16724 29699
rect 16672 29656 16724 29665
rect 16948 29699 17000 29708
rect 16948 29665 16982 29699
rect 16982 29665 17000 29699
rect 16948 29656 17000 29665
rect 19340 29656 19392 29708
rect 21272 29656 21324 29708
rect 22744 29724 22796 29776
rect 25596 29792 25648 29844
rect 28172 29792 28224 29844
rect 29184 29792 29236 29844
rect 27160 29724 27212 29776
rect 27804 29724 27856 29776
rect 22192 29699 22244 29708
rect 22192 29665 22201 29699
rect 22201 29665 22235 29699
rect 22235 29665 22244 29699
rect 22192 29656 22244 29665
rect 22468 29656 22520 29708
rect 24860 29656 24912 29708
rect 26056 29656 26108 29708
rect 26240 29656 26292 29708
rect 26608 29656 26660 29708
rect 13360 29631 13412 29640
rect 13360 29597 13363 29631
rect 13363 29597 13397 29631
rect 13397 29597 13412 29631
rect 13360 29588 13412 29597
rect 13820 29588 13872 29640
rect 15200 29588 15252 29640
rect 18972 29588 19024 29640
rect 20168 29631 20220 29640
rect 20168 29597 20177 29631
rect 20177 29597 20211 29631
rect 20211 29597 20220 29631
rect 20168 29588 20220 29597
rect 20444 29631 20496 29640
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 22100 29631 22152 29640
rect 20444 29588 20496 29597
rect 22100 29597 22109 29631
rect 22109 29597 22143 29631
rect 22143 29597 22152 29631
rect 22100 29588 22152 29597
rect 22284 29588 22336 29640
rect 27988 29656 28040 29708
rect 30380 29699 30432 29708
rect 30380 29665 30398 29699
rect 30398 29665 30432 29699
rect 30380 29656 30432 29665
rect 30656 29699 30708 29708
rect 30656 29665 30665 29699
rect 30665 29665 30699 29699
rect 30699 29665 30708 29699
rect 30656 29656 30708 29665
rect 12348 29520 12400 29572
rect 13452 29520 13504 29572
rect 3056 29495 3108 29504
rect 3056 29461 3065 29495
rect 3065 29461 3099 29495
rect 3099 29461 3108 29495
rect 3056 29452 3108 29461
rect 3148 29495 3200 29504
rect 3148 29461 3157 29495
rect 3157 29461 3191 29495
rect 3191 29461 3200 29495
rect 3148 29452 3200 29461
rect 3608 29452 3660 29504
rect 5356 29452 5408 29504
rect 5724 29452 5776 29504
rect 7012 29452 7064 29504
rect 8024 29452 8076 29504
rect 8852 29495 8904 29504
rect 8852 29461 8861 29495
rect 8861 29461 8895 29495
rect 8895 29461 8904 29495
rect 8852 29452 8904 29461
rect 12072 29452 12124 29504
rect 13084 29452 13136 29504
rect 13268 29452 13320 29504
rect 15200 29452 15252 29504
rect 20720 29520 20772 29572
rect 17868 29452 17920 29504
rect 21088 29452 21140 29504
rect 21180 29452 21232 29504
rect 23112 29520 23164 29572
rect 22560 29495 22612 29504
rect 22560 29461 22569 29495
rect 22569 29461 22603 29495
rect 22603 29461 22612 29495
rect 22560 29452 22612 29461
rect 26056 29495 26108 29504
rect 26056 29461 26065 29495
rect 26065 29461 26099 29495
rect 26099 29461 26108 29495
rect 26056 29452 26108 29461
rect 27620 29452 27672 29504
rect 28816 29452 28868 29504
rect 6102 29350 6154 29402
rect 6166 29350 6218 29402
rect 6230 29350 6282 29402
rect 6294 29350 6346 29402
rect 6358 29350 6410 29402
rect 16405 29350 16457 29402
rect 16469 29350 16521 29402
rect 16533 29350 16585 29402
rect 16597 29350 16649 29402
rect 16661 29350 16713 29402
rect 26709 29350 26761 29402
rect 26773 29350 26825 29402
rect 26837 29350 26889 29402
rect 26901 29350 26953 29402
rect 26965 29350 27017 29402
rect 1400 29248 1452 29300
rect 1768 29291 1820 29300
rect 1768 29257 1777 29291
rect 1777 29257 1811 29291
rect 1811 29257 1820 29291
rect 1768 29248 1820 29257
rect 3792 29248 3844 29300
rect 4252 29248 4304 29300
rect 4436 29248 4488 29300
rect 2964 29180 3016 29232
rect 2504 29155 2556 29164
rect 2504 29121 2513 29155
rect 2513 29121 2547 29155
rect 2547 29121 2556 29155
rect 2504 29112 2556 29121
rect 2688 29112 2740 29164
rect 4988 29180 5040 29232
rect 3516 29112 3568 29164
rect 3332 29044 3384 29096
rect 3608 29044 3660 29096
rect 4344 29112 4396 29164
rect 4068 29044 4120 29096
rect 5264 29087 5316 29096
rect 5264 29053 5273 29087
rect 5273 29053 5307 29087
rect 5307 29053 5316 29087
rect 5264 29044 5316 29053
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 5724 29180 5776 29232
rect 5816 29180 5868 29232
rect 6092 29180 6144 29232
rect 6644 29248 6696 29300
rect 7196 29180 7248 29232
rect 5908 29087 5960 29096
rect 5908 29053 5917 29087
rect 5917 29053 5951 29087
rect 5951 29053 5960 29087
rect 5908 29044 5960 29053
rect 10324 29248 10376 29300
rect 10508 29291 10560 29300
rect 10508 29257 10517 29291
rect 10517 29257 10551 29291
rect 10551 29257 10560 29291
rect 10508 29248 10560 29257
rect 11428 29248 11480 29300
rect 11704 29291 11756 29300
rect 8392 29155 8444 29164
rect 8392 29121 8401 29155
rect 8401 29121 8435 29155
rect 8435 29121 8444 29155
rect 8392 29112 8444 29121
rect 8852 29044 8904 29096
rect 5816 28976 5868 29028
rect 6000 28976 6052 29028
rect 6552 28976 6604 29028
rect 6920 28976 6972 29028
rect 7196 28976 7248 29028
rect 9680 28976 9732 29028
rect 2688 28951 2740 28960
rect 2688 28917 2697 28951
rect 2697 28917 2731 28951
rect 2731 28917 2740 28951
rect 2688 28908 2740 28917
rect 3792 28908 3844 28960
rect 4160 28908 4212 28960
rect 7840 28908 7892 28960
rect 9496 28908 9548 28960
rect 10600 29112 10652 29164
rect 10876 29087 10928 29096
rect 10876 29053 10885 29087
rect 10885 29053 10919 29087
rect 10919 29053 10928 29087
rect 10876 29044 10928 29053
rect 11060 29087 11112 29096
rect 11060 29053 11069 29087
rect 11069 29053 11103 29087
rect 11103 29053 11112 29087
rect 11060 29044 11112 29053
rect 11704 29257 11713 29291
rect 11713 29257 11747 29291
rect 11747 29257 11756 29291
rect 11704 29248 11756 29257
rect 12532 29291 12584 29300
rect 12532 29257 12541 29291
rect 12541 29257 12575 29291
rect 12575 29257 12584 29291
rect 12532 29248 12584 29257
rect 16304 29248 16356 29300
rect 19340 29291 19392 29300
rect 11888 29180 11940 29232
rect 12072 29180 12124 29232
rect 18420 29223 18472 29232
rect 12348 29112 12400 29164
rect 13360 29112 13412 29164
rect 15108 29112 15160 29164
rect 16120 29112 16172 29164
rect 16856 29112 16908 29164
rect 18420 29189 18429 29223
rect 18429 29189 18463 29223
rect 18463 29189 18472 29223
rect 18420 29180 18472 29189
rect 19340 29257 19349 29291
rect 19349 29257 19383 29291
rect 19383 29257 19392 29291
rect 19340 29248 19392 29257
rect 19800 29291 19852 29300
rect 19800 29257 19809 29291
rect 19809 29257 19843 29291
rect 19843 29257 19852 29291
rect 19800 29248 19852 29257
rect 21180 29248 21232 29300
rect 22100 29291 22152 29300
rect 22100 29257 22109 29291
rect 22109 29257 22143 29291
rect 22143 29257 22152 29291
rect 22100 29248 22152 29257
rect 23296 29248 23348 29300
rect 26240 29248 26292 29300
rect 30656 29248 30708 29300
rect 17684 29155 17736 29164
rect 11336 29044 11388 29096
rect 12716 29087 12768 29096
rect 11152 28976 11204 29028
rect 12716 29053 12725 29087
rect 12725 29053 12759 29087
rect 12759 29053 12768 29087
rect 12716 29044 12768 29053
rect 13176 29044 13228 29096
rect 14280 29087 14332 29096
rect 14280 29053 14289 29087
rect 14289 29053 14323 29087
rect 14323 29053 14332 29087
rect 14280 29044 14332 29053
rect 14464 29087 14516 29096
rect 14464 29053 14473 29087
rect 14473 29053 14507 29087
rect 14507 29053 14516 29087
rect 14464 29044 14516 29053
rect 14832 29087 14884 29096
rect 14832 29053 14841 29087
rect 14841 29053 14875 29087
rect 14875 29053 14884 29087
rect 14832 29044 14884 29053
rect 15016 29087 15068 29096
rect 15016 29053 15025 29087
rect 15025 29053 15059 29087
rect 15059 29053 15068 29087
rect 15016 29044 15068 29053
rect 15568 29087 15620 29096
rect 15568 29053 15577 29087
rect 15577 29053 15611 29087
rect 15611 29053 15620 29087
rect 15568 29044 15620 29053
rect 16672 29044 16724 29096
rect 17040 29044 17092 29096
rect 10968 28908 11020 28960
rect 11060 28908 11112 28960
rect 12256 28908 12308 28960
rect 14096 28976 14148 29028
rect 15844 28976 15896 29028
rect 16304 28951 16356 28960
rect 16304 28917 16313 28951
rect 16313 28917 16347 28951
rect 16347 28917 16356 28951
rect 16304 28908 16356 28917
rect 17684 29121 17693 29155
rect 17693 29121 17727 29155
rect 17727 29121 17736 29155
rect 17684 29112 17736 29121
rect 18972 29112 19024 29164
rect 26148 29112 26200 29164
rect 28172 29155 28224 29164
rect 28172 29121 28181 29155
rect 28181 29121 28215 29155
rect 28215 29121 28224 29155
rect 28172 29112 28224 29121
rect 17500 28976 17552 29028
rect 20168 29044 20220 29096
rect 22008 29044 22060 29096
rect 22192 29044 22244 29096
rect 23204 29087 23256 29096
rect 23204 29053 23222 29087
rect 23222 29053 23256 29087
rect 23204 29044 23256 29053
rect 23388 29044 23440 29096
rect 29000 29112 29052 29164
rect 31208 29112 31260 29164
rect 19984 28976 20036 29028
rect 24584 28976 24636 29028
rect 24860 28976 24912 29028
rect 25320 28976 25372 29028
rect 28632 29044 28684 29096
rect 26516 29019 26568 29028
rect 26516 28985 26550 29019
rect 26550 28985 26568 29019
rect 26516 28976 26568 28985
rect 30288 28976 30340 29028
rect 18512 28908 18564 28960
rect 19892 28908 19944 28960
rect 23204 28908 23256 28960
rect 23388 28908 23440 28960
rect 25044 28908 25096 28960
rect 29092 28908 29144 28960
rect 11253 28806 11305 28858
rect 11317 28806 11369 28858
rect 11381 28806 11433 28858
rect 11445 28806 11497 28858
rect 11509 28806 11561 28858
rect 21557 28806 21609 28858
rect 21621 28806 21673 28858
rect 21685 28806 21737 28858
rect 21749 28806 21801 28858
rect 21813 28806 21865 28858
rect 3884 28704 3936 28756
rect 4068 28704 4120 28756
rect 4344 28704 4396 28756
rect 5908 28704 5960 28756
rect 8852 28704 8904 28756
rect 9220 28704 9272 28756
rect 1952 28611 2004 28620
rect 1952 28577 1961 28611
rect 1961 28577 1995 28611
rect 1995 28577 2004 28611
rect 1952 28568 2004 28577
rect 3056 28611 3108 28620
rect 3056 28577 3065 28611
rect 3065 28577 3099 28611
rect 3099 28577 3108 28611
rect 3056 28568 3108 28577
rect 1676 28543 1728 28552
rect 1676 28509 1685 28543
rect 1685 28509 1719 28543
rect 1719 28509 1728 28543
rect 1676 28500 1728 28509
rect 2320 28432 2372 28484
rect 4160 28636 4212 28688
rect 4988 28636 5040 28688
rect 3332 28611 3384 28620
rect 3332 28577 3341 28611
rect 3341 28577 3375 28611
rect 3375 28577 3384 28611
rect 3332 28568 3384 28577
rect 2412 28364 2464 28416
rect 6460 28568 6512 28620
rect 6828 28611 6880 28620
rect 6828 28577 6837 28611
rect 6837 28577 6871 28611
rect 6871 28577 6880 28611
rect 6828 28568 6880 28577
rect 3884 28500 3936 28552
rect 4712 28500 4764 28552
rect 6920 28500 6972 28552
rect 7932 28568 7984 28620
rect 8576 28568 8628 28620
rect 9680 28568 9732 28620
rect 11060 28704 11112 28756
rect 11888 28704 11940 28756
rect 12992 28704 13044 28756
rect 13176 28704 13228 28756
rect 14280 28704 14332 28756
rect 14464 28704 14516 28756
rect 10600 28636 10652 28688
rect 11152 28636 11204 28688
rect 13268 28679 13320 28688
rect 13268 28645 13302 28679
rect 13302 28645 13320 28679
rect 13268 28636 13320 28645
rect 15936 28636 15988 28688
rect 10968 28611 11020 28620
rect 7196 28500 7248 28552
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 4160 28364 4212 28416
rect 4804 28364 4856 28416
rect 5632 28364 5684 28416
rect 6092 28432 6144 28484
rect 7288 28432 7340 28484
rect 7840 28432 7892 28484
rect 10968 28577 10977 28611
rect 10977 28577 11011 28611
rect 11011 28577 11020 28611
rect 10968 28568 11020 28577
rect 12072 28611 12124 28620
rect 12072 28577 12081 28611
rect 12081 28577 12115 28611
rect 12115 28577 12124 28611
rect 12072 28568 12124 28577
rect 12256 28611 12308 28620
rect 12256 28577 12265 28611
rect 12265 28577 12299 28611
rect 12299 28577 12308 28611
rect 12256 28568 12308 28577
rect 15016 28611 15068 28620
rect 15016 28577 15025 28611
rect 15025 28577 15059 28611
rect 15059 28577 15068 28611
rect 15016 28568 15068 28577
rect 16856 28704 16908 28756
rect 18144 28704 18196 28756
rect 19984 28747 20036 28756
rect 19984 28713 19993 28747
rect 19993 28713 20027 28747
rect 20027 28713 20036 28747
rect 19984 28704 20036 28713
rect 17684 28636 17736 28688
rect 9864 28432 9916 28484
rect 11796 28500 11848 28552
rect 9220 28364 9272 28416
rect 10232 28407 10284 28416
rect 10232 28373 10241 28407
rect 10241 28373 10275 28407
rect 10275 28373 10284 28407
rect 10232 28364 10284 28373
rect 10876 28432 10928 28484
rect 12164 28500 12216 28552
rect 12992 28543 13044 28552
rect 12992 28509 13001 28543
rect 13001 28509 13035 28543
rect 13035 28509 13044 28543
rect 12992 28500 13044 28509
rect 14832 28543 14884 28552
rect 14832 28509 14841 28543
rect 14841 28509 14875 28543
rect 14875 28509 14884 28543
rect 14832 28500 14884 28509
rect 15936 28500 15988 28552
rect 17132 28543 17184 28552
rect 17132 28509 17141 28543
rect 17141 28509 17175 28543
rect 17175 28509 17184 28543
rect 17132 28500 17184 28509
rect 17316 28568 17368 28620
rect 18236 28636 18288 28688
rect 17960 28568 18012 28620
rect 19800 28568 19852 28620
rect 20168 28611 20220 28620
rect 20168 28577 20177 28611
rect 20177 28577 20211 28611
rect 20211 28577 20220 28611
rect 20168 28568 20220 28577
rect 20444 28611 20496 28620
rect 20444 28577 20453 28611
rect 20453 28577 20487 28611
rect 20487 28577 20496 28611
rect 20444 28568 20496 28577
rect 20628 28636 20680 28688
rect 22100 28636 22152 28688
rect 22192 28636 22244 28688
rect 23204 28636 23256 28688
rect 24308 28704 24360 28756
rect 26148 28704 26200 28756
rect 26516 28704 26568 28756
rect 30380 28704 30432 28756
rect 24768 28636 24820 28688
rect 21272 28568 21324 28620
rect 22560 28568 22612 28620
rect 23756 28568 23808 28620
rect 24952 28636 25004 28688
rect 25044 28611 25096 28620
rect 12348 28432 12400 28484
rect 16672 28432 16724 28484
rect 17040 28432 17092 28484
rect 11796 28364 11848 28416
rect 11888 28364 11940 28416
rect 14648 28364 14700 28416
rect 16856 28364 16908 28416
rect 17776 28500 17828 28552
rect 20352 28543 20404 28552
rect 20352 28509 20361 28543
rect 20361 28509 20395 28543
rect 20395 28509 20404 28543
rect 20352 28500 20404 28509
rect 25044 28577 25053 28611
rect 25053 28577 25087 28611
rect 25087 28577 25096 28611
rect 25044 28568 25096 28577
rect 25688 28609 25740 28620
rect 25688 28575 25697 28609
rect 25697 28575 25731 28609
rect 25731 28575 25740 28609
rect 25688 28568 25740 28575
rect 25872 28611 25924 28620
rect 25872 28577 25881 28611
rect 25881 28577 25915 28611
rect 25915 28577 25924 28611
rect 26240 28611 26292 28620
rect 25872 28568 25924 28577
rect 26240 28577 26249 28611
rect 26249 28577 26283 28611
rect 26283 28577 26292 28611
rect 26240 28568 26292 28577
rect 27620 28611 27672 28620
rect 27620 28577 27629 28611
rect 27629 28577 27663 28611
rect 27663 28577 27672 28611
rect 27620 28568 27672 28577
rect 28632 28611 28684 28620
rect 17776 28364 17828 28416
rect 18052 28364 18104 28416
rect 19156 28364 19208 28416
rect 22284 28364 22336 28416
rect 22468 28364 22520 28416
rect 22744 28364 22796 28416
rect 24492 28407 24544 28416
rect 24492 28373 24501 28407
rect 24501 28373 24535 28407
rect 24535 28373 24544 28407
rect 24492 28364 24544 28373
rect 25872 28432 25924 28484
rect 26148 28500 26200 28552
rect 28632 28577 28641 28611
rect 28641 28577 28675 28611
rect 28675 28577 28684 28611
rect 28632 28568 28684 28577
rect 29092 28568 29144 28620
rect 31208 28611 31260 28620
rect 27528 28432 27580 28484
rect 28724 28500 28776 28552
rect 28908 28543 28960 28552
rect 28908 28509 28917 28543
rect 28917 28509 28951 28543
rect 28951 28509 28960 28543
rect 28908 28500 28960 28509
rect 29000 28543 29052 28552
rect 29000 28509 29009 28543
rect 29009 28509 29043 28543
rect 29043 28509 29052 28543
rect 31208 28577 31217 28611
rect 31217 28577 31251 28611
rect 31251 28577 31260 28611
rect 31208 28568 31260 28577
rect 29000 28500 29052 28509
rect 24952 28364 25004 28416
rect 28540 28364 28592 28416
rect 29736 28364 29788 28416
rect 6102 28262 6154 28314
rect 6166 28262 6218 28314
rect 6230 28262 6282 28314
rect 6294 28262 6346 28314
rect 6358 28262 6410 28314
rect 16405 28262 16457 28314
rect 16469 28262 16521 28314
rect 16533 28262 16585 28314
rect 16597 28262 16649 28314
rect 16661 28262 16713 28314
rect 26709 28262 26761 28314
rect 26773 28262 26825 28314
rect 26837 28262 26889 28314
rect 26901 28262 26953 28314
rect 26965 28262 27017 28314
rect 1308 28160 1360 28212
rect 2412 28160 2464 28212
rect 3884 28203 3936 28212
rect 1216 28092 1268 28144
rect 2688 28024 2740 28076
rect 3332 28092 3384 28144
rect 3884 28169 3893 28203
rect 3893 28169 3927 28203
rect 3927 28169 3936 28203
rect 3884 28160 3936 28169
rect 4896 28203 4948 28212
rect 4896 28169 4905 28203
rect 4905 28169 4939 28203
rect 4939 28169 4948 28203
rect 4896 28160 4948 28169
rect 4988 28160 5040 28212
rect 7104 28203 7156 28212
rect 4160 28092 4212 28144
rect 4436 28024 4488 28076
rect 4804 28024 4856 28076
rect 1492 27999 1544 28008
rect 1492 27965 1501 27999
rect 1501 27965 1535 27999
rect 1535 27965 1544 27999
rect 1492 27956 1544 27965
rect 2780 27999 2832 28008
rect 2780 27965 2789 27999
rect 2789 27965 2823 27999
rect 2823 27965 2832 27999
rect 2780 27956 2832 27965
rect 2964 27956 3016 28008
rect 3792 27999 3844 28008
rect 3792 27965 3801 27999
rect 3801 27965 3835 27999
rect 3835 27965 3844 27999
rect 3792 27956 3844 27965
rect 4896 27999 4948 28008
rect 4896 27965 4905 27999
rect 4905 27965 4939 27999
rect 4939 27965 4948 27999
rect 4896 27956 4948 27965
rect 6184 28135 6236 28144
rect 6184 28101 6193 28135
rect 6193 28101 6227 28135
rect 6227 28101 6236 28135
rect 6184 28092 6236 28101
rect 7104 28169 7113 28203
rect 7113 28169 7147 28203
rect 7147 28169 7156 28203
rect 7104 28160 7156 28169
rect 11060 28160 11112 28212
rect 14832 28203 14884 28212
rect 14832 28169 14841 28203
rect 14841 28169 14875 28203
rect 14875 28169 14884 28203
rect 14832 28160 14884 28169
rect 16764 28160 16816 28212
rect 17776 28160 17828 28212
rect 17960 28160 18012 28212
rect 18236 28160 18288 28212
rect 18512 28160 18564 28212
rect 20536 28160 20588 28212
rect 24676 28160 24728 28212
rect 29000 28160 29052 28212
rect 29920 28160 29972 28212
rect 30288 28203 30340 28212
rect 30288 28169 30297 28203
rect 30297 28169 30331 28203
rect 30331 28169 30340 28203
rect 30288 28160 30340 28169
rect 8300 28092 8352 28144
rect 6460 28024 6512 28076
rect 7196 28024 7248 28076
rect 7564 28067 7616 28076
rect 7564 28033 7573 28067
rect 7573 28033 7607 28067
rect 7607 28033 7616 28067
rect 7564 28024 7616 28033
rect 8208 28024 8260 28076
rect 13452 28024 13504 28076
rect 19432 28092 19484 28144
rect 20076 28092 20128 28144
rect 24400 28092 24452 28144
rect 17500 28024 17552 28076
rect 17776 28024 17828 28076
rect 17960 28024 18012 28076
rect 18052 28024 18104 28076
rect 4252 27888 4304 27940
rect 2780 27820 2832 27872
rect 3240 27820 3292 27872
rect 4528 27820 4580 27872
rect 4804 27820 4856 27872
rect 5428 27888 5480 27940
rect 7104 27956 7156 28008
rect 7288 27999 7340 28008
rect 7288 27965 7297 27999
rect 7297 27965 7331 27999
rect 7331 27965 7340 27999
rect 7288 27956 7340 27965
rect 7840 27999 7892 28008
rect 6460 27888 6512 27940
rect 7840 27965 7849 27999
rect 7849 27965 7883 27999
rect 7883 27965 7892 27999
rect 7840 27956 7892 27965
rect 9036 27956 9088 28008
rect 9404 27999 9456 28008
rect 9404 27965 9413 27999
rect 9413 27965 9447 27999
rect 9447 27965 9456 27999
rect 9404 27956 9456 27965
rect 10232 27956 10284 28008
rect 12348 27956 12400 28008
rect 12624 27956 12676 28008
rect 14096 27999 14148 28008
rect 14096 27965 14105 27999
rect 14105 27965 14139 27999
rect 14139 27965 14148 27999
rect 14096 27956 14148 27965
rect 14280 27999 14332 28008
rect 14280 27965 14289 27999
rect 14289 27965 14323 27999
rect 14323 27965 14332 27999
rect 14280 27956 14332 27965
rect 14648 27999 14700 28008
rect 11152 27888 11204 27940
rect 12808 27888 12860 27940
rect 12992 27931 13044 27940
rect 12992 27897 13001 27931
rect 13001 27897 13035 27931
rect 13035 27897 13044 27931
rect 12992 27888 13044 27897
rect 13912 27888 13964 27940
rect 14188 27888 14240 27940
rect 14648 27965 14657 27999
rect 14657 27965 14691 27999
rect 14691 27965 14700 27999
rect 14648 27956 14700 27965
rect 15292 27956 15344 28008
rect 16304 27956 16356 28008
rect 17132 27956 17184 28008
rect 18144 27956 18196 28008
rect 22928 28024 22980 28076
rect 19616 27999 19668 28008
rect 19616 27965 19625 27999
rect 19625 27965 19659 27999
rect 19659 27965 19668 27999
rect 19616 27956 19668 27965
rect 19800 27999 19852 28008
rect 19800 27965 19809 27999
rect 19809 27965 19843 27999
rect 19843 27965 19852 27999
rect 19800 27956 19852 27965
rect 21180 27999 21232 28008
rect 17960 27888 18012 27940
rect 21180 27965 21189 27999
rect 21189 27965 21223 27999
rect 21223 27965 21232 27999
rect 21180 27956 21232 27965
rect 21272 27956 21324 28008
rect 22008 27999 22060 28008
rect 22008 27965 22017 27999
rect 22017 27965 22051 27999
rect 22051 27965 22060 27999
rect 23848 28024 23900 28076
rect 24860 28067 24912 28076
rect 24860 28033 24869 28067
rect 24869 28033 24903 28067
rect 24903 28033 24912 28067
rect 24860 28024 24912 28033
rect 27528 28067 27580 28076
rect 27528 28033 27537 28067
rect 27537 28033 27571 28067
rect 27571 28033 27580 28067
rect 27528 28024 27580 28033
rect 29092 28024 29144 28076
rect 22008 27956 22060 27965
rect 8208 27820 8260 27872
rect 9496 27820 9548 27872
rect 11796 27820 11848 27872
rect 14740 27820 14792 27872
rect 15936 27820 15988 27872
rect 23664 27888 23716 27940
rect 24492 27956 24544 28008
rect 27620 27956 27672 28008
rect 28632 27956 28684 28008
rect 29552 27999 29604 28008
rect 29552 27965 29561 27999
rect 29561 27965 29595 27999
rect 29595 27965 29604 27999
rect 29552 27956 29604 27965
rect 19248 27820 19300 27872
rect 25688 27820 25740 27872
rect 25780 27820 25832 27872
rect 26424 27820 26476 27872
rect 26608 27820 26660 27872
rect 27620 27820 27672 27872
rect 28264 27820 28316 27872
rect 28816 27820 28868 27872
rect 29920 27999 29972 28008
rect 29920 27965 29929 27999
rect 29929 27965 29963 27999
rect 29963 27965 29972 27999
rect 29920 27956 29972 27965
rect 31116 27999 31168 28008
rect 31116 27965 31125 27999
rect 31125 27965 31159 27999
rect 31159 27965 31168 27999
rect 31116 27956 31168 27965
rect 30012 27888 30064 27940
rect 11253 27718 11305 27770
rect 11317 27718 11369 27770
rect 11381 27718 11433 27770
rect 11445 27718 11497 27770
rect 11509 27718 11561 27770
rect 21557 27718 21609 27770
rect 21621 27718 21673 27770
rect 21685 27718 21737 27770
rect 21749 27718 21801 27770
rect 21813 27718 21865 27770
rect 1492 27616 1544 27668
rect 2688 27616 2740 27668
rect 1584 27591 1636 27600
rect 1584 27557 1593 27591
rect 1593 27557 1627 27591
rect 1627 27557 1636 27591
rect 1584 27548 1636 27557
rect 1952 27548 2004 27600
rect 2780 27548 2832 27600
rect 3608 27548 3660 27600
rect 6000 27548 6052 27600
rect 1400 27412 1452 27464
rect 2044 27480 2096 27532
rect 2228 27480 2280 27532
rect 3332 27523 3384 27532
rect 3332 27489 3341 27523
rect 3341 27489 3375 27523
rect 3375 27489 3384 27523
rect 3332 27480 3384 27489
rect 3516 27523 3568 27532
rect 3516 27489 3525 27523
rect 3525 27489 3559 27523
rect 3559 27489 3568 27523
rect 3516 27480 3568 27489
rect 3884 27523 3936 27532
rect 3884 27489 3893 27523
rect 3893 27489 3927 27523
rect 3927 27489 3936 27523
rect 3884 27480 3936 27489
rect 4896 27480 4948 27532
rect 2504 27412 2556 27464
rect 3240 27412 3292 27464
rect 4160 27412 4212 27464
rect 4344 27412 4396 27464
rect 1676 27344 1728 27396
rect 4712 27344 4764 27396
rect 7104 27616 7156 27668
rect 6644 27548 6696 27600
rect 6276 27412 6328 27464
rect 6460 27412 6512 27464
rect 6920 27480 6972 27532
rect 7748 27548 7800 27600
rect 9680 27616 9732 27668
rect 10968 27548 11020 27600
rect 11244 27548 11296 27600
rect 7564 27455 7616 27464
rect 7564 27421 7573 27455
rect 7573 27421 7607 27455
rect 7607 27421 7616 27455
rect 7564 27412 7616 27421
rect 7196 27344 7248 27396
rect 7840 27523 7892 27532
rect 7840 27489 7849 27523
rect 7849 27489 7883 27523
rect 7883 27489 7892 27523
rect 7840 27480 7892 27489
rect 8392 27480 8444 27532
rect 8576 27480 8628 27532
rect 10232 27480 10284 27532
rect 11980 27480 12032 27532
rect 15016 27616 15068 27668
rect 12992 27480 13044 27532
rect 14096 27480 14148 27532
rect 14648 27480 14700 27532
rect 15660 27523 15712 27532
rect 15660 27489 15669 27523
rect 15669 27489 15703 27523
rect 15703 27489 15712 27523
rect 15660 27480 15712 27489
rect 9496 27344 9548 27396
rect 15936 27455 15988 27464
rect 15936 27421 15945 27455
rect 15945 27421 15979 27455
rect 15979 27421 15988 27455
rect 15936 27412 15988 27421
rect 17684 27548 17736 27600
rect 18604 27591 18656 27600
rect 16856 27523 16908 27532
rect 16856 27489 16865 27523
rect 16865 27489 16899 27523
rect 16899 27489 16908 27523
rect 16856 27480 16908 27489
rect 17132 27523 17184 27532
rect 17132 27489 17141 27523
rect 17141 27489 17175 27523
rect 17175 27489 17184 27523
rect 17132 27480 17184 27489
rect 17316 27480 17368 27532
rect 17776 27480 17828 27532
rect 18052 27523 18104 27532
rect 18052 27489 18061 27523
rect 18061 27489 18095 27523
rect 18095 27489 18104 27523
rect 18052 27480 18104 27489
rect 18604 27557 18613 27591
rect 18613 27557 18647 27591
rect 18647 27557 18656 27591
rect 18604 27548 18656 27557
rect 18788 27616 18840 27668
rect 19524 27616 19576 27668
rect 19616 27616 19668 27668
rect 21180 27659 21232 27668
rect 21180 27625 21189 27659
rect 21189 27625 21223 27659
rect 21223 27625 21232 27659
rect 21180 27616 21232 27625
rect 18972 27548 19024 27600
rect 19156 27548 19208 27600
rect 19064 27523 19116 27532
rect 19064 27489 19073 27523
rect 19073 27489 19107 27523
rect 19107 27489 19116 27523
rect 19064 27480 19116 27489
rect 19248 27523 19300 27532
rect 19248 27489 19257 27523
rect 19257 27489 19291 27523
rect 19291 27489 19300 27523
rect 19248 27480 19300 27489
rect 19984 27548 20036 27600
rect 1308 27276 1360 27328
rect 3792 27276 3844 27328
rect 4528 27276 4580 27328
rect 4896 27276 4948 27328
rect 8760 27276 8812 27328
rect 16212 27344 16264 27396
rect 17684 27412 17736 27464
rect 18144 27455 18196 27464
rect 18144 27421 18153 27455
rect 18153 27421 18187 27455
rect 18187 27421 18196 27455
rect 18144 27412 18196 27421
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 20168 27480 20220 27532
rect 20628 27523 20680 27532
rect 20628 27489 20637 27523
rect 20637 27489 20671 27523
rect 20671 27489 20680 27523
rect 20628 27480 20680 27489
rect 22100 27480 22152 27532
rect 23112 27548 23164 27600
rect 24400 27616 24452 27668
rect 24308 27591 24360 27600
rect 19984 27412 20036 27464
rect 20076 27412 20128 27464
rect 20812 27455 20864 27464
rect 20812 27421 20821 27455
rect 20821 27421 20855 27455
rect 20855 27421 20864 27455
rect 20812 27412 20864 27421
rect 22744 27412 22796 27464
rect 22928 27412 22980 27464
rect 23756 27480 23808 27532
rect 24308 27557 24317 27591
rect 24317 27557 24351 27591
rect 24351 27557 24360 27591
rect 24308 27548 24360 27557
rect 27528 27616 27580 27668
rect 31116 27616 31168 27668
rect 24768 27548 24820 27600
rect 25228 27548 25280 27600
rect 25412 27548 25464 27600
rect 26148 27548 26200 27600
rect 29000 27548 29052 27600
rect 25688 27412 25740 27464
rect 28908 27480 28960 27532
rect 29552 27523 29604 27532
rect 27988 27412 28040 27464
rect 28724 27412 28776 27464
rect 29552 27489 29561 27523
rect 29561 27489 29595 27523
rect 29595 27489 29604 27523
rect 29552 27480 29604 27489
rect 29736 27523 29788 27532
rect 29736 27489 29745 27523
rect 29745 27489 29779 27523
rect 29779 27489 29788 27523
rect 29736 27480 29788 27489
rect 29644 27412 29696 27464
rect 30012 27480 30064 27532
rect 30472 27480 30524 27532
rect 31300 27480 31352 27532
rect 29920 27455 29972 27464
rect 29920 27421 29929 27455
rect 29929 27421 29963 27455
rect 29963 27421 29972 27455
rect 29920 27412 29972 27421
rect 13268 27319 13320 27328
rect 13268 27285 13277 27319
rect 13277 27285 13311 27319
rect 13311 27285 13320 27319
rect 13268 27276 13320 27285
rect 14280 27276 14332 27328
rect 16304 27276 16356 27328
rect 23572 27344 23624 27396
rect 24308 27344 24360 27396
rect 27252 27344 27304 27396
rect 30840 27344 30892 27396
rect 17316 27276 17368 27328
rect 18604 27276 18656 27328
rect 27620 27276 27672 27328
rect 28172 27276 28224 27328
rect 28724 27276 28776 27328
rect 30932 27276 30984 27328
rect 6102 27174 6154 27226
rect 6166 27174 6218 27226
rect 6230 27174 6282 27226
rect 6294 27174 6346 27226
rect 6358 27174 6410 27226
rect 16405 27174 16457 27226
rect 16469 27174 16521 27226
rect 16533 27174 16585 27226
rect 16597 27174 16649 27226
rect 16661 27174 16713 27226
rect 26709 27174 26761 27226
rect 26773 27174 26825 27226
rect 26837 27174 26889 27226
rect 26901 27174 26953 27226
rect 26965 27174 27017 27226
rect 1768 27115 1820 27124
rect 1768 27081 1777 27115
rect 1777 27081 1811 27115
rect 1811 27081 1820 27115
rect 1768 27072 1820 27081
rect 4252 27072 4304 27124
rect 4068 27004 4120 27056
rect 4712 27004 4764 27056
rect 6736 27072 6788 27124
rect 8392 27072 8444 27124
rect 10232 27072 10284 27124
rect 11980 27115 12032 27124
rect 11980 27081 11989 27115
rect 11989 27081 12023 27115
rect 12023 27081 12032 27115
rect 11980 27072 12032 27081
rect 16856 27072 16908 27124
rect 5264 27004 5316 27056
rect 7564 27004 7616 27056
rect 10600 27004 10652 27056
rect 7012 26936 7064 26988
rect 11060 26936 11112 26988
rect 12900 27004 12952 27056
rect 2504 26868 2556 26920
rect 1952 26800 2004 26852
rect 3332 26868 3384 26920
rect 3884 26868 3936 26920
rect 4160 26911 4212 26920
rect 4160 26877 4169 26911
rect 4169 26877 4203 26911
rect 4203 26877 4212 26911
rect 4160 26868 4212 26877
rect 4344 26911 4396 26920
rect 4344 26877 4353 26911
rect 4353 26877 4387 26911
rect 4387 26877 4396 26911
rect 4344 26868 4396 26877
rect 4804 26868 4856 26920
rect 5172 26911 5224 26920
rect 5172 26877 5181 26911
rect 5181 26877 5215 26911
rect 5215 26877 5224 26911
rect 5172 26868 5224 26877
rect 8208 26868 8260 26920
rect 9036 26868 9088 26920
rect 4988 26843 5040 26852
rect 4988 26809 4997 26843
rect 4997 26809 5031 26843
rect 5031 26809 5040 26843
rect 4988 26800 5040 26809
rect 11152 26868 11204 26920
rect 11244 26911 11296 26920
rect 11244 26877 11253 26911
rect 11253 26877 11287 26911
rect 11287 26877 11296 26911
rect 14924 26936 14976 26988
rect 11244 26868 11296 26877
rect 11796 26911 11848 26920
rect 9220 26843 9272 26852
rect 9220 26809 9254 26843
rect 9254 26809 9272 26843
rect 9220 26800 9272 26809
rect 11060 26800 11112 26852
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 11980 26868 12032 26920
rect 11888 26800 11940 26852
rect 12348 26800 12400 26852
rect 13268 26868 13320 26920
rect 13544 26911 13596 26920
rect 13544 26877 13553 26911
rect 13553 26877 13587 26911
rect 13587 26877 13596 26911
rect 13544 26868 13596 26877
rect 13636 26868 13688 26920
rect 14280 26868 14332 26920
rect 16764 26868 16816 26920
rect 14464 26800 14516 26852
rect 14648 26800 14700 26852
rect 15016 26800 15068 26852
rect 2596 26732 2648 26784
rect 2780 26732 2832 26784
rect 3240 26775 3292 26784
rect 3240 26741 3249 26775
rect 3249 26741 3283 26775
rect 3283 26741 3292 26775
rect 3240 26732 3292 26741
rect 3700 26732 3752 26784
rect 4068 26732 4120 26784
rect 16028 26732 16080 26784
rect 16304 26800 16356 26852
rect 16580 26800 16632 26852
rect 17684 26936 17736 26988
rect 18144 26868 18196 26920
rect 19156 27072 19208 27124
rect 19800 27115 19852 27124
rect 19800 27081 19809 27115
rect 19809 27081 19843 27115
rect 19843 27081 19852 27115
rect 19800 27072 19852 27081
rect 20076 27072 20128 27124
rect 19064 27004 19116 27056
rect 20168 27004 20220 27056
rect 20628 27072 20680 27124
rect 21272 27072 21324 27124
rect 23020 27004 23072 27056
rect 23664 27004 23716 27056
rect 24400 27004 24452 27056
rect 24768 27072 24820 27124
rect 25136 27072 25188 27124
rect 27620 27115 27672 27124
rect 27620 27081 27629 27115
rect 27629 27081 27663 27115
rect 27663 27081 27672 27115
rect 27620 27072 27672 27081
rect 28448 27004 28500 27056
rect 20720 26936 20772 26988
rect 22008 26936 22060 26988
rect 22560 26911 22612 26920
rect 18236 26800 18288 26852
rect 17684 26732 17736 26784
rect 17776 26732 17828 26784
rect 18052 26732 18104 26784
rect 18420 26732 18472 26784
rect 18880 26800 18932 26852
rect 19064 26800 19116 26852
rect 19524 26800 19576 26852
rect 20720 26843 20772 26852
rect 20720 26809 20729 26843
rect 20729 26809 20763 26843
rect 20763 26809 20772 26843
rect 20720 26800 20772 26809
rect 20904 26800 20956 26852
rect 21456 26843 21508 26852
rect 21456 26809 21465 26843
rect 21465 26809 21499 26843
rect 21499 26809 21508 26843
rect 21456 26800 21508 26809
rect 22560 26877 22569 26911
rect 22569 26877 22603 26911
rect 22603 26877 22612 26911
rect 22560 26868 22612 26877
rect 22744 26911 22796 26920
rect 22744 26877 22753 26911
rect 22753 26877 22787 26911
rect 22787 26877 22796 26911
rect 22744 26868 22796 26877
rect 23204 26911 23256 26920
rect 23204 26877 23213 26911
rect 23213 26877 23247 26911
rect 23247 26877 23256 26911
rect 23204 26868 23256 26877
rect 25136 26936 25188 26988
rect 25228 26868 25280 26920
rect 26608 26868 26660 26920
rect 26976 26911 27028 26920
rect 26976 26877 26985 26911
rect 26985 26877 27019 26911
rect 27019 26877 27028 26911
rect 26976 26868 27028 26877
rect 27436 26868 27488 26920
rect 29736 26936 29788 26988
rect 31208 26979 31260 26988
rect 31208 26945 31217 26979
rect 31217 26945 31251 26979
rect 31251 26945 31260 26979
rect 31208 26936 31260 26945
rect 29092 26868 29144 26920
rect 30932 26911 30984 26920
rect 30932 26877 30950 26911
rect 30950 26877 30984 26911
rect 30932 26868 30984 26877
rect 23756 26800 23808 26852
rect 25688 26800 25740 26852
rect 27528 26800 27580 26852
rect 31024 26800 31076 26852
rect 21088 26732 21140 26784
rect 24400 26775 24452 26784
rect 24400 26741 24409 26775
rect 24409 26741 24443 26775
rect 24443 26741 24452 26775
rect 24400 26732 24452 26741
rect 24492 26732 24544 26784
rect 26332 26732 26384 26784
rect 27896 26732 27948 26784
rect 28908 26775 28960 26784
rect 28908 26741 28917 26775
rect 28917 26741 28951 26775
rect 28951 26741 28960 26775
rect 28908 26732 28960 26741
rect 30472 26732 30524 26784
rect 11253 26630 11305 26682
rect 11317 26630 11369 26682
rect 11381 26630 11433 26682
rect 11445 26630 11497 26682
rect 11509 26630 11561 26682
rect 21557 26630 21609 26682
rect 21621 26630 21673 26682
rect 21685 26630 21737 26682
rect 21749 26630 21801 26682
rect 21813 26630 21865 26682
rect 2044 26528 2096 26580
rect 3884 26528 3936 26580
rect 5540 26528 5592 26580
rect 6828 26528 6880 26580
rect 7840 26528 7892 26580
rect 8760 26528 8812 26580
rect 15660 26528 15712 26580
rect 17132 26528 17184 26580
rect 17408 26528 17460 26580
rect 17684 26528 17736 26580
rect 20812 26528 20864 26580
rect 22560 26528 22612 26580
rect 28724 26528 28776 26580
rect 1952 26392 2004 26444
rect 4160 26460 4212 26512
rect 4528 26503 4580 26512
rect 4528 26469 4546 26503
rect 4546 26469 4580 26503
rect 4528 26460 4580 26469
rect 7196 26460 7248 26512
rect 2596 26435 2648 26444
rect 2596 26401 2605 26435
rect 2605 26401 2639 26435
rect 2639 26401 2648 26435
rect 2596 26392 2648 26401
rect 5908 26392 5960 26444
rect 6736 26435 6788 26444
rect 6736 26401 6745 26435
rect 6745 26401 6779 26435
rect 6779 26401 6788 26435
rect 6736 26392 6788 26401
rect 6828 26392 6880 26444
rect 7748 26392 7800 26444
rect 8760 26435 8812 26444
rect 8760 26401 8769 26435
rect 8769 26401 8803 26435
rect 8803 26401 8812 26435
rect 8760 26392 8812 26401
rect 9496 26392 9548 26444
rect 11152 26392 11204 26444
rect 11520 26435 11572 26444
rect 11520 26401 11529 26435
rect 11529 26401 11563 26435
rect 11563 26401 11572 26435
rect 11520 26392 11572 26401
rect 11796 26460 11848 26512
rect 11888 26435 11940 26444
rect 11888 26401 11897 26435
rect 11897 26401 11931 26435
rect 11931 26401 11940 26435
rect 11888 26392 11940 26401
rect 11980 26392 12032 26444
rect 12532 26460 12584 26512
rect 16212 26460 16264 26512
rect 16580 26460 16632 26512
rect 12716 26435 12768 26444
rect 12716 26401 12725 26435
rect 12725 26401 12759 26435
rect 12759 26401 12768 26435
rect 12716 26392 12768 26401
rect 12900 26392 12952 26444
rect 13544 26435 13596 26444
rect 13544 26401 13553 26435
rect 13553 26401 13587 26435
rect 13587 26401 13596 26435
rect 13544 26392 13596 26401
rect 13636 26392 13688 26444
rect 15568 26392 15620 26444
rect 15844 26435 15896 26444
rect 15844 26401 15853 26435
rect 15853 26401 15887 26435
rect 15887 26401 15896 26435
rect 15844 26392 15896 26401
rect 16856 26392 16908 26444
rect 3240 26324 3292 26376
rect 4804 26367 4856 26376
rect 4804 26333 4813 26367
rect 4813 26333 4847 26367
rect 4847 26333 4856 26367
rect 4804 26324 4856 26333
rect 8208 26324 8260 26376
rect 10600 26324 10652 26376
rect 12348 26324 12400 26376
rect 2504 26256 2556 26308
rect 8300 26256 8352 26308
rect 1860 26188 1912 26240
rect 2320 26188 2372 26240
rect 5908 26188 5960 26240
rect 6460 26188 6512 26240
rect 7012 26188 7064 26240
rect 9312 26231 9364 26240
rect 9312 26197 9321 26231
rect 9321 26197 9355 26231
rect 9355 26197 9364 26231
rect 9312 26188 9364 26197
rect 11520 26188 11572 26240
rect 12072 26188 12124 26240
rect 12440 26256 12492 26308
rect 12532 26256 12584 26308
rect 13268 26324 13320 26376
rect 14464 26324 14516 26376
rect 16304 26324 16356 26376
rect 16948 26367 17000 26376
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 16948 26324 17000 26333
rect 17132 26435 17184 26444
rect 17132 26401 17141 26435
rect 17141 26401 17175 26435
rect 17175 26401 17184 26435
rect 17132 26392 17184 26401
rect 17868 26435 17920 26444
rect 17868 26401 17877 26435
rect 17877 26401 17911 26435
rect 17911 26401 17920 26435
rect 17868 26392 17920 26401
rect 17960 26392 18012 26444
rect 20720 26460 20772 26512
rect 22652 26460 22704 26512
rect 19708 26392 19760 26444
rect 20444 26435 20496 26444
rect 20444 26401 20453 26435
rect 20453 26401 20487 26435
rect 20487 26401 20496 26435
rect 20444 26392 20496 26401
rect 20536 26435 20588 26444
rect 20536 26401 20545 26435
rect 20545 26401 20579 26435
rect 20579 26401 20588 26435
rect 20536 26392 20588 26401
rect 13084 26256 13136 26308
rect 18420 26324 18472 26376
rect 19984 26324 20036 26376
rect 20168 26324 20220 26376
rect 13820 26188 13872 26240
rect 15384 26188 15436 26240
rect 16212 26188 16264 26240
rect 16304 26188 16356 26240
rect 19340 26256 19392 26308
rect 20720 26256 20772 26308
rect 22284 26392 22336 26444
rect 23204 26460 23256 26512
rect 22008 26256 22060 26308
rect 23112 26392 23164 26444
rect 20812 26188 20864 26240
rect 20996 26231 21048 26240
rect 20996 26197 21005 26231
rect 21005 26197 21039 26231
rect 21039 26197 21048 26231
rect 20996 26188 21048 26197
rect 21088 26188 21140 26240
rect 23204 26324 23256 26376
rect 22652 26256 22704 26308
rect 24032 26460 24084 26512
rect 24400 26460 24452 26512
rect 23572 26435 23624 26444
rect 23572 26401 23581 26435
rect 23581 26401 23615 26435
rect 23615 26401 23624 26435
rect 23572 26392 23624 26401
rect 23848 26392 23900 26444
rect 24676 26392 24728 26444
rect 26240 26460 26292 26512
rect 25136 26392 25188 26444
rect 26148 26392 26200 26444
rect 27712 26435 27764 26444
rect 27712 26401 27721 26435
rect 27721 26401 27755 26435
rect 27755 26401 27764 26435
rect 27712 26392 27764 26401
rect 27896 26435 27948 26444
rect 27896 26401 27905 26435
rect 27905 26401 27939 26435
rect 27939 26401 27948 26435
rect 27896 26392 27948 26401
rect 28908 26392 28960 26444
rect 29276 26392 29328 26444
rect 29552 26392 29604 26444
rect 24032 26324 24084 26376
rect 24952 26324 25004 26376
rect 24308 26256 24360 26308
rect 24584 26299 24636 26308
rect 24584 26265 24593 26299
rect 24593 26265 24627 26299
rect 24627 26265 24636 26299
rect 24584 26256 24636 26265
rect 23020 26188 23072 26240
rect 27252 26324 27304 26376
rect 27528 26324 27580 26376
rect 28080 26367 28132 26376
rect 28080 26333 28089 26367
rect 28089 26333 28123 26367
rect 28123 26333 28132 26367
rect 28080 26324 28132 26333
rect 27160 26256 27212 26308
rect 30012 26435 30064 26444
rect 30012 26401 30021 26435
rect 30021 26401 30055 26435
rect 30055 26401 30064 26435
rect 30012 26392 30064 26401
rect 30564 26392 30616 26444
rect 31024 26392 31076 26444
rect 25872 26231 25924 26240
rect 25872 26197 25881 26231
rect 25881 26197 25915 26231
rect 25915 26197 25924 26231
rect 25872 26188 25924 26197
rect 26516 26188 26568 26240
rect 29552 26256 29604 26308
rect 30472 26324 30524 26376
rect 30656 26324 30708 26376
rect 29920 26256 29972 26308
rect 31024 26256 31076 26308
rect 6102 26086 6154 26138
rect 6166 26086 6218 26138
rect 6230 26086 6282 26138
rect 6294 26086 6346 26138
rect 6358 26086 6410 26138
rect 16405 26086 16457 26138
rect 16469 26086 16521 26138
rect 16533 26086 16585 26138
rect 16597 26086 16649 26138
rect 16661 26086 16713 26138
rect 26709 26086 26761 26138
rect 26773 26086 26825 26138
rect 26837 26086 26889 26138
rect 26901 26086 26953 26138
rect 26965 26086 27017 26138
rect 1400 26027 1452 26036
rect 1400 25993 1409 26027
rect 1409 25993 1443 26027
rect 1443 25993 1452 26027
rect 1400 25984 1452 25993
rect 5172 26027 5224 26036
rect 5172 25993 5181 26027
rect 5181 25993 5215 26027
rect 5215 25993 5224 26027
rect 5172 25984 5224 25993
rect 6828 26027 6880 26036
rect 6828 25993 6837 26027
rect 6837 25993 6871 26027
rect 6871 25993 6880 26027
rect 6828 25984 6880 25993
rect 8208 26027 8260 26036
rect 8208 25993 8217 26027
rect 8217 25993 8251 26027
rect 8251 25993 8260 26027
rect 8208 25984 8260 25993
rect 12808 25984 12860 26036
rect 13084 25984 13136 26036
rect 14280 25984 14332 26036
rect 14372 25984 14424 26036
rect 16120 26027 16172 26036
rect 16120 25993 16129 26027
rect 16129 25993 16163 26027
rect 16163 25993 16172 26027
rect 16120 25984 16172 25993
rect 16948 25984 17000 26036
rect 19708 26027 19760 26036
rect 19708 25993 19717 26027
rect 19717 25993 19751 26027
rect 19751 25993 19760 26027
rect 19708 25984 19760 25993
rect 21456 25984 21508 26036
rect 22560 25984 22612 26036
rect 22744 25984 22796 26036
rect 10876 25916 10928 25968
rect 11980 25916 12032 25968
rect 14924 25916 14976 25968
rect 15476 25916 15528 25968
rect 18052 25916 18104 25968
rect 6644 25848 6696 25900
rect 7748 25848 7800 25900
rect 9036 25891 9088 25900
rect 9036 25857 9045 25891
rect 9045 25857 9079 25891
rect 9079 25857 9088 25891
rect 9036 25848 9088 25857
rect 18512 25916 18564 25968
rect 22100 25916 22152 25968
rect 26424 25916 26476 25968
rect 26700 25916 26752 25968
rect 2504 25823 2556 25832
rect 2504 25789 2522 25823
rect 2522 25789 2556 25823
rect 2504 25780 2556 25789
rect 2780 25823 2832 25832
rect 2780 25789 2789 25823
rect 2789 25789 2823 25823
rect 2823 25789 2832 25823
rect 2780 25780 2832 25789
rect 4804 25780 4856 25832
rect 7012 25823 7064 25832
rect 7012 25789 7021 25823
rect 7021 25789 7055 25823
rect 7055 25789 7064 25823
rect 7012 25780 7064 25789
rect 7196 25823 7248 25832
rect 7196 25789 7205 25823
rect 7205 25789 7239 25823
rect 7239 25789 7248 25823
rect 7196 25780 7248 25789
rect 8024 25823 8076 25832
rect 8024 25789 8033 25823
rect 8033 25789 8067 25823
rect 8067 25789 8076 25823
rect 8024 25780 8076 25789
rect 9312 25823 9364 25832
rect 9312 25789 9346 25823
rect 9346 25789 9364 25823
rect 9312 25780 9364 25789
rect 12440 25780 12492 25832
rect 12992 25823 13044 25832
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 13544 25780 13596 25832
rect 4068 25755 4120 25764
rect 4068 25721 4102 25755
rect 4102 25721 4120 25755
rect 4068 25712 4120 25721
rect 6920 25712 6972 25764
rect 7288 25712 7340 25764
rect 7748 25712 7800 25764
rect 14648 25823 14700 25832
rect 14648 25789 14657 25823
rect 14657 25789 14691 25823
rect 14691 25789 14700 25823
rect 14648 25780 14700 25789
rect 18144 25780 18196 25832
rect 18420 25823 18472 25832
rect 18420 25789 18429 25823
rect 18429 25789 18463 25823
rect 18463 25789 18472 25823
rect 18420 25780 18472 25789
rect 18604 25823 18656 25832
rect 18604 25789 18613 25823
rect 18613 25789 18647 25823
rect 18647 25789 18656 25823
rect 18604 25780 18656 25789
rect 22192 25848 22244 25900
rect 22744 25848 22796 25900
rect 25688 25848 25740 25900
rect 26516 25848 26568 25900
rect 27528 25984 27580 26036
rect 27712 26027 27764 26036
rect 27712 25993 27721 26027
rect 27721 25993 27755 26027
rect 27755 25993 27764 26027
rect 27712 25984 27764 25993
rect 20260 25780 20312 25832
rect 22284 25780 22336 25832
rect 23296 25780 23348 25832
rect 15016 25755 15068 25764
rect 15016 25721 15025 25755
rect 15025 25721 15059 25755
rect 15059 25721 15068 25755
rect 15016 25712 15068 25721
rect 5540 25644 5592 25696
rect 6828 25644 6880 25696
rect 8208 25644 8260 25696
rect 8484 25644 8536 25696
rect 10416 25687 10468 25696
rect 10416 25653 10425 25687
rect 10425 25653 10459 25687
rect 10459 25653 10468 25687
rect 10416 25644 10468 25653
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 13268 25644 13320 25696
rect 14464 25644 14516 25696
rect 15384 25644 15436 25696
rect 18880 25712 18932 25764
rect 20076 25712 20128 25764
rect 21916 25712 21968 25764
rect 24676 25823 24728 25832
rect 24676 25789 24685 25823
rect 24685 25789 24719 25823
rect 24719 25789 24728 25823
rect 24676 25780 24728 25789
rect 25044 25780 25096 25832
rect 25872 25780 25924 25832
rect 26056 25780 26108 25832
rect 27344 25916 27396 25968
rect 27436 25916 27488 25968
rect 27252 25848 27304 25900
rect 28816 25848 28868 25900
rect 28264 25823 28316 25832
rect 24768 25712 24820 25764
rect 26516 25712 26568 25764
rect 28264 25789 28273 25823
rect 28273 25789 28307 25823
rect 28307 25789 28316 25823
rect 28264 25780 28316 25789
rect 31024 25823 31076 25832
rect 31024 25789 31042 25823
rect 31042 25789 31076 25823
rect 31024 25780 31076 25789
rect 31208 25780 31260 25832
rect 20168 25644 20220 25696
rect 20536 25644 20588 25696
rect 22008 25644 22060 25696
rect 24032 25644 24084 25696
rect 24584 25644 24636 25696
rect 25964 25687 26016 25696
rect 25964 25653 25973 25687
rect 25973 25653 26007 25687
rect 26007 25653 26016 25687
rect 25964 25644 26016 25653
rect 26424 25687 26476 25696
rect 26424 25653 26433 25687
rect 26433 25653 26467 25687
rect 26467 25653 26476 25687
rect 26424 25644 26476 25653
rect 29460 25644 29512 25696
rect 30012 25644 30064 25696
rect 11253 25542 11305 25594
rect 11317 25542 11369 25594
rect 11381 25542 11433 25594
rect 11445 25542 11497 25594
rect 11509 25542 11561 25594
rect 21557 25542 21609 25594
rect 21621 25542 21673 25594
rect 21685 25542 21737 25594
rect 21749 25542 21801 25594
rect 21813 25542 21865 25594
rect 3424 25440 3476 25492
rect 4068 25440 4120 25492
rect 5080 25440 5132 25492
rect 5908 25440 5960 25492
rect 6552 25440 6604 25492
rect 13636 25440 13688 25492
rect 15660 25440 15712 25492
rect 17132 25440 17184 25492
rect 3332 25372 3384 25424
rect 5724 25372 5776 25424
rect 8484 25372 8536 25424
rect 9496 25415 9548 25424
rect 9496 25381 9505 25415
rect 9505 25381 9539 25415
rect 9539 25381 9548 25415
rect 9496 25372 9548 25381
rect 9680 25415 9732 25424
rect 9680 25381 9689 25415
rect 9689 25381 9723 25415
rect 9723 25381 9732 25415
rect 9680 25372 9732 25381
rect 10416 25372 10468 25424
rect 10600 25372 10652 25424
rect 12900 25372 12952 25424
rect 13176 25415 13228 25424
rect 13176 25381 13185 25415
rect 13185 25381 13219 25415
rect 13219 25381 13228 25415
rect 13176 25372 13228 25381
rect 17776 25415 17828 25424
rect 2872 25304 2924 25356
rect 6828 25347 6880 25356
rect 6828 25313 6837 25347
rect 6837 25313 6871 25347
rect 6871 25313 6880 25347
rect 6828 25304 6880 25313
rect 7840 25304 7892 25356
rect 8300 25347 8352 25356
rect 8300 25313 8309 25347
rect 8309 25313 8343 25347
rect 8343 25313 8352 25347
rect 8300 25304 8352 25313
rect 9588 25304 9640 25356
rect 11060 25304 11112 25356
rect 11980 25304 12032 25356
rect 13452 25304 13504 25356
rect 13636 25304 13688 25356
rect 14188 25347 14240 25356
rect 1952 25168 2004 25220
rect 9036 25236 9088 25288
rect 12072 25279 12124 25288
rect 12072 25245 12081 25279
rect 12081 25245 12115 25279
rect 12115 25245 12124 25279
rect 12072 25236 12124 25245
rect 13912 25236 13964 25288
rect 3700 25168 3752 25220
rect 9772 25168 9824 25220
rect 1492 25100 1544 25152
rect 3424 25100 3476 25152
rect 4344 25100 4396 25152
rect 5264 25100 5316 25152
rect 7748 25100 7800 25152
rect 12716 25100 12768 25152
rect 14188 25313 14197 25347
rect 14197 25313 14231 25347
rect 14231 25313 14240 25347
rect 14188 25304 14240 25313
rect 14372 25347 14424 25356
rect 14372 25313 14381 25347
rect 14381 25313 14415 25347
rect 14415 25313 14424 25347
rect 14372 25304 14424 25313
rect 17776 25381 17810 25415
rect 17810 25381 17828 25415
rect 17776 25372 17828 25381
rect 18144 25440 18196 25492
rect 21272 25440 21324 25492
rect 24492 25483 24544 25492
rect 20720 25372 20772 25424
rect 15384 25347 15436 25356
rect 14096 25236 14148 25288
rect 14464 25236 14516 25288
rect 15384 25313 15393 25347
rect 15393 25313 15427 25347
rect 15427 25313 15436 25347
rect 15384 25304 15436 25313
rect 14648 25236 14700 25288
rect 15568 25236 15620 25288
rect 14188 25168 14240 25220
rect 15936 25304 15988 25356
rect 16764 25304 16816 25356
rect 18788 25304 18840 25356
rect 20996 25304 21048 25356
rect 15936 25211 15988 25220
rect 15936 25177 15945 25211
rect 15945 25177 15979 25211
rect 15979 25177 15988 25211
rect 15936 25168 15988 25177
rect 18604 25168 18656 25220
rect 20904 25236 20956 25288
rect 22284 25304 22336 25356
rect 24124 25372 24176 25424
rect 24492 25449 24501 25483
rect 24501 25449 24535 25483
rect 24535 25449 24544 25483
rect 24492 25440 24544 25449
rect 25964 25440 26016 25492
rect 24400 25304 24452 25356
rect 24768 25372 24820 25424
rect 24952 25347 25004 25356
rect 24952 25313 24961 25347
rect 24961 25313 24995 25347
rect 24995 25313 25004 25347
rect 24952 25304 25004 25313
rect 25044 25304 25096 25356
rect 25320 25304 25372 25356
rect 25412 25304 25464 25356
rect 25872 25236 25924 25288
rect 22100 25168 22152 25220
rect 16764 25100 16816 25152
rect 16948 25100 17000 25152
rect 25964 25168 26016 25220
rect 26148 25304 26200 25356
rect 27252 25347 27304 25356
rect 27252 25313 27261 25347
rect 27261 25313 27295 25347
rect 27295 25313 27304 25347
rect 27252 25304 27304 25313
rect 28816 25304 28868 25356
rect 29276 25347 29328 25356
rect 29276 25313 29285 25347
rect 29285 25313 29319 25347
rect 29319 25313 29328 25347
rect 29276 25304 29328 25313
rect 29460 25347 29512 25356
rect 29460 25313 29469 25347
rect 29469 25313 29503 25347
rect 29503 25313 29512 25347
rect 29460 25304 29512 25313
rect 29552 25347 29604 25356
rect 29552 25313 29561 25347
rect 29561 25313 29595 25347
rect 29595 25313 29604 25347
rect 29552 25304 29604 25313
rect 29736 25304 29788 25356
rect 30472 25347 30524 25356
rect 30472 25313 30481 25347
rect 30481 25313 30515 25347
rect 30515 25313 30524 25347
rect 30472 25304 30524 25313
rect 31300 25304 31352 25356
rect 27988 25279 28040 25288
rect 27988 25245 27997 25279
rect 27997 25245 28031 25279
rect 28031 25245 28040 25279
rect 27988 25236 28040 25245
rect 28540 25236 28592 25288
rect 25228 25143 25280 25152
rect 25228 25109 25237 25143
rect 25237 25109 25271 25143
rect 25271 25109 25280 25143
rect 25228 25100 25280 25109
rect 25412 25100 25464 25152
rect 26700 25168 26752 25220
rect 27436 25100 27488 25152
rect 27620 25100 27672 25152
rect 30380 25100 30432 25152
rect 6102 24998 6154 25050
rect 6166 24998 6218 25050
rect 6230 24998 6282 25050
rect 6294 24998 6346 25050
rect 6358 24998 6410 25050
rect 16405 24998 16457 25050
rect 16469 24998 16521 25050
rect 16533 24998 16585 25050
rect 16597 24998 16649 25050
rect 16661 24998 16713 25050
rect 26709 24998 26761 25050
rect 26773 24998 26825 25050
rect 26837 24998 26889 25050
rect 26901 24998 26953 25050
rect 26965 24998 27017 25050
rect 5356 24896 5408 24948
rect 4344 24828 4396 24880
rect 2780 24803 2832 24812
rect 2780 24769 2789 24803
rect 2789 24769 2823 24803
rect 2823 24769 2832 24803
rect 2780 24760 2832 24769
rect 1952 24692 2004 24744
rect 4804 24760 4856 24812
rect 1860 24624 1912 24676
rect 2136 24624 2188 24676
rect 2504 24667 2556 24676
rect 2504 24633 2522 24667
rect 2522 24633 2556 24667
rect 2504 24624 2556 24633
rect 3700 24624 3752 24676
rect 4160 24735 4212 24744
rect 4160 24701 4169 24735
rect 4169 24701 4203 24735
rect 4203 24701 4212 24735
rect 4160 24692 4212 24701
rect 10416 24896 10468 24948
rect 11336 24896 11388 24948
rect 13912 24896 13964 24948
rect 15200 24896 15252 24948
rect 16212 24896 16264 24948
rect 22284 24896 22336 24948
rect 22468 24896 22520 24948
rect 23296 24896 23348 24948
rect 23572 24896 23624 24948
rect 24400 24939 24452 24948
rect 24400 24905 24409 24939
rect 24409 24905 24443 24939
rect 24443 24905 24452 24939
rect 24400 24896 24452 24905
rect 24492 24896 24544 24948
rect 10324 24828 10376 24880
rect 10784 24828 10836 24880
rect 14096 24828 14148 24880
rect 6552 24760 6604 24812
rect 7472 24760 7524 24812
rect 9588 24760 9640 24812
rect 10600 24760 10652 24812
rect 8024 24692 8076 24744
rect 8760 24692 8812 24744
rect 9496 24692 9548 24744
rect 9956 24692 10008 24744
rect 10232 24692 10284 24744
rect 10968 24735 11020 24744
rect 2044 24556 2096 24608
rect 2412 24556 2464 24608
rect 2780 24556 2832 24608
rect 3516 24556 3568 24608
rect 5080 24624 5132 24676
rect 10968 24701 10977 24735
rect 10977 24701 11011 24735
rect 11011 24701 11020 24735
rect 10968 24692 11020 24701
rect 11152 24735 11204 24744
rect 11152 24701 11161 24735
rect 11161 24701 11195 24735
rect 11195 24701 11204 24735
rect 11152 24692 11204 24701
rect 11336 24735 11388 24744
rect 11336 24701 11345 24735
rect 11345 24701 11379 24735
rect 11379 24701 11388 24735
rect 12348 24735 12400 24744
rect 11336 24692 11388 24701
rect 12348 24701 12357 24735
rect 12357 24701 12391 24735
rect 12391 24701 12400 24735
rect 12348 24692 12400 24701
rect 12532 24735 12584 24744
rect 12532 24701 12541 24735
rect 12541 24701 12575 24735
rect 12575 24701 12584 24735
rect 12532 24692 12584 24701
rect 12072 24624 12124 24676
rect 4528 24599 4580 24608
rect 4528 24565 4537 24599
rect 4537 24565 4571 24599
rect 4571 24565 4580 24599
rect 4528 24556 4580 24565
rect 6368 24599 6420 24608
rect 6368 24565 6377 24599
rect 6377 24565 6411 24599
rect 6411 24565 6420 24599
rect 6368 24556 6420 24565
rect 9036 24599 9088 24608
rect 9036 24565 9045 24599
rect 9045 24565 9079 24599
rect 9079 24565 9088 24599
rect 9036 24556 9088 24565
rect 10784 24556 10836 24608
rect 11704 24556 11756 24608
rect 11796 24556 11848 24608
rect 18328 24760 18380 24812
rect 20904 24828 20956 24880
rect 23204 24871 23256 24880
rect 23204 24837 23213 24871
rect 23213 24837 23247 24871
rect 23247 24837 23256 24871
rect 23204 24828 23256 24837
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 20444 24760 20496 24812
rect 22744 24760 22796 24812
rect 25136 24803 25188 24812
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25136 24760 25188 24769
rect 12808 24692 12860 24744
rect 13452 24692 13504 24744
rect 13544 24692 13596 24744
rect 14740 24692 14792 24744
rect 17684 24692 17736 24744
rect 18696 24735 18748 24744
rect 18696 24701 18705 24735
rect 18705 24701 18739 24735
rect 18739 24701 18748 24735
rect 18696 24692 18748 24701
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 14464 24624 14516 24676
rect 15108 24624 15160 24676
rect 17040 24667 17092 24676
rect 17040 24633 17049 24667
rect 17049 24633 17083 24667
rect 17083 24633 17092 24667
rect 17040 24624 17092 24633
rect 19616 24735 19668 24744
rect 19616 24701 19625 24735
rect 19625 24701 19659 24735
rect 19659 24701 19668 24735
rect 19616 24692 19668 24701
rect 19800 24692 19852 24744
rect 20812 24692 20864 24744
rect 21088 24624 21140 24676
rect 12992 24556 13044 24608
rect 15568 24556 15620 24608
rect 21364 24624 21416 24676
rect 23112 24692 23164 24744
rect 24584 24735 24636 24744
rect 24584 24701 24593 24735
rect 24593 24701 24627 24735
rect 24627 24701 24636 24735
rect 24584 24692 24636 24701
rect 21916 24556 21968 24608
rect 24124 24624 24176 24676
rect 24952 24624 25004 24676
rect 26608 24896 26660 24948
rect 26424 24828 26476 24880
rect 27528 24760 27580 24812
rect 26424 24735 26476 24744
rect 26424 24701 26433 24735
rect 26433 24701 26467 24735
rect 26467 24701 26476 24735
rect 26424 24692 26476 24701
rect 26608 24735 26660 24744
rect 26608 24701 26617 24735
rect 26617 24701 26651 24735
rect 26651 24701 26660 24735
rect 26608 24692 26660 24701
rect 27068 24692 27120 24744
rect 27620 24735 27672 24744
rect 27620 24701 27629 24735
rect 27629 24701 27663 24735
rect 27663 24701 27672 24735
rect 27620 24692 27672 24701
rect 27804 24735 27856 24744
rect 27804 24701 27813 24735
rect 27813 24701 27847 24735
rect 27847 24701 27856 24735
rect 27804 24692 27856 24701
rect 26240 24624 26292 24676
rect 22468 24556 22520 24608
rect 23388 24556 23440 24608
rect 27160 24624 27212 24676
rect 27344 24624 27396 24676
rect 28080 24760 28132 24812
rect 31208 24760 31260 24812
rect 29000 24735 29052 24744
rect 29000 24701 29009 24735
rect 29009 24701 29043 24735
rect 29043 24701 29052 24735
rect 29000 24692 29052 24701
rect 30380 24692 30432 24744
rect 26700 24556 26752 24608
rect 29000 24556 29052 24608
rect 29736 24556 29788 24608
rect 11253 24454 11305 24506
rect 11317 24454 11369 24506
rect 11381 24454 11433 24506
rect 11445 24454 11497 24506
rect 11509 24454 11561 24506
rect 21557 24454 21609 24506
rect 21621 24454 21673 24506
rect 21685 24454 21737 24506
rect 21749 24454 21801 24506
rect 21813 24454 21865 24506
rect 1952 24352 2004 24404
rect 2044 24352 2096 24404
rect 2504 24352 2556 24404
rect 5080 24395 5132 24404
rect 5080 24361 5089 24395
rect 5089 24361 5123 24395
rect 5123 24361 5132 24395
rect 5080 24352 5132 24361
rect 7932 24352 7984 24404
rect 2044 24259 2096 24268
rect 2044 24225 2053 24259
rect 2053 24225 2087 24259
rect 2087 24225 2096 24259
rect 2044 24216 2096 24225
rect 2136 24191 2188 24200
rect 2136 24157 2145 24191
rect 2145 24157 2179 24191
rect 2179 24157 2188 24191
rect 2136 24148 2188 24157
rect 4160 24284 4212 24336
rect 4804 24284 4856 24336
rect 8116 24352 8168 24404
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 2044 24080 2096 24132
rect 4252 24080 4304 24132
rect 5448 24259 5500 24268
rect 5448 24225 5457 24259
rect 5457 24225 5491 24259
rect 5491 24225 5500 24259
rect 5632 24259 5684 24268
rect 5448 24216 5500 24225
rect 5632 24225 5641 24259
rect 5641 24225 5675 24259
rect 5675 24225 5684 24259
rect 5632 24216 5684 24225
rect 6000 24216 6052 24268
rect 7840 24216 7892 24268
rect 6552 24148 6604 24200
rect 8576 24148 8628 24200
rect 5816 24080 5868 24132
rect 6368 24080 6420 24132
rect 7012 24012 7064 24064
rect 9496 24284 9548 24336
rect 9588 24216 9640 24268
rect 9956 24259 10008 24268
rect 9956 24225 9965 24259
rect 9965 24225 9999 24259
rect 9999 24225 10008 24259
rect 9956 24216 10008 24225
rect 11152 24352 11204 24404
rect 15292 24352 15344 24404
rect 16028 24395 16080 24404
rect 16028 24361 16037 24395
rect 16037 24361 16071 24395
rect 16071 24361 16080 24395
rect 16028 24352 16080 24361
rect 18788 24352 18840 24404
rect 19340 24352 19392 24404
rect 19524 24352 19576 24404
rect 10968 24284 11020 24336
rect 12532 24284 12584 24336
rect 12716 24284 12768 24336
rect 13268 24284 13320 24336
rect 15108 24284 15160 24336
rect 10784 24216 10836 24268
rect 11060 24216 11112 24268
rect 11520 24259 11572 24268
rect 11520 24225 11529 24259
rect 11529 24225 11563 24259
rect 11563 24225 11572 24259
rect 11520 24216 11572 24225
rect 12992 24259 13044 24268
rect 12992 24225 13001 24259
rect 13001 24225 13035 24259
rect 13035 24225 13044 24259
rect 12992 24216 13044 24225
rect 13176 24259 13228 24268
rect 13176 24225 13185 24259
rect 13185 24225 13219 24259
rect 13219 24225 13228 24259
rect 13176 24216 13228 24225
rect 13820 24216 13872 24268
rect 14188 24216 14240 24268
rect 16948 24216 17000 24268
rect 17408 24216 17460 24268
rect 18144 24259 18196 24268
rect 18144 24225 18153 24259
rect 18153 24225 18187 24259
rect 18187 24225 18196 24259
rect 18144 24216 18196 24225
rect 18236 24259 18288 24268
rect 18236 24225 18245 24259
rect 18245 24225 18279 24259
rect 18279 24225 18288 24259
rect 18236 24216 18288 24225
rect 18604 24216 18656 24268
rect 19432 24259 19484 24268
rect 19432 24225 19441 24259
rect 19441 24225 19475 24259
rect 19475 24225 19484 24259
rect 19432 24216 19484 24225
rect 14648 24191 14700 24200
rect 11612 24080 11664 24132
rect 9220 24012 9272 24064
rect 9956 24055 10008 24064
rect 9956 24021 9965 24055
rect 9965 24021 9999 24055
rect 9999 24021 10008 24055
rect 9956 24012 10008 24021
rect 10600 24012 10652 24064
rect 11060 24012 11112 24064
rect 14648 24157 14657 24191
rect 14657 24157 14691 24191
rect 14691 24157 14700 24191
rect 14648 24148 14700 24157
rect 16212 24148 16264 24200
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 19156 24148 19208 24200
rect 18788 24080 18840 24132
rect 16304 24012 16356 24064
rect 19892 24216 19944 24268
rect 20812 24284 20864 24336
rect 21364 24352 21416 24404
rect 23848 24352 23900 24404
rect 24124 24352 24176 24404
rect 20628 24216 20680 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21088 24259 21140 24268
rect 21088 24225 21097 24259
rect 21097 24225 21131 24259
rect 21131 24225 21140 24259
rect 21088 24216 21140 24225
rect 19616 24148 19668 24200
rect 19984 24148 20036 24200
rect 22284 24080 22336 24132
rect 21548 24012 21600 24064
rect 23388 24284 23440 24336
rect 22560 24259 22612 24268
rect 22560 24225 22569 24259
rect 22569 24225 22603 24259
rect 22603 24225 22612 24259
rect 22560 24216 22612 24225
rect 23204 24216 23256 24268
rect 23020 24148 23072 24200
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 22744 24012 22796 24064
rect 24308 24284 24360 24336
rect 25688 24284 25740 24336
rect 24860 24259 24912 24268
rect 24860 24225 24869 24259
rect 24869 24225 24903 24259
rect 24903 24225 24912 24259
rect 24860 24216 24912 24225
rect 25320 24216 25372 24268
rect 25964 24216 26016 24268
rect 26424 24352 26476 24404
rect 27068 24352 27120 24404
rect 27804 24352 27856 24404
rect 28816 24395 28868 24404
rect 28816 24361 28825 24395
rect 28825 24361 28859 24395
rect 28859 24361 28868 24395
rect 28816 24352 28868 24361
rect 29828 24352 29880 24404
rect 30564 24395 30616 24404
rect 30564 24361 30573 24395
rect 30573 24361 30607 24395
rect 30607 24361 30616 24395
rect 30564 24352 30616 24361
rect 30840 24352 30892 24404
rect 26332 24284 26384 24336
rect 27160 24327 27212 24336
rect 27160 24293 27169 24327
rect 27169 24293 27203 24327
rect 27203 24293 27212 24327
rect 27160 24284 27212 24293
rect 30288 24284 30340 24336
rect 31300 24284 31352 24336
rect 26700 24216 26752 24268
rect 28816 24216 28868 24268
rect 29460 24216 29512 24268
rect 31116 24259 31168 24268
rect 31116 24225 31125 24259
rect 31125 24225 31159 24259
rect 31159 24225 31168 24259
rect 31116 24216 31168 24225
rect 24216 24148 24268 24200
rect 24768 24148 24820 24200
rect 25136 24148 25188 24200
rect 25412 24148 25464 24200
rect 31024 24080 31076 24132
rect 23204 24012 23256 24064
rect 24584 24012 24636 24064
rect 24952 24012 25004 24064
rect 26332 24055 26384 24064
rect 26332 24021 26341 24055
rect 26341 24021 26375 24055
rect 26375 24021 26384 24055
rect 26332 24012 26384 24021
rect 6102 23910 6154 23962
rect 6166 23910 6218 23962
rect 6230 23910 6282 23962
rect 6294 23910 6346 23962
rect 6358 23910 6410 23962
rect 16405 23910 16457 23962
rect 16469 23910 16521 23962
rect 16533 23910 16585 23962
rect 16597 23910 16649 23962
rect 16661 23910 16713 23962
rect 26709 23910 26761 23962
rect 26773 23910 26825 23962
rect 26837 23910 26889 23962
rect 26901 23910 26953 23962
rect 26965 23910 27017 23962
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 1584 23468 1636 23520
rect 3516 23808 3568 23860
rect 3148 23740 3200 23792
rect 5540 23808 5592 23860
rect 7840 23808 7892 23860
rect 6736 23740 6788 23792
rect 6000 23672 6052 23724
rect 4528 23604 4580 23656
rect 5172 23647 5224 23656
rect 5172 23613 5181 23647
rect 5181 23613 5215 23647
rect 5215 23613 5224 23647
rect 5172 23604 5224 23613
rect 5908 23604 5960 23656
rect 5540 23536 5592 23588
rect 6736 23604 6788 23656
rect 7472 23672 7524 23724
rect 8208 23740 8260 23792
rect 12348 23740 12400 23792
rect 12716 23808 12768 23860
rect 13176 23808 13228 23860
rect 13268 23808 13320 23860
rect 13912 23808 13964 23860
rect 17960 23808 18012 23860
rect 19156 23808 19208 23860
rect 19432 23851 19484 23860
rect 19432 23817 19441 23851
rect 19441 23817 19475 23851
rect 19475 23817 19484 23851
rect 19432 23808 19484 23817
rect 19616 23851 19668 23860
rect 19616 23817 19625 23851
rect 19625 23817 19659 23851
rect 19659 23817 19668 23851
rect 19616 23808 19668 23817
rect 13360 23740 13412 23792
rect 14648 23740 14700 23792
rect 16304 23740 16356 23792
rect 21548 23783 21600 23792
rect 9036 23672 9088 23724
rect 7196 23536 7248 23588
rect 7840 23604 7892 23656
rect 9220 23647 9272 23656
rect 9220 23613 9229 23647
rect 9229 23613 9263 23647
rect 9263 23613 9272 23647
rect 9220 23604 9272 23613
rect 12532 23672 12584 23724
rect 12808 23672 12860 23724
rect 13268 23672 13320 23724
rect 13820 23672 13872 23724
rect 15752 23672 15804 23724
rect 9128 23536 9180 23588
rect 9864 23604 9916 23656
rect 11704 23647 11756 23656
rect 11704 23613 11722 23647
rect 11722 23613 11756 23647
rect 11704 23604 11756 23613
rect 11888 23604 11940 23656
rect 14372 23604 14424 23656
rect 14740 23604 14792 23656
rect 11520 23536 11572 23588
rect 12348 23536 12400 23588
rect 15384 23604 15436 23656
rect 15844 23604 15896 23656
rect 16856 23604 16908 23656
rect 17132 23604 17184 23656
rect 16304 23536 16356 23588
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 2780 23468 2832 23477
rect 2964 23468 3016 23520
rect 7380 23468 7432 23520
rect 8392 23468 8444 23520
rect 10416 23468 10468 23520
rect 11980 23468 12032 23520
rect 13820 23468 13872 23520
rect 14924 23468 14976 23520
rect 15016 23468 15068 23520
rect 15660 23468 15712 23520
rect 17132 23468 17184 23520
rect 21548 23749 21557 23783
rect 21557 23749 21591 23783
rect 21591 23749 21600 23783
rect 21548 23740 21600 23749
rect 23296 23808 23348 23860
rect 24492 23808 24544 23860
rect 27252 23808 27304 23860
rect 20444 23672 20496 23724
rect 20996 23672 21048 23724
rect 18144 23647 18196 23656
rect 18144 23613 18153 23647
rect 18153 23613 18187 23647
rect 18187 23613 18196 23647
rect 18144 23604 18196 23613
rect 17592 23536 17644 23588
rect 17684 23468 17736 23520
rect 19616 23604 19668 23656
rect 20628 23604 20680 23656
rect 20812 23604 20864 23656
rect 23112 23672 23164 23724
rect 22100 23604 22152 23656
rect 24584 23647 24636 23656
rect 20076 23536 20128 23588
rect 19340 23468 19392 23520
rect 22468 23536 22520 23588
rect 22560 23536 22612 23588
rect 23112 23536 23164 23588
rect 24584 23613 24593 23647
rect 24593 23613 24627 23647
rect 24627 23613 24636 23647
rect 24584 23604 24636 23613
rect 27068 23740 27120 23792
rect 27344 23740 27396 23792
rect 25044 23604 25096 23656
rect 25320 23536 25372 23588
rect 28172 23647 28224 23656
rect 28172 23613 28181 23647
rect 28181 23613 28215 23647
rect 28215 23613 28224 23647
rect 28172 23604 28224 23613
rect 29000 23672 29052 23724
rect 22284 23468 22336 23520
rect 26056 23536 26108 23588
rect 27160 23536 27212 23588
rect 28540 23647 28592 23656
rect 28540 23613 28549 23647
rect 28549 23613 28583 23647
rect 28583 23613 28592 23647
rect 28540 23604 28592 23613
rect 28816 23604 28868 23656
rect 30932 23647 30984 23656
rect 30932 23613 30941 23647
rect 30941 23613 30975 23647
rect 30975 23613 30984 23647
rect 30932 23604 30984 23613
rect 26332 23468 26384 23520
rect 26700 23468 26752 23520
rect 28448 23468 28500 23520
rect 28816 23468 28868 23520
rect 11253 23366 11305 23418
rect 11317 23366 11369 23418
rect 11381 23366 11433 23418
rect 11445 23366 11497 23418
rect 11509 23366 11561 23418
rect 21557 23366 21609 23418
rect 21621 23366 21673 23418
rect 21685 23366 21737 23418
rect 21749 23366 21801 23418
rect 21813 23366 21865 23418
rect 2228 23264 2280 23316
rect 2412 23264 2464 23316
rect 4436 23264 4488 23316
rect 6828 23264 6880 23316
rect 7472 23264 7524 23316
rect 8024 23264 8076 23316
rect 12992 23264 13044 23316
rect 16948 23264 17000 23316
rect 18236 23264 18288 23316
rect 18880 23307 18932 23316
rect 18880 23273 18889 23307
rect 18889 23273 18923 23307
rect 18923 23273 18932 23307
rect 18880 23264 18932 23273
rect 19984 23307 20036 23316
rect 19984 23273 19993 23307
rect 19993 23273 20027 23307
rect 20027 23273 20036 23307
rect 19984 23264 20036 23273
rect 1400 23060 1452 23112
rect 2596 23128 2648 23180
rect 5172 23196 5224 23248
rect 3240 23060 3292 23112
rect 6000 23128 6052 23180
rect 7012 23196 7064 23248
rect 7840 23196 7892 23248
rect 8944 23196 8996 23248
rect 20444 23196 20496 23248
rect 6736 23171 6788 23180
rect 6736 23137 6745 23171
rect 6745 23137 6779 23171
rect 6779 23137 6788 23171
rect 6736 23128 6788 23137
rect 6920 23171 6972 23180
rect 6920 23137 6929 23171
rect 6929 23137 6963 23171
rect 6963 23137 6972 23171
rect 6920 23128 6972 23137
rect 7472 23128 7524 23180
rect 8484 23128 8536 23180
rect 9312 23171 9364 23180
rect 9312 23137 9321 23171
rect 9321 23137 9355 23171
rect 9355 23137 9364 23171
rect 9312 23128 9364 23137
rect 9496 23128 9548 23180
rect 10048 23128 10100 23180
rect 12440 23128 12492 23180
rect 8116 23060 8168 23112
rect 8576 23103 8628 23112
rect 4252 22924 4304 22976
rect 5908 22992 5960 23044
rect 6552 22992 6604 23044
rect 5724 22967 5776 22976
rect 5724 22933 5733 22967
rect 5733 22933 5767 22967
rect 5767 22933 5776 22967
rect 5724 22924 5776 22933
rect 6828 22924 6880 22976
rect 8576 23069 8585 23103
rect 8585 23069 8619 23103
rect 8619 23069 8628 23103
rect 8576 23060 8628 23069
rect 10508 22992 10560 23044
rect 8576 22924 8628 22976
rect 12992 23128 13044 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 13820 23171 13872 23180
rect 13820 23137 13854 23171
rect 13854 23137 13872 23171
rect 13820 23128 13872 23137
rect 14372 23128 14424 23180
rect 15384 23171 15436 23180
rect 15384 23137 15393 23171
rect 15393 23137 15427 23171
rect 15427 23137 15436 23171
rect 15384 23128 15436 23137
rect 15568 23171 15620 23180
rect 15568 23137 15577 23171
rect 15577 23137 15611 23171
rect 15611 23137 15620 23171
rect 15568 23128 15620 23137
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 15844 23128 15896 23180
rect 16028 23128 16080 23180
rect 14188 22924 14240 22976
rect 14740 22924 14792 22976
rect 15108 22924 15160 22976
rect 16028 22924 16080 22976
rect 18052 23060 18104 23112
rect 18512 23060 18564 23112
rect 18604 22924 18656 22976
rect 20628 23128 20680 23180
rect 20904 23264 20956 23316
rect 22560 23307 22612 23316
rect 21272 23171 21324 23180
rect 21272 23137 21281 23171
rect 21281 23137 21315 23171
rect 21315 23137 21324 23171
rect 21272 23128 21324 23137
rect 21824 23171 21876 23180
rect 21824 23137 21833 23171
rect 21833 23137 21867 23171
rect 21867 23137 21876 23171
rect 21824 23128 21876 23137
rect 22008 23171 22060 23180
rect 22008 23137 22017 23171
rect 22017 23137 22051 23171
rect 22051 23137 22060 23171
rect 22008 23128 22060 23137
rect 22560 23273 22569 23307
rect 22569 23273 22603 23307
rect 22603 23273 22612 23307
rect 22560 23264 22612 23273
rect 24952 23307 25004 23316
rect 24952 23273 24961 23307
rect 24961 23273 24995 23307
rect 24995 23273 25004 23307
rect 24952 23264 25004 23273
rect 25228 23264 25280 23316
rect 26516 23264 26568 23316
rect 30288 23307 30340 23316
rect 24492 23196 24544 23248
rect 30288 23273 30297 23307
rect 30297 23273 30331 23307
rect 30331 23273 30340 23307
rect 30288 23264 30340 23273
rect 31116 23264 31168 23316
rect 22744 23128 22796 23180
rect 24400 23128 24452 23180
rect 25780 23128 25832 23180
rect 30196 23196 30248 23248
rect 23296 23060 23348 23112
rect 27160 23060 27212 23112
rect 27252 23060 27304 23112
rect 28632 23128 28684 23180
rect 31024 23128 31076 23180
rect 31300 23128 31352 23180
rect 28724 23060 28776 23112
rect 21824 22992 21876 23044
rect 22008 22992 22060 23044
rect 23112 22992 23164 23044
rect 26700 22992 26752 23044
rect 27436 22992 27488 23044
rect 20904 22924 20956 22976
rect 26056 22967 26108 22976
rect 26056 22933 26065 22967
rect 26065 22933 26099 22967
rect 26099 22933 26108 22967
rect 26056 22924 26108 22933
rect 27252 22924 27304 22976
rect 6102 22822 6154 22874
rect 6166 22822 6218 22874
rect 6230 22822 6282 22874
rect 6294 22822 6346 22874
rect 6358 22822 6410 22874
rect 16405 22822 16457 22874
rect 16469 22822 16521 22874
rect 16533 22822 16585 22874
rect 16597 22822 16649 22874
rect 16661 22822 16713 22874
rect 26709 22822 26761 22874
rect 26773 22822 26825 22874
rect 26837 22822 26889 22874
rect 26901 22822 26953 22874
rect 26965 22822 27017 22874
rect 1952 22720 2004 22772
rect 2596 22763 2648 22772
rect 2596 22729 2605 22763
rect 2605 22729 2639 22763
rect 2639 22729 2648 22763
rect 2596 22720 2648 22729
rect 5172 22720 5224 22772
rect 5908 22763 5960 22772
rect 5908 22729 5917 22763
rect 5917 22729 5951 22763
rect 5951 22729 5960 22763
rect 5908 22720 5960 22729
rect 9312 22720 9364 22772
rect 10048 22763 10100 22772
rect 10048 22729 10057 22763
rect 10057 22729 10091 22763
rect 10091 22729 10100 22763
rect 10048 22720 10100 22729
rect 5632 22652 5684 22704
rect 6736 22652 6788 22704
rect 6276 22584 6328 22636
rect 6552 22584 6604 22636
rect 7564 22584 7616 22636
rect 2044 22559 2096 22568
rect 2044 22525 2057 22559
rect 2057 22525 2091 22559
rect 2091 22525 2096 22559
rect 2044 22516 2096 22525
rect 2139 22559 2191 22568
rect 2139 22525 2154 22559
rect 2154 22525 2188 22559
rect 2188 22525 2191 22559
rect 2412 22559 2464 22568
rect 2139 22516 2191 22525
rect 2412 22525 2421 22559
rect 2421 22525 2455 22559
rect 2455 22525 2464 22559
rect 2412 22516 2464 22525
rect 4252 22516 4304 22568
rect 4620 22559 4672 22568
rect 4620 22525 4629 22559
rect 4629 22525 4663 22559
rect 4663 22525 4672 22559
rect 4620 22516 4672 22525
rect 5448 22516 5500 22568
rect 6000 22516 6052 22568
rect 6460 22516 6512 22568
rect 6920 22516 6972 22568
rect 7656 22516 7708 22568
rect 2228 22380 2280 22432
rect 4160 22380 4212 22432
rect 4804 22380 4856 22432
rect 7748 22448 7800 22500
rect 8484 22652 8536 22704
rect 9128 22652 9180 22704
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 9680 22652 9732 22704
rect 9956 22584 10008 22636
rect 8760 22516 8812 22568
rect 9772 22516 9824 22568
rect 10232 22516 10284 22568
rect 10876 22720 10928 22772
rect 11060 22584 11112 22636
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 12716 22720 12768 22772
rect 13360 22720 13412 22772
rect 13544 22720 13596 22772
rect 19524 22720 19576 22772
rect 19708 22720 19760 22772
rect 18420 22652 18472 22704
rect 21364 22720 21416 22772
rect 14924 22584 14976 22636
rect 18696 22584 18748 22636
rect 22100 22720 22152 22772
rect 22376 22720 22428 22772
rect 22928 22720 22980 22772
rect 23112 22763 23164 22772
rect 23112 22729 23121 22763
rect 23121 22729 23155 22763
rect 23155 22729 23164 22763
rect 23112 22720 23164 22729
rect 24860 22720 24912 22772
rect 25044 22720 25096 22772
rect 26608 22720 26660 22772
rect 26424 22652 26476 22704
rect 27528 22652 27580 22704
rect 28724 22652 28776 22704
rect 10968 22516 11020 22525
rect 11612 22516 11664 22568
rect 11888 22516 11940 22568
rect 15292 22516 15344 22568
rect 15752 22559 15804 22568
rect 15752 22525 15761 22559
rect 15761 22525 15795 22559
rect 15795 22525 15804 22559
rect 15752 22516 15804 22525
rect 16028 22559 16080 22568
rect 16028 22525 16062 22559
rect 16062 22525 16080 22559
rect 16028 22516 16080 22525
rect 17500 22516 17552 22568
rect 17960 22559 18012 22568
rect 17960 22525 17969 22559
rect 17969 22525 18003 22559
rect 18003 22525 18012 22559
rect 17960 22516 18012 22525
rect 18420 22559 18472 22568
rect 18420 22525 18429 22559
rect 18429 22525 18463 22559
rect 18463 22525 18472 22559
rect 18420 22516 18472 22525
rect 26240 22516 26292 22568
rect 15844 22448 15896 22500
rect 16304 22448 16356 22500
rect 19800 22448 19852 22500
rect 7104 22380 7156 22432
rect 7564 22423 7616 22432
rect 7564 22389 7573 22423
rect 7573 22389 7607 22423
rect 7607 22389 7616 22423
rect 7564 22380 7616 22389
rect 7656 22380 7708 22432
rect 8024 22380 8076 22432
rect 8300 22380 8352 22432
rect 9588 22380 9640 22432
rect 13360 22380 13412 22432
rect 15292 22380 15344 22432
rect 15476 22380 15528 22432
rect 17316 22380 17368 22432
rect 19432 22380 19484 22432
rect 21272 22448 21324 22500
rect 25136 22448 25188 22500
rect 28448 22627 28500 22636
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 28448 22584 28500 22593
rect 28540 22627 28592 22636
rect 28540 22593 28549 22627
rect 28549 22593 28583 22627
rect 28583 22593 28592 22627
rect 30932 22627 30984 22636
rect 28540 22584 28592 22593
rect 30932 22593 30941 22627
rect 30941 22593 30975 22627
rect 30975 22593 30984 22627
rect 30932 22584 30984 22593
rect 26884 22559 26936 22568
rect 26884 22525 26893 22559
rect 26893 22525 26927 22559
rect 26927 22525 26936 22559
rect 26884 22516 26936 22525
rect 27068 22559 27120 22568
rect 27068 22525 27077 22559
rect 27077 22525 27111 22559
rect 27111 22525 27120 22559
rect 27252 22559 27304 22568
rect 27068 22516 27120 22525
rect 27252 22525 27261 22559
rect 27261 22525 27295 22559
rect 27295 22525 27304 22559
rect 27252 22516 27304 22525
rect 28172 22559 28224 22568
rect 28172 22525 28181 22559
rect 28181 22525 28215 22559
rect 28215 22525 28224 22559
rect 28172 22516 28224 22525
rect 28724 22559 28776 22568
rect 28264 22448 28316 22500
rect 28724 22525 28733 22559
rect 28733 22525 28767 22559
rect 28767 22525 28776 22559
rect 28724 22516 28776 22525
rect 28816 22448 28868 22500
rect 29368 22380 29420 22432
rect 11253 22278 11305 22330
rect 11317 22278 11369 22330
rect 11381 22278 11433 22330
rect 11445 22278 11497 22330
rect 11509 22278 11561 22330
rect 21557 22278 21609 22330
rect 21621 22278 21673 22330
rect 21685 22278 21737 22330
rect 21749 22278 21801 22330
rect 21813 22278 21865 22330
rect 7472 22176 7524 22228
rect 7656 22176 7708 22228
rect 9496 22176 9548 22228
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 1676 22083 1728 22092
rect 1676 22049 1710 22083
rect 1710 22049 1728 22083
rect 3240 22083 3292 22092
rect 1676 22040 1728 22049
rect 3240 22049 3249 22083
rect 3249 22049 3283 22083
rect 3283 22049 3292 22083
rect 3240 22040 3292 22049
rect 3424 22083 3476 22092
rect 3424 22049 3433 22083
rect 3433 22049 3467 22083
rect 3467 22049 3476 22083
rect 3424 22040 3476 22049
rect 3608 22083 3660 22092
rect 3608 22049 3617 22083
rect 3617 22049 3651 22083
rect 3651 22049 3660 22083
rect 3608 22040 3660 22049
rect 4068 22040 4120 22092
rect 5264 22040 5316 22092
rect 5724 22040 5776 22092
rect 5908 22108 5960 22160
rect 6828 22083 6880 22092
rect 4436 21972 4488 22024
rect 6828 22049 6862 22083
rect 6862 22049 6880 22083
rect 6828 22040 6880 22049
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 8944 21972 8996 22024
rect 2320 21836 2372 21888
rect 4436 21879 4488 21888
rect 4436 21845 4445 21879
rect 4445 21845 4479 21879
rect 4479 21845 4488 21879
rect 4436 21836 4488 21845
rect 5908 21904 5960 21956
rect 6276 21904 6328 21956
rect 9128 21904 9180 21956
rect 9956 22040 10008 22092
rect 10232 22083 10284 22092
rect 10232 22049 10241 22083
rect 10241 22049 10275 22083
rect 10275 22049 10284 22083
rect 10232 22040 10284 22049
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 11060 22176 11112 22228
rect 15844 22176 15896 22228
rect 19248 22176 19300 22228
rect 20996 22219 21048 22228
rect 11152 22108 11204 22160
rect 11612 22040 11664 22092
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 13452 22083 13504 22092
rect 13452 22049 13461 22083
rect 13461 22049 13495 22083
rect 13495 22049 13504 22083
rect 16304 22108 16356 22160
rect 13452 22040 13504 22049
rect 16212 22040 16264 22092
rect 16856 22040 16908 22092
rect 5816 21836 5868 21888
rect 7748 21836 7800 21888
rect 8852 21836 8904 21888
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 11060 21972 11112 22024
rect 15568 21972 15620 22024
rect 16488 21972 16540 22024
rect 17224 22040 17276 22092
rect 17316 22083 17368 22092
rect 17316 22049 17325 22083
rect 17325 22049 17359 22083
rect 17359 22049 17368 22083
rect 17500 22083 17552 22092
rect 17316 22040 17368 22049
rect 17500 22049 17509 22083
rect 17509 22049 17543 22083
rect 17543 22049 17552 22083
rect 17500 22040 17552 22049
rect 19340 22108 19392 22160
rect 18604 22083 18656 22092
rect 18604 22049 18613 22083
rect 18613 22049 18647 22083
rect 18647 22049 18656 22083
rect 18604 22040 18656 22049
rect 20996 22185 21005 22219
rect 21005 22185 21039 22219
rect 21039 22185 21048 22219
rect 20996 22176 21048 22185
rect 22100 22176 22152 22228
rect 23296 22176 23348 22228
rect 24952 22176 25004 22228
rect 25136 22219 25188 22228
rect 25136 22185 25145 22219
rect 25145 22185 25179 22219
rect 25179 22185 25188 22219
rect 25136 22176 25188 22185
rect 26424 22219 26476 22228
rect 26424 22185 26433 22219
rect 26433 22185 26467 22219
rect 26467 22185 26476 22219
rect 26424 22176 26476 22185
rect 27160 22176 27212 22228
rect 19892 22083 19944 22092
rect 19892 22049 19926 22083
rect 19926 22049 19944 22083
rect 23020 22108 23072 22160
rect 19892 22040 19944 22049
rect 22100 22040 22152 22092
rect 18052 21972 18104 22024
rect 17960 21904 18012 21956
rect 18788 22015 18840 22024
rect 18788 21981 18797 22015
rect 18797 21981 18831 22015
rect 18831 21981 18840 22015
rect 19616 22015 19668 22024
rect 18788 21972 18840 21981
rect 19616 21981 19625 22015
rect 19625 21981 19659 22015
rect 19659 21981 19668 22015
rect 19616 21972 19668 21981
rect 25964 22108 26016 22160
rect 26332 22108 26384 22160
rect 25044 22040 25096 22092
rect 27528 22040 27580 22092
rect 28172 22040 28224 22092
rect 28724 22108 28776 22160
rect 28632 22083 28684 22092
rect 22284 21972 22336 22024
rect 23848 21972 23900 22024
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 28356 22015 28408 22024
rect 24768 21972 24820 21981
rect 28356 21981 28365 22015
rect 28365 21981 28399 22015
rect 28399 21981 28408 22015
rect 28356 21972 28408 21981
rect 28632 22049 28641 22083
rect 28641 22049 28675 22083
rect 28675 22049 28684 22083
rect 28632 22040 28684 22049
rect 28540 21972 28592 22024
rect 24860 21904 24912 21956
rect 26056 21904 26108 21956
rect 28172 21904 28224 21956
rect 28724 21904 28776 21956
rect 29368 22083 29420 22092
rect 29368 22049 29377 22083
rect 29377 22049 29411 22083
rect 29411 22049 29420 22083
rect 29368 22040 29420 22049
rect 31300 22083 31352 22092
rect 11888 21836 11940 21888
rect 12440 21836 12492 21888
rect 19892 21836 19944 21888
rect 20352 21836 20404 21888
rect 23664 21836 23716 21888
rect 23940 21836 23992 21888
rect 27068 21836 27120 21888
rect 28816 21879 28868 21888
rect 28816 21845 28825 21879
rect 28825 21845 28859 21879
rect 28859 21845 28868 21879
rect 28816 21836 28868 21845
rect 28908 21836 28960 21888
rect 31300 22049 31309 22083
rect 31309 22049 31343 22083
rect 31343 22049 31352 22083
rect 31300 22040 31352 22049
rect 6102 21734 6154 21786
rect 6166 21734 6218 21786
rect 6230 21734 6282 21786
rect 6294 21734 6346 21786
rect 6358 21734 6410 21786
rect 16405 21734 16457 21786
rect 16469 21734 16521 21786
rect 16533 21734 16585 21786
rect 16597 21734 16649 21786
rect 16661 21734 16713 21786
rect 26709 21734 26761 21786
rect 26773 21734 26825 21786
rect 26837 21734 26889 21786
rect 26901 21734 26953 21786
rect 26965 21734 27017 21786
rect 1676 21632 1728 21684
rect 2412 21632 2464 21684
rect 4620 21632 4672 21684
rect 4712 21675 4764 21684
rect 4712 21641 4721 21675
rect 4721 21641 4755 21675
rect 4755 21641 4764 21675
rect 5264 21675 5316 21684
rect 4712 21632 4764 21641
rect 5264 21641 5273 21675
rect 5273 21641 5307 21675
rect 5307 21641 5316 21675
rect 5264 21632 5316 21641
rect 8576 21632 8628 21684
rect 13176 21632 13228 21684
rect 13636 21632 13688 21684
rect 14464 21675 14516 21684
rect 14464 21641 14473 21675
rect 14473 21641 14507 21675
rect 14507 21641 14516 21675
rect 14464 21632 14516 21641
rect 5816 21564 5868 21616
rect 8944 21564 8996 21616
rect 11980 21564 12032 21616
rect 18144 21632 18196 21684
rect 18328 21632 18380 21684
rect 19432 21675 19484 21684
rect 19432 21641 19441 21675
rect 19441 21641 19475 21675
rect 19475 21641 19484 21675
rect 19432 21632 19484 21641
rect 1952 21539 2004 21548
rect 1952 21505 1961 21539
rect 1961 21505 1995 21539
rect 1995 21505 2004 21539
rect 1952 21496 2004 21505
rect 2044 21471 2096 21480
rect 2044 21437 2053 21471
rect 2053 21437 2087 21471
rect 2087 21437 2096 21471
rect 2044 21428 2096 21437
rect 2504 21496 2556 21548
rect 4804 21496 4856 21548
rect 5080 21496 5132 21548
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 6552 21496 6604 21548
rect 9128 21496 9180 21548
rect 9312 21496 9364 21548
rect 9588 21496 9640 21548
rect 10140 21496 10192 21548
rect 10600 21496 10652 21548
rect 10968 21496 11020 21548
rect 2228 21428 2280 21480
rect 3608 21428 3660 21480
rect 3792 21428 3844 21480
rect 4436 21428 4488 21480
rect 5448 21471 5500 21480
rect 5448 21437 5457 21471
rect 5457 21437 5491 21471
rect 5491 21437 5500 21471
rect 5448 21428 5500 21437
rect 5816 21471 5868 21480
rect 5816 21437 5825 21471
rect 5825 21437 5859 21471
rect 5859 21437 5868 21471
rect 5816 21428 5868 21437
rect 6000 21471 6052 21480
rect 6000 21437 6009 21471
rect 6009 21437 6043 21471
rect 6043 21437 6052 21471
rect 6000 21428 6052 21437
rect 6460 21428 6512 21480
rect 7564 21428 7616 21480
rect 10232 21471 10284 21480
rect 10232 21437 10241 21471
rect 10241 21437 10275 21471
rect 10275 21437 10284 21471
rect 10232 21428 10284 21437
rect 10876 21428 10928 21480
rect 13268 21496 13320 21548
rect 14924 21539 14976 21548
rect 11704 21428 11756 21480
rect 12900 21428 12952 21480
rect 13360 21428 13412 21480
rect 2412 21360 2464 21412
rect 3056 21292 3108 21344
rect 4896 21360 4948 21412
rect 9128 21360 9180 21412
rect 9864 21360 9916 21412
rect 12164 21360 12216 21412
rect 13636 21360 13688 21412
rect 3332 21292 3384 21344
rect 3884 21292 3936 21344
rect 4620 21292 4672 21344
rect 7196 21292 7248 21344
rect 7656 21292 7708 21344
rect 8392 21335 8444 21344
rect 8392 21301 8401 21335
rect 8401 21301 8435 21335
rect 8435 21301 8444 21335
rect 8392 21292 8444 21301
rect 13084 21292 13136 21344
rect 13268 21292 13320 21344
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 14372 21428 14424 21480
rect 15016 21471 15068 21480
rect 15016 21437 15021 21471
rect 15021 21437 15055 21471
rect 15055 21437 15068 21471
rect 15016 21428 15068 21437
rect 15384 21496 15436 21548
rect 15568 21496 15620 21548
rect 15476 21428 15528 21480
rect 15752 21471 15804 21480
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 17684 21496 17736 21548
rect 18328 21496 18380 21548
rect 18788 21496 18840 21548
rect 19984 21564 20036 21616
rect 21456 21632 21508 21684
rect 22192 21632 22244 21684
rect 22468 21632 22520 21684
rect 23940 21632 23992 21684
rect 24400 21675 24452 21684
rect 24400 21641 24409 21675
rect 24409 21641 24443 21675
rect 24443 21641 24452 21675
rect 24400 21632 24452 21641
rect 25320 21632 25372 21684
rect 27528 21632 27580 21684
rect 16396 21428 16448 21480
rect 16580 21428 16632 21480
rect 14464 21292 14516 21344
rect 16856 21360 16908 21412
rect 15660 21292 15712 21344
rect 16948 21292 17000 21344
rect 17132 21335 17184 21344
rect 17132 21301 17141 21335
rect 17141 21301 17175 21335
rect 17175 21301 17184 21335
rect 17132 21292 17184 21301
rect 18604 21428 18656 21480
rect 19708 21428 19760 21480
rect 21088 21496 21140 21548
rect 22100 21496 22152 21548
rect 24400 21496 24452 21548
rect 23664 21471 23716 21480
rect 18512 21403 18564 21412
rect 18512 21369 18521 21403
rect 18521 21369 18555 21403
rect 18555 21369 18564 21403
rect 18512 21360 18564 21369
rect 19340 21360 19392 21412
rect 20168 21360 20220 21412
rect 20260 21292 20312 21344
rect 20812 21292 20864 21344
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 24952 21564 25004 21616
rect 25780 21564 25832 21616
rect 28448 21564 28500 21616
rect 24860 21471 24912 21480
rect 24860 21437 24869 21471
rect 24869 21437 24903 21471
rect 24903 21437 24912 21471
rect 24860 21428 24912 21437
rect 24952 21471 25004 21480
rect 24952 21437 24961 21471
rect 24961 21437 24995 21471
rect 24995 21437 25004 21471
rect 24952 21428 25004 21437
rect 25136 21471 25188 21480
rect 25136 21437 25145 21471
rect 25145 21437 25179 21471
rect 25179 21437 25188 21471
rect 25136 21428 25188 21437
rect 23572 21360 23624 21412
rect 25504 21292 25556 21344
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 27528 21471 27580 21480
rect 26056 21360 26108 21412
rect 27528 21437 27537 21471
rect 27537 21437 27571 21471
rect 27571 21437 27580 21471
rect 27528 21428 27580 21437
rect 28172 21471 28224 21480
rect 28172 21437 28181 21471
rect 28181 21437 28215 21471
rect 28215 21437 28224 21471
rect 28172 21428 28224 21437
rect 28448 21471 28500 21480
rect 28448 21437 28457 21471
rect 28457 21437 28491 21471
rect 28491 21437 28500 21471
rect 28448 21428 28500 21437
rect 28540 21471 28592 21480
rect 28540 21437 28549 21471
rect 28549 21437 28583 21471
rect 28583 21437 28592 21471
rect 29460 21632 29512 21684
rect 31300 21632 31352 21684
rect 31024 21564 31076 21616
rect 30656 21496 30708 21548
rect 31392 21496 31444 21548
rect 31576 21496 31628 21548
rect 28540 21428 28592 21437
rect 30840 21428 30892 21480
rect 30288 21403 30340 21412
rect 30288 21369 30297 21403
rect 30297 21369 30331 21403
rect 30331 21369 30340 21403
rect 30288 21360 30340 21369
rect 31208 21428 31260 21480
rect 31576 21360 31628 21412
rect 26332 21335 26384 21344
rect 26332 21301 26341 21335
rect 26341 21301 26375 21335
rect 26375 21301 26384 21335
rect 26332 21292 26384 21301
rect 26608 21292 26660 21344
rect 27988 21335 28040 21344
rect 27988 21301 27997 21335
rect 27997 21301 28031 21335
rect 28031 21301 28040 21335
rect 27988 21292 28040 21301
rect 28080 21292 28132 21344
rect 30472 21292 30524 21344
rect 31208 21292 31260 21344
rect 11253 21190 11305 21242
rect 11317 21190 11369 21242
rect 11381 21190 11433 21242
rect 11445 21190 11497 21242
rect 11509 21190 11561 21242
rect 21557 21190 21609 21242
rect 21621 21190 21673 21242
rect 21685 21190 21737 21242
rect 21749 21190 21801 21242
rect 21813 21190 21865 21242
rect 3424 21088 3476 21140
rect 6736 21088 6788 21140
rect 7288 21088 7340 21140
rect 8300 21088 8352 21140
rect 9128 21088 9180 21140
rect 12900 21131 12952 21140
rect 12900 21097 12909 21131
rect 12909 21097 12943 21131
rect 12943 21097 12952 21131
rect 12900 21088 12952 21097
rect 1860 21020 1912 21072
rect 2688 21020 2740 21072
rect 2412 20952 2464 21004
rect 3240 21020 3292 21072
rect 3792 21063 3844 21072
rect 3792 21029 3817 21063
rect 3817 21029 3844 21063
rect 3792 21020 3844 21029
rect 5908 21020 5960 21072
rect 7012 21020 7064 21072
rect 16580 21088 16632 21140
rect 16764 21131 16816 21140
rect 16764 21097 16773 21131
rect 16773 21097 16807 21131
rect 16807 21097 16816 21131
rect 16764 21088 16816 21097
rect 18144 21088 18196 21140
rect 21916 21088 21968 21140
rect 3516 20952 3568 21004
rect 3148 20927 3200 20936
rect 3148 20893 3157 20927
rect 3157 20893 3191 20927
rect 3191 20893 3200 20927
rect 3148 20884 3200 20893
rect 3332 20884 3384 20936
rect 3884 20884 3936 20936
rect 4068 20884 4120 20936
rect 4528 20952 4580 21004
rect 6000 20952 6052 21004
rect 8024 20952 8076 21004
rect 8392 20995 8444 21004
rect 8392 20961 8401 20995
rect 8401 20961 8435 20995
rect 8435 20961 8444 20995
rect 8392 20952 8444 20961
rect 8944 20952 8996 21004
rect 9772 20952 9824 21004
rect 10968 20952 11020 21004
rect 11152 20952 11204 21004
rect 11520 20995 11572 21004
rect 11520 20961 11529 20995
rect 11529 20961 11563 20995
rect 11563 20961 11572 20995
rect 11520 20952 11572 20961
rect 12440 20952 12492 21004
rect 13084 20995 13136 21004
rect 13084 20961 13093 20995
rect 13093 20961 13127 20995
rect 13127 20961 13136 20995
rect 13084 20952 13136 20961
rect 13268 20995 13320 21004
rect 13268 20961 13277 20995
rect 13277 20961 13311 20995
rect 13311 20961 13320 20995
rect 13268 20952 13320 20961
rect 13452 20995 13504 21004
rect 13452 20961 13461 20995
rect 13461 20961 13495 20995
rect 13495 20961 13504 20995
rect 13452 20952 13504 20961
rect 14280 20995 14332 21004
rect 4712 20884 4764 20936
rect 5172 20884 5224 20936
rect 5908 20884 5960 20936
rect 9220 20884 9272 20936
rect 1400 20816 1452 20868
rect 2780 20816 2832 20868
rect 4896 20816 4948 20868
rect 9956 20816 10008 20868
rect 11980 20884 12032 20936
rect 13544 20884 13596 20936
rect 12992 20816 13044 20868
rect 14280 20961 14289 20995
rect 14289 20961 14323 20995
rect 14323 20961 14332 20995
rect 14280 20952 14332 20961
rect 14464 20995 14516 21004
rect 14464 20961 14473 20995
rect 14473 20961 14507 20995
rect 14507 20961 14516 20995
rect 14464 20952 14516 20961
rect 14924 21020 14976 21072
rect 15016 21020 15068 21072
rect 15384 20952 15436 21004
rect 15936 20952 15988 21004
rect 17316 21020 17368 21072
rect 16764 20952 16816 21004
rect 17408 20952 17460 21004
rect 18604 20952 18656 21004
rect 18788 20952 18840 21004
rect 20904 20952 20956 21004
rect 15568 20884 15620 20936
rect 15660 20884 15712 20936
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 16120 20927 16172 20936
rect 16120 20893 16129 20927
rect 16129 20893 16163 20927
rect 16163 20893 16172 20927
rect 16120 20884 16172 20893
rect 16212 20884 16264 20936
rect 2320 20791 2372 20800
rect 2320 20757 2329 20791
rect 2329 20757 2363 20791
rect 2363 20757 2372 20791
rect 2320 20748 2372 20757
rect 2964 20791 3016 20800
rect 2964 20757 2973 20791
rect 2973 20757 3007 20791
rect 3007 20757 3016 20791
rect 2964 20748 3016 20757
rect 3332 20748 3384 20800
rect 3884 20748 3936 20800
rect 4160 20748 4212 20800
rect 4436 20748 4488 20800
rect 10876 20748 10928 20800
rect 11980 20748 12032 20800
rect 13544 20748 13596 20800
rect 14372 20748 14424 20800
rect 15108 20748 15160 20800
rect 15660 20748 15712 20800
rect 16396 20816 16448 20868
rect 18512 20884 18564 20936
rect 20076 20884 20128 20936
rect 20168 20884 20220 20936
rect 21364 21020 21416 21072
rect 23112 21020 23164 21072
rect 23848 21088 23900 21140
rect 25136 21088 25188 21140
rect 25872 21088 25924 21140
rect 22560 20952 22612 21004
rect 23296 20952 23348 21004
rect 23664 21020 23716 21072
rect 25964 21020 26016 21072
rect 28540 21088 28592 21140
rect 29552 21088 29604 21140
rect 30748 21131 30800 21140
rect 30748 21097 30757 21131
rect 30757 21097 30791 21131
rect 30791 21097 30800 21131
rect 30748 21088 30800 21097
rect 28816 21020 28868 21072
rect 24032 20952 24084 21004
rect 24308 20952 24360 21004
rect 24768 20952 24820 21004
rect 25780 20952 25832 21004
rect 28356 20952 28408 21004
rect 31024 20995 31076 21004
rect 31024 20961 31033 20995
rect 31033 20961 31067 20995
rect 31067 20961 31076 20995
rect 31024 20952 31076 20961
rect 31208 20995 31260 21004
rect 31208 20961 31217 20995
rect 31217 20961 31251 20995
rect 31251 20961 31260 20995
rect 31208 20952 31260 20961
rect 22468 20927 22520 20936
rect 22468 20893 22477 20927
rect 22477 20893 22511 20927
rect 22511 20893 22520 20927
rect 22468 20884 22520 20893
rect 25596 20927 25648 20936
rect 25596 20893 25605 20927
rect 25605 20893 25639 20927
rect 25639 20893 25648 20927
rect 25596 20884 25648 20893
rect 28080 20884 28132 20936
rect 30380 20884 30432 20936
rect 30840 20884 30892 20936
rect 30932 20927 30984 20936
rect 30932 20893 30941 20927
rect 30941 20893 30975 20927
rect 30975 20893 30984 20927
rect 30932 20884 30984 20893
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 17316 20748 17368 20800
rect 22928 20816 22980 20868
rect 19156 20748 19208 20800
rect 19800 20748 19852 20800
rect 24124 20748 24176 20800
rect 24584 20791 24636 20800
rect 24584 20757 24593 20791
rect 24593 20757 24627 20791
rect 24627 20757 24636 20791
rect 24584 20748 24636 20757
rect 24952 20748 25004 20800
rect 25136 20791 25188 20800
rect 25136 20757 25145 20791
rect 25145 20757 25179 20791
rect 25179 20757 25188 20791
rect 25136 20748 25188 20757
rect 27160 20748 27212 20800
rect 6102 20646 6154 20698
rect 6166 20646 6218 20698
rect 6230 20646 6282 20698
rect 6294 20646 6346 20698
rect 6358 20646 6410 20698
rect 16405 20646 16457 20698
rect 16469 20646 16521 20698
rect 16533 20646 16585 20698
rect 16597 20646 16649 20698
rect 16661 20646 16713 20698
rect 26709 20646 26761 20698
rect 26773 20646 26825 20698
rect 26837 20646 26889 20698
rect 26901 20646 26953 20698
rect 26965 20646 27017 20698
rect 7656 20544 7708 20596
rect 8852 20544 8904 20596
rect 13084 20544 13136 20596
rect 13360 20587 13412 20596
rect 2688 20476 2740 20528
rect 5172 20476 5224 20528
rect 9956 20476 10008 20528
rect 10968 20476 11020 20528
rect 11152 20476 11204 20528
rect 13360 20553 13369 20587
rect 13369 20553 13403 20587
rect 13403 20553 13412 20587
rect 13360 20544 13412 20553
rect 15016 20544 15068 20596
rect 2964 20451 3016 20460
rect 2964 20417 2973 20451
rect 2973 20417 3007 20451
rect 3007 20417 3016 20451
rect 2964 20408 3016 20417
rect 4436 20451 4488 20460
rect 4436 20417 4445 20451
rect 4445 20417 4479 20451
rect 4479 20417 4488 20451
rect 4436 20408 4488 20417
rect 5816 20408 5868 20460
rect 2044 20340 2096 20392
rect 2412 20340 2464 20392
rect 3240 20383 3292 20392
rect 3240 20349 3249 20383
rect 3249 20349 3283 20383
rect 3283 20349 3292 20383
rect 4252 20383 4304 20392
rect 3240 20340 3292 20349
rect 4252 20349 4261 20383
rect 4261 20349 4295 20383
rect 4295 20349 4304 20383
rect 4252 20340 4304 20349
rect 4896 20383 4948 20392
rect 4896 20349 4905 20383
rect 4905 20349 4939 20383
rect 4939 20349 4948 20383
rect 4896 20340 4948 20349
rect 5448 20340 5500 20392
rect 7564 20408 7616 20460
rect 8208 20451 8260 20460
rect 6552 20340 6604 20392
rect 7012 20383 7064 20392
rect 7012 20349 7021 20383
rect 7021 20349 7055 20383
rect 7055 20349 7064 20383
rect 7012 20340 7064 20349
rect 7932 20383 7984 20392
rect 7932 20349 7941 20383
rect 7941 20349 7975 20383
rect 7975 20349 7984 20383
rect 7932 20340 7984 20349
rect 8208 20417 8217 20451
rect 8217 20417 8251 20451
rect 8251 20417 8260 20451
rect 8208 20408 8260 20417
rect 11888 20451 11940 20460
rect 11888 20417 11897 20451
rect 11897 20417 11931 20451
rect 11931 20417 11940 20451
rect 11888 20408 11940 20417
rect 8484 20340 8536 20392
rect 8944 20383 8996 20392
rect 8944 20349 8953 20383
rect 8953 20349 8987 20383
rect 8987 20349 8996 20383
rect 8944 20340 8996 20349
rect 11060 20340 11112 20392
rect 11520 20340 11572 20392
rect 5172 20272 5224 20324
rect 1584 20204 1636 20256
rect 1768 20247 1820 20256
rect 1768 20213 1777 20247
rect 1777 20213 1811 20247
rect 1811 20213 1820 20247
rect 1768 20204 1820 20213
rect 3424 20204 3476 20256
rect 5448 20204 5500 20256
rect 6000 20204 6052 20256
rect 7932 20204 7984 20256
rect 11704 20340 11756 20392
rect 12440 20408 12492 20460
rect 13360 20408 13412 20460
rect 12072 20340 12124 20392
rect 12992 20340 13044 20392
rect 15476 20340 15528 20392
rect 15936 20383 15988 20392
rect 15936 20349 15945 20383
rect 15945 20349 15979 20383
rect 15979 20349 15988 20383
rect 15936 20340 15988 20349
rect 16304 20476 16356 20528
rect 16856 20544 16908 20596
rect 20260 20544 20312 20596
rect 21456 20544 21508 20596
rect 22468 20587 22520 20596
rect 16488 20476 16540 20528
rect 17224 20476 17276 20528
rect 17684 20476 17736 20528
rect 18512 20476 18564 20528
rect 18880 20476 18932 20528
rect 21364 20476 21416 20528
rect 22468 20553 22477 20587
rect 22477 20553 22511 20587
rect 22511 20553 22520 20587
rect 22468 20544 22520 20553
rect 23112 20587 23164 20596
rect 23112 20553 23121 20587
rect 23121 20553 23155 20587
rect 23155 20553 23164 20587
rect 23112 20544 23164 20553
rect 25504 20587 25556 20596
rect 17960 20408 18012 20460
rect 19708 20408 19760 20460
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22100 20408 22152 20417
rect 14372 20315 14424 20324
rect 14372 20281 14406 20315
rect 14406 20281 14424 20315
rect 14372 20272 14424 20281
rect 14464 20272 14516 20324
rect 14832 20272 14884 20324
rect 15384 20272 15436 20324
rect 15844 20272 15896 20324
rect 16580 20340 16632 20392
rect 17224 20340 17276 20392
rect 18512 20383 18564 20392
rect 17592 20272 17644 20324
rect 18512 20349 18521 20383
rect 18521 20349 18555 20383
rect 18555 20349 18564 20383
rect 18512 20340 18564 20349
rect 18880 20272 18932 20324
rect 8852 20204 8904 20256
rect 10416 20204 10468 20256
rect 11612 20204 11664 20256
rect 12716 20204 12768 20256
rect 13268 20204 13320 20256
rect 15108 20204 15160 20256
rect 16672 20204 16724 20256
rect 20168 20340 20220 20392
rect 20904 20383 20956 20392
rect 20904 20349 20913 20383
rect 20913 20349 20947 20383
rect 20947 20349 20956 20383
rect 20904 20340 20956 20349
rect 21088 20383 21140 20392
rect 21088 20349 21097 20383
rect 21097 20349 21131 20383
rect 21131 20349 21140 20383
rect 21088 20340 21140 20349
rect 21916 20383 21968 20392
rect 21916 20349 21925 20383
rect 21925 20349 21959 20383
rect 21959 20349 21968 20383
rect 21916 20340 21968 20349
rect 24584 20476 24636 20528
rect 25504 20553 25513 20587
rect 25513 20553 25547 20587
rect 25547 20553 25556 20587
rect 25504 20544 25556 20553
rect 28724 20587 28776 20596
rect 28724 20553 28733 20587
rect 28733 20553 28767 20587
rect 28767 20553 28776 20587
rect 28724 20544 28776 20553
rect 31668 20544 31720 20596
rect 30196 20476 30248 20528
rect 23388 20408 23440 20460
rect 30472 20451 30524 20460
rect 30472 20417 30481 20451
rect 30481 20417 30515 20451
rect 30515 20417 30524 20451
rect 30472 20408 30524 20417
rect 30656 20451 30708 20460
rect 30656 20417 30665 20451
rect 30665 20417 30699 20451
rect 30699 20417 30708 20451
rect 30656 20408 30708 20417
rect 21180 20272 21232 20324
rect 22008 20272 22060 20324
rect 23664 20383 23716 20392
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 23848 20383 23900 20392
rect 23848 20349 23857 20383
rect 23857 20349 23891 20383
rect 23891 20349 23900 20383
rect 23848 20340 23900 20349
rect 24768 20340 24820 20392
rect 26240 20340 26292 20392
rect 27988 20340 28040 20392
rect 28724 20340 28776 20392
rect 30288 20340 30340 20392
rect 25136 20272 25188 20324
rect 26608 20315 26660 20324
rect 26608 20281 26626 20315
rect 26626 20281 26660 20315
rect 26608 20272 26660 20281
rect 30472 20272 30524 20324
rect 30932 20340 30984 20392
rect 20812 20204 20864 20256
rect 21272 20247 21324 20256
rect 21272 20213 21281 20247
rect 21281 20213 21315 20247
rect 21315 20213 21324 20247
rect 21272 20204 21324 20213
rect 21364 20204 21416 20256
rect 24952 20247 25004 20256
rect 24952 20213 24961 20247
rect 24961 20213 24995 20247
rect 24995 20213 25004 20247
rect 24952 20204 25004 20213
rect 11253 20102 11305 20154
rect 11317 20102 11369 20154
rect 11381 20102 11433 20154
rect 11445 20102 11497 20154
rect 11509 20102 11561 20154
rect 21557 20102 21609 20154
rect 21621 20102 21673 20154
rect 21685 20102 21737 20154
rect 21749 20102 21801 20154
rect 21813 20102 21865 20154
rect 1308 20000 1360 20052
rect 1492 20000 1544 20052
rect 2964 20043 3016 20052
rect 2964 20009 2973 20043
rect 2973 20009 3007 20043
rect 3007 20009 3016 20043
rect 2964 20000 3016 20009
rect 4252 20043 4304 20052
rect 4252 20009 4261 20043
rect 4261 20009 4295 20043
rect 4295 20009 4304 20043
rect 4252 20000 4304 20009
rect 5356 20000 5408 20052
rect 8208 20043 8260 20052
rect 1492 19907 1544 19916
rect 1492 19873 1501 19907
rect 1501 19873 1535 19907
rect 1535 19873 1544 19907
rect 1492 19864 1544 19873
rect 1676 19864 1728 19916
rect 2412 19932 2464 19984
rect 4620 19932 4672 19984
rect 4896 19932 4948 19984
rect 8208 20009 8217 20043
rect 8217 20009 8251 20043
rect 8251 20009 8260 20043
rect 8208 20000 8260 20009
rect 10508 20000 10560 20052
rect 10968 20000 11020 20052
rect 12624 20000 12676 20052
rect 13452 20043 13504 20052
rect 2504 19907 2556 19916
rect 2504 19873 2513 19907
rect 2513 19873 2547 19907
rect 2547 19873 2556 19907
rect 2504 19864 2556 19873
rect 3424 19907 3476 19916
rect 3424 19873 3433 19907
rect 3433 19873 3467 19907
rect 3467 19873 3476 19907
rect 3424 19864 3476 19873
rect 3608 19907 3660 19916
rect 3608 19873 3617 19907
rect 3617 19873 3651 19907
rect 3651 19873 3660 19907
rect 3608 19864 3660 19873
rect 4160 19907 4212 19916
rect 4160 19873 4169 19907
rect 4169 19873 4203 19907
rect 4203 19873 4212 19907
rect 4160 19864 4212 19873
rect 7656 19932 7708 19984
rect 1768 19703 1820 19712
rect 1768 19669 1777 19703
rect 1777 19669 1811 19703
rect 1811 19669 1820 19703
rect 1768 19660 1820 19669
rect 2872 19728 2924 19780
rect 6552 19907 6604 19916
rect 5172 19796 5224 19848
rect 6552 19873 6561 19907
rect 6561 19873 6595 19907
rect 6595 19873 6604 19907
rect 6552 19864 6604 19873
rect 7748 19907 7800 19916
rect 5264 19728 5316 19780
rect 6000 19728 6052 19780
rect 7748 19873 7757 19907
rect 7757 19873 7791 19907
rect 7791 19873 7800 19907
rect 7748 19864 7800 19873
rect 8024 19932 8076 19984
rect 7932 19907 7984 19916
rect 7932 19873 7941 19907
rect 7941 19873 7975 19907
rect 7975 19873 7984 19907
rect 7932 19864 7984 19873
rect 9128 19864 9180 19916
rect 10416 19907 10468 19916
rect 10416 19873 10425 19907
rect 10425 19873 10459 19907
rect 10459 19873 10468 19907
rect 10416 19864 10468 19873
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 12900 19932 12952 19984
rect 13452 20009 13461 20043
rect 13461 20009 13495 20043
rect 13495 20009 13504 20043
rect 13452 20000 13504 20009
rect 14188 20000 14240 20052
rect 14832 20000 14884 20052
rect 18972 20000 19024 20052
rect 13360 19907 13412 19916
rect 8116 19796 8168 19848
rect 8484 19728 8536 19780
rect 13360 19873 13369 19907
rect 13369 19873 13403 19907
rect 13403 19873 13412 19907
rect 13360 19864 13412 19873
rect 14280 19864 14332 19916
rect 15108 19864 15160 19916
rect 15384 19907 15436 19916
rect 15384 19873 15393 19907
rect 15393 19873 15427 19907
rect 15427 19873 15436 19907
rect 15384 19864 15436 19873
rect 16120 19932 16172 19984
rect 17684 19932 17736 19984
rect 21180 20000 21232 20052
rect 23664 20000 23716 20052
rect 26148 20000 26200 20052
rect 31116 20000 31168 20052
rect 22100 19932 22152 19984
rect 26332 19932 26384 19984
rect 13176 19796 13228 19848
rect 15844 19864 15896 19916
rect 15292 19728 15344 19780
rect 15844 19728 15896 19780
rect 16212 19864 16264 19916
rect 16580 19864 16632 19916
rect 17132 19864 17184 19916
rect 18604 19907 18656 19916
rect 3332 19660 3384 19712
rect 4988 19703 5040 19712
rect 4988 19669 4997 19703
rect 4997 19669 5031 19703
rect 5031 19669 5040 19703
rect 4988 19660 5040 19669
rect 6828 19660 6880 19712
rect 7012 19703 7064 19712
rect 7012 19669 7021 19703
rect 7021 19669 7055 19703
rect 7055 19669 7064 19703
rect 7012 19660 7064 19669
rect 8576 19660 8628 19712
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 9404 19660 9456 19712
rect 9772 19660 9824 19712
rect 11152 19660 11204 19712
rect 13820 19660 13872 19712
rect 16672 19796 16724 19848
rect 18144 19839 18196 19848
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 18972 19907 19024 19916
rect 18972 19873 18981 19907
rect 18981 19873 19015 19907
rect 19015 19873 19024 19907
rect 18972 19864 19024 19873
rect 16856 19728 16908 19780
rect 18696 19728 18748 19780
rect 17408 19660 17460 19712
rect 19616 19864 19668 19916
rect 20904 19864 20956 19916
rect 22284 19864 22336 19916
rect 22468 19907 22520 19916
rect 22468 19873 22502 19907
rect 22502 19873 22520 19907
rect 27528 19907 27580 19916
rect 22468 19864 22520 19873
rect 27528 19873 27537 19907
rect 27537 19873 27571 19907
rect 27571 19873 27580 19907
rect 27528 19864 27580 19873
rect 28080 19864 28132 19916
rect 31024 19932 31076 19984
rect 26240 19796 26292 19848
rect 19156 19660 19208 19712
rect 21364 19660 21416 19712
rect 23296 19660 23348 19712
rect 24400 19660 24452 19712
rect 28908 19796 28960 19848
rect 30748 19864 30800 19916
rect 31392 19932 31444 19984
rect 31300 19907 31352 19916
rect 31300 19873 31309 19907
rect 31309 19873 31343 19907
rect 31343 19873 31352 19907
rect 31300 19864 31352 19873
rect 28356 19703 28408 19712
rect 28356 19669 28365 19703
rect 28365 19669 28399 19703
rect 28399 19669 28408 19703
rect 28356 19660 28408 19669
rect 29920 19660 29972 19712
rect 6102 19558 6154 19610
rect 6166 19558 6218 19610
rect 6230 19558 6282 19610
rect 6294 19558 6346 19610
rect 6358 19558 6410 19610
rect 16405 19558 16457 19610
rect 16469 19558 16521 19610
rect 16533 19558 16585 19610
rect 16597 19558 16649 19610
rect 16661 19558 16713 19610
rect 26709 19558 26761 19610
rect 26773 19558 26825 19610
rect 26837 19558 26889 19610
rect 26901 19558 26953 19610
rect 26965 19558 27017 19610
rect 1768 19456 1820 19508
rect 2688 19456 2740 19508
rect 3608 19456 3660 19508
rect 7012 19456 7064 19508
rect 7288 19456 7340 19508
rect 12440 19456 12492 19508
rect 1492 19388 1544 19440
rect 2412 19388 2464 19440
rect 2780 19388 2832 19440
rect 3424 19388 3476 19440
rect 3884 19363 3936 19372
rect 2044 19252 2096 19304
rect 2320 19252 2372 19304
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 4620 19388 4672 19440
rect 5172 19388 5224 19440
rect 5448 19388 5500 19440
rect 4252 19320 4304 19372
rect 8024 19363 8076 19372
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 8392 19363 8444 19372
rect 8392 19329 8401 19363
rect 8401 19329 8435 19363
rect 8435 19329 8444 19363
rect 8392 19320 8444 19329
rect 9404 19320 9456 19372
rect 9772 19363 9824 19372
rect 9772 19329 9781 19363
rect 9781 19329 9815 19363
rect 9815 19329 9824 19363
rect 9772 19320 9824 19329
rect 2872 19252 2924 19261
rect 3424 19252 3476 19304
rect 4436 19252 4488 19304
rect 5632 19295 5684 19304
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 6000 19295 6052 19304
rect 6000 19261 6009 19295
rect 6009 19261 6043 19295
rect 6043 19261 6052 19295
rect 6000 19252 6052 19261
rect 6736 19252 6788 19304
rect 7656 19295 7708 19304
rect 3148 19227 3200 19236
rect 3148 19193 3157 19227
rect 3157 19193 3191 19227
rect 3191 19193 3200 19227
rect 3148 19184 3200 19193
rect 2688 19116 2740 19168
rect 3056 19116 3108 19168
rect 3792 19116 3844 19168
rect 4528 19159 4580 19168
rect 4528 19125 4537 19159
rect 4537 19125 4571 19159
rect 4571 19125 4580 19159
rect 4528 19116 4580 19125
rect 6552 19116 6604 19168
rect 6828 19184 6880 19236
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 8852 19252 8904 19304
rect 11704 19388 11756 19440
rect 12624 19388 12676 19440
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 10508 19252 10560 19304
rect 11520 19252 11572 19304
rect 11796 19184 11848 19236
rect 11980 19252 12032 19304
rect 13360 19456 13412 19508
rect 12900 19388 12952 19440
rect 13544 19388 13596 19440
rect 14740 19388 14792 19440
rect 15384 19456 15436 19508
rect 15108 19388 15160 19440
rect 15936 19388 15988 19440
rect 15844 19320 15896 19372
rect 8116 19116 8168 19168
rect 8760 19116 8812 19168
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 10876 19116 10928 19125
rect 11152 19116 11204 19168
rect 12072 19184 12124 19236
rect 12164 19116 12216 19168
rect 13084 19184 13136 19236
rect 14280 19184 14332 19236
rect 14924 19184 14976 19236
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 16120 19252 16172 19304
rect 17960 19456 18012 19508
rect 18604 19456 18656 19508
rect 21180 19456 21232 19508
rect 17132 19388 17184 19440
rect 17316 19388 17368 19440
rect 19248 19388 19300 19440
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 17868 19320 17920 19372
rect 18512 19320 18564 19372
rect 16580 19184 16632 19236
rect 17592 19184 17644 19236
rect 18604 19184 18656 19236
rect 15936 19116 15988 19168
rect 16396 19116 16448 19168
rect 17316 19116 17368 19168
rect 17500 19116 17552 19168
rect 17776 19116 17828 19168
rect 17868 19116 17920 19168
rect 20352 19388 20404 19440
rect 22008 19456 22060 19508
rect 20260 19252 20312 19304
rect 21272 19295 21324 19304
rect 21272 19261 21290 19295
rect 21290 19261 21324 19295
rect 21272 19252 21324 19261
rect 22284 19252 22336 19304
rect 22376 19252 22428 19304
rect 22744 19252 22796 19304
rect 23296 19295 23348 19304
rect 23296 19261 23305 19295
rect 23305 19261 23339 19295
rect 23339 19261 23348 19295
rect 23296 19252 23348 19261
rect 23480 19320 23532 19372
rect 23848 19320 23900 19372
rect 23756 19295 23808 19304
rect 23756 19261 23765 19295
rect 23765 19261 23799 19295
rect 23799 19261 23808 19295
rect 23756 19252 23808 19261
rect 24400 19295 24452 19304
rect 24400 19261 24409 19295
rect 24409 19261 24443 19295
rect 24443 19261 24452 19295
rect 24400 19252 24452 19261
rect 25596 19252 25648 19304
rect 30748 19456 30800 19508
rect 27344 19363 27396 19372
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 28172 19388 28224 19440
rect 27252 19295 27304 19304
rect 27252 19261 27261 19295
rect 27261 19261 27295 19295
rect 27295 19261 27304 19295
rect 27252 19252 27304 19261
rect 28908 19320 28960 19372
rect 30472 19320 30524 19372
rect 22560 19159 22612 19168
rect 22560 19125 22569 19159
rect 22569 19125 22603 19159
rect 22603 19125 22612 19159
rect 22560 19116 22612 19125
rect 22928 19116 22980 19168
rect 25504 19116 25556 19168
rect 27528 19184 27580 19236
rect 27712 19252 27764 19304
rect 28356 19252 28408 19304
rect 28724 19252 28776 19304
rect 29000 19252 29052 19304
rect 30656 19184 30708 19236
rect 26332 19116 26384 19168
rect 27804 19159 27856 19168
rect 27804 19125 27813 19159
rect 27813 19125 27847 19159
rect 27847 19125 27856 19159
rect 27804 19116 27856 19125
rect 28816 19116 28868 19168
rect 29736 19116 29788 19168
rect 30380 19116 30432 19168
rect 11253 19014 11305 19066
rect 11317 19014 11369 19066
rect 11381 19014 11433 19066
rect 11445 19014 11497 19066
rect 11509 19014 11561 19066
rect 21557 19014 21609 19066
rect 21621 19014 21673 19066
rect 21685 19014 21737 19066
rect 21749 19014 21801 19066
rect 21813 19014 21865 19066
rect 1400 18776 1452 18828
rect 2228 18912 2280 18964
rect 3056 18912 3108 18964
rect 3240 18912 3292 18964
rect 4436 18955 4488 18964
rect 4436 18921 4445 18955
rect 4445 18921 4479 18955
rect 4479 18921 4488 18955
rect 6828 18955 6880 18964
rect 4436 18912 4488 18921
rect 1676 18819 1728 18828
rect 1676 18785 1685 18819
rect 1685 18785 1719 18819
rect 1719 18785 1728 18819
rect 1676 18776 1728 18785
rect 2136 18844 2188 18896
rect 2320 18844 2372 18896
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 9128 18912 9180 18964
rect 10600 18912 10652 18964
rect 13084 18912 13136 18964
rect 13360 18912 13412 18964
rect 14096 18912 14148 18964
rect 15292 18912 15344 18964
rect 15476 18912 15528 18964
rect 16672 18912 16724 18964
rect 17684 18912 17736 18964
rect 18328 18912 18380 18964
rect 19248 18912 19300 18964
rect 2044 18819 2096 18828
rect 2044 18785 2053 18819
rect 2053 18785 2087 18819
rect 2087 18785 2096 18819
rect 2044 18776 2096 18785
rect 2688 18819 2740 18828
rect 2688 18785 2697 18819
rect 2697 18785 2731 18819
rect 2731 18785 2740 18819
rect 2688 18776 2740 18785
rect 3240 18776 3292 18828
rect 3608 18776 3660 18828
rect 3884 18819 3936 18828
rect 3884 18785 3893 18819
rect 3893 18785 3927 18819
rect 3927 18785 3936 18819
rect 3884 18776 3936 18785
rect 4252 18776 4304 18828
rect 4620 18776 4672 18828
rect 5264 18819 5316 18828
rect 5264 18785 5273 18819
rect 5273 18785 5307 18819
rect 5307 18785 5316 18819
rect 5264 18776 5316 18785
rect 8116 18844 8168 18896
rect 10876 18844 10928 18896
rect 11796 18844 11848 18896
rect 12348 18844 12400 18896
rect 12900 18844 12952 18896
rect 19340 18844 19392 18896
rect 19800 18912 19852 18964
rect 20904 18955 20956 18964
rect 20904 18921 20913 18955
rect 20913 18921 20947 18955
rect 20947 18921 20956 18955
rect 20904 18912 20956 18921
rect 21916 18955 21968 18964
rect 21916 18921 21925 18955
rect 21925 18921 21959 18955
rect 21959 18921 21968 18955
rect 21916 18912 21968 18921
rect 22468 18912 22520 18964
rect 23572 18912 23624 18964
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 1952 18708 2004 18760
rect 2320 18708 2372 18760
rect 2780 18708 2832 18760
rect 4804 18708 4856 18760
rect 5816 18776 5868 18828
rect 7012 18776 7064 18828
rect 7656 18776 7708 18828
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 7472 18708 7524 18760
rect 7840 18776 7892 18828
rect 8024 18776 8076 18828
rect 8208 18776 8260 18828
rect 10968 18776 11020 18828
rect 11244 18776 11296 18828
rect 8944 18708 8996 18760
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 10876 18708 10928 18760
rect 11152 18708 11204 18760
rect 3332 18640 3384 18692
rect 7840 18640 7892 18692
rect 10968 18640 11020 18692
rect 13452 18776 13504 18828
rect 14372 18776 14424 18828
rect 14556 18819 14608 18828
rect 14556 18785 14590 18819
rect 14590 18785 14608 18819
rect 14556 18776 14608 18785
rect 14924 18776 14976 18828
rect 15936 18776 15988 18828
rect 16304 18776 16356 18828
rect 16856 18819 16908 18828
rect 12348 18708 12400 18760
rect 1492 18572 1544 18624
rect 1676 18572 1728 18624
rect 2228 18615 2280 18624
rect 2228 18581 2237 18615
rect 2237 18581 2271 18615
rect 2271 18581 2280 18615
rect 2228 18572 2280 18581
rect 5172 18572 5224 18624
rect 6460 18572 6512 18624
rect 8116 18572 8168 18624
rect 8760 18572 8812 18624
rect 10508 18572 10560 18624
rect 15292 18708 15344 18760
rect 15844 18708 15896 18760
rect 16856 18785 16865 18819
rect 16865 18785 16899 18819
rect 16899 18785 16908 18819
rect 16856 18776 16908 18785
rect 17224 18776 17276 18828
rect 17316 18776 17368 18828
rect 18144 18776 18196 18828
rect 18604 18819 18656 18828
rect 18604 18785 18638 18819
rect 18638 18785 18656 18819
rect 18604 18776 18656 18785
rect 18880 18776 18932 18828
rect 17132 18708 17184 18760
rect 16580 18640 16632 18692
rect 16948 18640 17000 18692
rect 17224 18640 17276 18692
rect 18328 18640 18380 18692
rect 19432 18776 19484 18828
rect 20168 18819 20220 18828
rect 20168 18785 20177 18819
rect 20177 18785 20211 18819
rect 20211 18785 20220 18819
rect 20168 18776 20220 18785
rect 21456 18844 21508 18896
rect 24584 18912 24636 18964
rect 20352 18819 20404 18828
rect 20352 18785 20361 18819
rect 20361 18785 20395 18819
rect 20395 18785 20404 18819
rect 20352 18776 20404 18785
rect 22008 18819 22060 18828
rect 22008 18785 22017 18819
rect 22017 18785 22051 18819
rect 22051 18785 22060 18819
rect 22008 18776 22060 18785
rect 22744 18819 22796 18828
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 23480 18776 23532 18828
rect 27804 18912 27856 18964
rect 27160 18844 27212 18896
rect 28080 18844 28132 18896
rect 28816 18887 28868 18896
rect 28816 18853 28834 18887
rect 28834 18853 28868 18887
rect 30656 18912 30708 18964
rect 28816 18844 28868 18853
rect 19616 18708 19668 18760
rect 20812 18708 20864 18760
rect 20904 18708 20956 18760
rect 24584 18751 24636 18760
rect 23664 18640 23716 18692
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 27988 18776 28040 18828
rect 29644 18776 29696 18828
rect 26424 18708 26476 18760
rect 26332 18640 26384 18692
rect 16120 18572 16172 18624
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 17316 18572 17368 18624
rect 17408 18572 17460 18624
rect 17592 18572 17644 18624
rect 19340 18572 19392 18624
rect 19800 18572 19852 18624
rect 19892 18572 19944 18624
rect 23112 18572 23164 18624
rect 25320 18572 25372 18624
rect 27160 18615 27212 18624
rect 27160 18581 27169 18615
rect 27169 18581 27203 18615
rect 27203 18581 27212 18615
rect 27160 18572 27212 18581
rect 28724 18572 28776 18624
rect 6102 18470 6154 18522
rect 6166 18470 6218 18522
rect 6230 18470 6282 18522
rect 6294 18470 6346 18522
rect 6358 18470 6410 18522
rect 16405 18470 16457 18522
rect 16469 18470 16521 18522
rect 16533 18470 16585 18522
rect 16597 18470 16649 18522
rect 16661 18470 16713 18522
rect 26709 18470 26761 18522
rect 26773 18470 26825 18522
rect 26837 18470 26889 18522
rect 26901 18470 26953 18522
rect 26965 18470 27017 18522
rect 4068 18368 4120 18420
rect 5632 18368 5684 18420
rect 8116 18411 8168 18420
rect 5540 18300 5592 18352
rect 8116 18377 8125 18411
rect 8125 18377 8159 18411
rect 8159 18377 8168 18411
rect 8116 18368 8168 18377
rect 8852 18368 8904 18420
rect 9404 18368 9456 18420
rect 11060 18368 11112 18420
rect 12348 18368 12400 18420
rect 14004 18368 14056 18420
rect 15936 18411 15988 18420
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 2228 18164 2280 18216
rect 2688 18164 2740 18216
rect 4528 18164 4580 18216
rect 5632 18232 5684 18284
rect 6736 18232 6788 18284
rect 9128 18300 9180 18352
rect 9496 18300 9548 18352
rect 10232 18300 10284 18352
rect 12808 18300 12860 18352
rect 13268 18300 13320 18352
rect 15568 18343 15620 18352
rect 15568 18309 15577 18343
rect 15577 18309 15611 18343
rect 15611 18309 15620 18343
rect 15568 18300 15620 18309
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16212 18368 16264 18420
rect 17316 18368 17368 18420
rect 18328 18368 18380 18420
rect 19248 18368 19300 18420
rect 9864 18275 9916 18284
rect 6460 18164 6512 18216
rect 7012 18207 7064 18216
rect 7012 18173 7021 18207
rect 7021 18173 7055 18207
rect 7055 18173 7064 18207
rect 7012 18164 7064 18173
rect 7472 18207 7524 18216
rect 7472 18173 7481 18207
rect 7481 18173 7515 18207
rect 7515 18173 7524 18207
rect 7472 18164 7524 18173
rect 7932 18164 7984 18216
rect 8484 18164 8536 18216
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 10416 18164 10468 18216
rect 11704 18164 11756 18216
rect 14648 18232 14700 18284
rect 14924 18232 14976 18284
rect 15476 18232 15528 18284
rect 17224 18300 17276 18352
rect 20444 18368 20496 18420
rect 23664 18368 23716 18420
rect 27068 18368 27120 18420
rect 14004 18164 14056 18216
rect 14096 18164 14148 18216
rect 8300 18096 8352 18148
rect 9496 18096 9548 18148
rect 14188 18096 14240 18148
rect 14924 18096 14976 18148
rect 16304 18096 16356 18148
rect 1492 18028 1544 18080
rect 2044 18028 2096 18080
rect 2780 18028 2832 18080
rect 4068 18028 4120 18080
rect 4252 18028 4304 18080
rect 4712 18028 4764 18080
rect 5724 18028 5776 18080
rect 6000 18071 6052 18080
rect 6000 18037 6009 18071
rect 6009 18037 6043 18071
rect 6043 18037 6052 18071
rect 6000 18028 6052 18037
rect 8208 18028 8260 18080
rect 10048 18028 10100 18080
rect 11612 18028 11664 18080
rect 11796 18028 11848 18080
rect 12808 18028 12860 18080
rect 14556 18028 14608 18080
rect 15752 18028 15804 18080
rect 16212 18028 16264 18080
rect 16672 18164 16724 18216
rect 16764 18164 16816 18216
rect 17224 18164 17276 18216
rect 17684 18164 17736 18216
rect 17776 18164 17828 18216
rect 18328 18207 18380 18216
rect 18328 18173 18337 18207
rect 18337 18173 18371 18207
rect 18371 18173 18380 18207
rect 18328 18164 18380 18173
rect 18696 18232 18748 18284
rect 19892 18300 19944 18352
rect 20536 18300 20588 18352
rect 28908 18368 28960 18420
rect 20812 18232 20864 18284
rect 19340 18164 19392 18216
rect 19800 18207 19852 18216
rect 18052 18096 18104 18148
rect 18512 18096 18564 18148
rect 18880 18096 18932 18148
rect 19156 18096 19208 18148
rect 19800 18173 19809 18207
rect 19809 18173 19843 18207
rect 19843 18173 19852 18207
rect 19800 18164 19852 18173
rect 19616 18096 19668 18148
rect 22652 18164 22704 18216
rect 23388 18164 23440 18216
rect 17592 18028 17644 18080
rect 19892 18028 19944 18080
rect 20536 18071 20588 18080
rect 20536 18037 20545 18071
rect 20545 18037 20579 18071
rect 20579 18037 20588 18071
rect 20536 18028 20588 18037
rect 21088 18028 21140 18080
rect 22008 18096 22060 18148
rect 23756 18139 23808 18148
rect 23756 18105 23765 18139
rect 23765 18105 23799 18139
rect 23799 18105 23808 18139
rect 23756 18096 23808 18105
rect 22192 18028 22244 18080
rect 22836 18028 22888 18080
rect 23664 18071 23716 18080
rect 23664 18037 23673 18071
rect 23673 18037 23707 18071
rect 23707 18037 23716 18071
rect 23664 18028 23716 18037
rect 25228 18028 25280 18080
rect 26240 18028 26292 18080
rect 29000 18164 29052 18216
rect 29736 18164 29788 18216
rect 27804 18139 27856 18148
rect 27804 18105 27838 18139
rect 27838 18105 27856 18139
rect 27804 18096 27856 18105
rect 30288 18096 30340 18148
rect 27252 18028 27304 18080
rect 30472 18028 30524 18080
rect 31300 18071 31352 18080
rect 31300 18037 31309 18071
rect 31309 18037 31343 18071
rect 31343 18037 31352 18071
rect 31300 18028 31352 18037
rect 11253 17926 11305 17978
rect 11317 17926 11369 17978
rect 11381 17926 11433 17978
rect 11445 17926 11497 17978
rect 11509 17926 11561 17978
rect 21557 17926 21609 17978
rect 21621 17926 21673 17978
rect 21685 17926 21737 17978
rect 21749 17926 21801 17978
rect 21813 17926 21865 17978
rect 1952 17824 2004 17876
rect 3884 17824 3936 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 1492 17688 1544 17740
rect 1768 17756 1820 17808
rect 8208 17867 8260 17876
rect 8208 17833 8233 17867
rect 8233 17833 8260 17867
rect 8392 17867 8444 17876
rect 8208 17824 8260 17833
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 7932 17756 7984 17808
rect 2688 17688 2740 17740
rect 5632 17688 5684 17740
rect 6920 17731 6972 17740
rect 6920 17697 6929 17731
rect 6929 17697 6963 17731
rect 6963 17697 6972 17731
rect 6920 17688 6972 17697
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 5540 17620 5592 17672
rect 10600 17824 10652 17876
rect 11612 17824 11664 17876
rect 12992 17824 13044 17876
rect 16948 17824 17000 17876
rect 8668 17756 8720 17808
rect 9864 17756 9916 17808
rect 10508 17756 10560 17808
rect 9956 17688 10008 17740
rect 10416 17688 10468 17740
rect 10876 17731 10928 17740
rect 10876 17697 10885 17731
rect 10885 17697 10919 17731
rect 10919 17697 10928 17731
rect 15752 17756 15804 17808
rect 16120 17756 16172 17808
rect 10876 17688 10928 17697
rect 12348 17731 12400 17740
rect 12348 17697 12357 17731
rect 12357 17697 12391 17731
rect 12391 17697 12400 17731
rect 12348 17688 12400 17697
rect 13084 17688 13136 17740
rect 14188 17731 14240 17740
rect 14188 17697 14197 17731
rect 14197 17697 14231 17731
rect 14231 17697 14240 17731
rect 14188 17688 14240 17697
rect 15108 17688 15160 17740
rect 17132 17756 17184 17808
rect 18604 17824 18656 17876
rect 18972 17824 19024 17876
rect 19524 17824 19576 17876
rect 17776 17799 17828 17808
rect 17776 17765 17785 17799
rect 17785 17765 17819 17799
rect 17819 17765 17828 17799
rect 17776 17756 17828 17765
rect 18236 17799 18288 17808
rect 18236 17765 18245 17799
rect 18245 17765 18279 17799
rect 18279 17765 18288 17799
rect 18236 17756 18288 17765
rect 20076 17824 20128 17876
rect 20628 17824 20680 17876
rect 20168 17756 20220 17808
rect 23020 17824 23072 17876
rect 23388 17824 23440 17876
rect 24216 17824 24268 17876
rect 27804 17824 27856 17876
rect 17592 17731 17644 17740
rect 9404 17620 9456 17672
rect 10048 17620 10100 17672
rect 11888 17620 11940 17672
rect 13544 17620 13596 17672
rect 15476 17620 15528 17672
rect 3884 17552 3936 17604
rect 6460 17552 6512 17604
rect 6920 17552 6972 17604
rect 7196 17552 7248 17604
rect 10416 17552 10468 17604
rect 10876 17552 10928 17604
rect 2872 17484 2924 17536
rect 5264 17527 5316 17536
rect 5264 17493 5273 17527
rect 5273 17493 5307 17527
rect 5307 17493 5316 17527
rect 5264 17484 5316 17493
rect 5908 17484 5960 17536
rect 7840 17484 7892 17536
rect 9588 17484 9640 17536
rect 10600 17484 10652 17536
rect 16856 17552 16908 17604
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 20352 17688 20404 17740
rect 25320 17799 25372 17808
rect 25320 17765 25354 17799
rect 25354 17765 25372 17799
rect 25320 17756 25372 17765
rect 25872 17756 25924 17808
rect 18052 17620 18104 17672
rect 20536 17620 20588 17672
rect 19800 17552 19852 17604
rect 20260 17552 20312 17604
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 20812 17620 20864 17629
rect 22284 17731 22336 17740
rect 22284 17697 22293 17731
rect 22293 17697 22327 17731
rect 22327 17697 22336 17731
rect 22284 17688 22336 17697
rect 22560 17731 22612 17740
rect 22560 17697 22594 17731
rect 22594 17697 22612 17731
rect 24216 17731 24268 17740
rect 22560 17688 22612 17697
rect 24216 17697 24225 17731
rect 24225 17697 24259 17731
rect 24259 17697 24268 17731
rect 24216 17688 24268 17697
rect 26516 17688 26568 17740
rect 21364 17620 21416 17672
rect 14464 17484 14516 17536
rect 18236 17484 18288 17536
rect 18512 17484 18564 17536
rect 18604 17484 18656 17536
rect 20996 17484 21048 17536
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 22100 17484 22152 17536
rect 23940 17484 23992 17536
rect 27252 17756 27304 17808
rect 27620 17756 27672 17808
rect 30840 17824 30892 17876
rect 30932 17824 30984 17876
rect 27252 17663 27304 17672
rect 27252 17629 27261 17663
rect 27261 17629 27295 17663
rect 27295 17629 27304 17663
rect 27252 17620 27304 17629
rect 25228 17484 25280 17536
rect 26424 17527 26476 17536
rect 26424 17493 26433 17527
rect 26433 17493 26467 17527
rect 26467 17493 26476 17527
rect 26424 17484 26476 17493
rect 28448 17527 28500 17536
rect 28448 17493 28457 17527
rect 28457 17493 28491 17527
rect 28491 17493 28500 17527
rect 28448 17484 28500 17493
rect 28632 17527 28684 17536
rect 28632 17493 28641 17527
rect 28641 17493 28675 17527
rect 28675 17493 28684 17527
rect 28632 17484 28684 17493
rect 29920 17756 29972 17808
rect 30196 17731 30248 17740
rect 30196 17697 30230 17731
rect 30230 17697 30248 17731
rect 30196 17688 30248 17697
rect 29736 17620 29788 17672
rect 30656 17484 30708 17536
rect 6102 17382 6154 17434
rect 6166 17382 6218 17434
rect 6230 17382 6282 17434
rect 6294 17382 6346 17434
rect 6358 17382 6410 17434
rect 16405 17382 16457 17434
rect 16469 17382 16521 17434
rect 16533 17382 16585 17434
rect 16597 17382 16649 17434
rect 16661 17382 16713 17434
rect 26709 17382 26761 17434
rect 26773 17382 26825 17434
rect 26837 17382 26889 17434
rect 26901 17382 26953 17434
rect 26965 17382 27017 17434
rect 1768 17280 1820 17332
rect 8484 17280 8536 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 9956 17280 10008 17332
rect 4068 17212 4120 17264
rect 5264 17212 5316 17264
rect 3608 17144 3660 17196
rect 3976 17144 4028 17196
rect 5540 17144 5592 17196
rect 6000 17212 6052 17264
rect 9864 17144 9916 17196
rect 10968 17212 11020 17264
rect 3056 17076 3108 17128
rect 4620 17119 4672 17128
rect 4620 17085 4629 17119
rect 4629 17085 4663 17119
rect 4663 17085 4672 17119
rect 4620 17076 4672 17085
rect 4804 17076 4856 17128
rect 5356 17076 5408 17128
rect 5724 17119 5776 17128
rect 5724 17085 5733 17119
rect 5733 17085 5767 17119
rect 5767 17085 5776 17119
rect 5724 17076 5776 17085
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 7472 17076 7524 17128
rect 9956 17119 10008 17128
rect 9956 17085 9965 17119
rect 9965 17085 9999 17119
rect 9999 17085 10008 17119
rect 9956 17076 10008 17085
rect 3148 17008 3200 17060
rect 6000 17008 6052 17060
rect 6460 17008 6512 17060
rect 10508 17085 10517 17106
rect 10517 17085 10551 17106
rect 10551 17085 10560 17106
rect 10508 17054 10560 17085
rect 2780 16940 2832 16992
rect 3424 16940 3476 16992
rect 3884 16940 3936 16992
rect 4160 16983 4212 16992
rect 4160 16949 4169 16983
rect 4169 16949 4203 16983
rect 4203 16949 4212 16983
rect 4160 16940 4212 16949
rect 5264 16940 5316 16992
rect 10876 17144 10928 17196
rect 11060 17076 11112 17128
rect 11612 17280 11664 17332
rect 12532 17280 12584 17332
rect 13084 17323 13136 17332
rect 11888 17212 11940 17264
rect 11612 17144 11664 17196
rect 11980 17144 12032 17196
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 12072 17076 12124 17128
rect 12348 17119 12400 17128
rect 12348 17085 12357 17119
rect 12357 17085 12391 17119
rect 12391 17085 12400 17119
rect 12348 17076 12400 17085
rect 12440 17076 12492 17128
rect 13084 17289 13093 17323
rect 13093 17289 13127 17323
rect 13127 17289 13136 17323
rect 13084 17280 13136 17289
rect 15292 17280 15344 17332
rect 16764 17280 16816 17332
rect 17224 17280 17276 17332
rect 17500 17280 17552 17332
rect 17592 17280 17644 17332
rect 19248 17280 19300 17332
rect 14280 17255 14332 17264
rect 14280 17221 14289 17255
rect 14289 17221 14323 17255
rect 14323 17221 14332 17255
rect 14280 17212 14332 17221
rect 12808 17144 12860 17196
rect 15476 17144 15528 17196
rect 16396 17144 16448 17196
rect 17868 17144 17920 17196
rect 18328 17212 18380 17264
rect 22468 17280 22520 17332
rect 24216 17280 24268 17332
rect 30104 17280 30156 17332
rect 30288 17323 30340 17332
rect 30288 17289 30297 17323
rect 30297 17289 30331 17323
rect 30331 17289 30340 17323
rect 30288 17280 30340 17289
rect 30656 17280 30708 17332
rect 20536 17144 20588 17196
rect 12992 17076 13044 17128
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 11980 16940 12032 16992
rect 14372 17076 14424 17128
rect 14464 17008 14516 17060
rect 14740 17008 14792 17060
rect 15476 17008 15528 17060
rect 15844 17008 15896 17060
rect 16304 17076 16356 17128
rect 17132 17119 17184 17128
rect 17132 17085 17141 17119
rect 17141 17085 17175 17119
rect 17175 17085 17184 17119
rect 17132 17076 17184 17085
rect 15752 16940 15804 16992
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 17132 16940 17184 16992
rect 17592 17076 17644 17128
rect 17960 17076 18012 17128
rect 18788 17076 18840 17128
rect 19616 17119 19668 17128
rect 18512 17051 18564 17060
rect 18512 17017 18521 17051
rect 18521 17017 18555 17051
rect 18555 17017 18564 17051
rect 18512 17008 18564 17017
rect 19064 17008 19116 17060
rect 19616 17085 19625 17119
rect 19625 17085 19659 17119
rect 19659 17085 19668 17119
rect 19616 17076 19668 17085
rect 20444 17076 20496 17128
rect 20812 17119 20864 17128
rect 20812 17085 20821 17119
rect 20821 17085 20855 17119
rect 20855 17085 20864 17119
rect 20812 17076 20864 17085
rect 23848 17144 23900 17196
rect 23480 17119 23532 17128
rect 23480 17085 23489 17119
rect 23489 17085 23523 17119
rect 23523 17085 23532 17119
rect 23480 17076 23532 17085
rect 28632 17212 28684 17264
rect 19524 17008 19576 17060
rect 17776 16940 17828 16992
rect 18880 16940 18932 16992
rect 21456 17008 21508 17060
rect 23204 17008 23256 17060
rect 25228 17076 25280 17128
rect 26148 17076 26200 17128
rect 27160 17144 27212 17196
rect 29276 17144 29328 17196
rect 26516 17119 26568 17128
rect 26516 17085 26525 17119
rect 26525 17085 26559 17119
rect 26559 17085 26568 17119
rect 26516 17076 26568 17085
rect 29644 17144 29696 17196
rect 30288 17144 30340 17196
rect 30932 17144 30984 17196
rect 29828 17119 29880 17128
rect 29828 17085 29837 17119
rect 29837 17085 29871 17119
rect 29871 17085 29880 17119
rect 29828 17076 29880 17085
rect 30012 17076 30064 17128
rect 30104 17119 30156 17128
rect 30104 17085 30113 17119
rect 30113 17085 30147 17119
rect 30147 17085 30156 17119
rect 30104 17076 30156 17085
rect 30472 17076 30524 17128
rect 30656 17076 30708 17128
rect 21916 16940 21968 16992
rect 22192 16983 22244 16992
rect 22192 16949 22201 16983
rect 22201 16949 22235 16983
rect 22235 16949 22244 16983
rect 22192 16940 22244 16949
rect 23112 16940 23164 16992
rect 26976 16940 27028 16992
rect 28816 16940 28868 16992
rect 11253 16838 11305 16890
rect 11317 16838 11369 16890
rect 11381 16838 11433 16890
rect 11445 16838 11497 16890
rect 11509 16838 11561 16890
rect 21557 16838 21609 16890
rect 21621 16838 21673 16890
rect 21685 16838 21737 16890
rect 21749 16838 21801 16890
rect 21813 16838 21865 16890
rect 1216 16736 1268 16788
rect 2596 16736 2648 16788
rect 3424 16736 3476 16788
rect 3700 16736 3752 16788
rect 4160 16736 4212 16788
rect 1400 16600 1452 16652
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 2136 16643 2188 16652
rect 2136 16609 2145 16643
rect 2145 16609 2179 16643
rect 2179 16609 2188 16643
rect 2136 16600 2188 16609
rect 2228 16643 2280 16652
rect 2228 16609 2237 16643
rect 2237 16609 2271 16643
rect 2271 16609 2280 16643
rect 2228 16600 2280 16609
rect 2044 16532 2096 16584
rect 3148 16643 3200 16652
rect 3148 16609 3157 16643
rect 3157 16609 3191 16643
rect 3191 16609 3200 16643
rect 5080 16668 5132 16720
rect 6736 16736 6788 16788
rect 7380 16736 7432 16788
rect 9220 16736 9272 16788
rect 3148 16600 3200 16609
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 7012 16600 7064 16652
rect 8944 16643 8996 16652
rect 8944 16609 8953 16643
rect 8953 16609 8987 16643
rect 8987 16609 8996 16643
rect 8944 16600 8996 16609
rect 9404 16643 9456 16652
rect 9404 16609 9413 16643
rect 9413 16609 9447 16643
rect 9447 16609 9456 16643
rect 9404 16600 9456 16609
rect 4252 16532 4304 16584
rect 8852 16532 8904 16584
rect 9220 16532 9272 16584
rect 9864 16736 9916 16788
rect 10600 16736 10652 16788
rect 11980 16736 12032 16788
rect 10232 16668 10284 16720
rect 11060 16668 11112 16720
rect 12348 16736 12400 16788
rect 12440 16736 12492 16788
rect 13544 16736 13596 16788
rect 14372 16736 14424 16788
rect 13912 16668 13964 16720
rect 14556 16668 14608 16720
rect 15568 16736 15620 16788
rect 15844 16736 15896 16788
rect 17408 16736 17460 16788
rect 17592 16736 17644 16788
rect 17868 16736 17920 16788
rect 20260 16736 20312 16788
rect 22468 16736 22520 16788
rect 22560 16736 22612 16788
rect 23756 16779 23808 16788
rect 23756 16745 23765 16779
rect 23765 16745 23799 16779
rect 23799 16745 23808 16779
rect 23756 16736 23808 16745
rect 2596 16464 2648 16516
rect 6552 16464 6604 16516
rect 10416 16532 10468 16584
rect 11704 16600 11756 16652
rect 11980 16600 12032 16652
rect 12164 16600 12216 16652
rect 12900 16600 12952 16652
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 14004 16600 14056 16652
rect 14924 16600 14976 16652
rect 15200 16600 15252 16652
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 18144 16668 18196 16720
rect 16948 16643 17000 16652
rect 16948 16609 16982 16643
rect 16982 16609 17000 16643
rect 16948 16600 17000 16609
rect 17408 16600 17460 16652
rect 17960 16600 18012 16652
rect 18604 16600 18656 16652
rect 18880 16643 18932 16652
rect 18880 16609 18889 16643
rect 18889 16609 18923 16643
rect 18923 16609 18932 16643
rect 18880 16600 18932 16609
rect 19064 16643 19116 16652
rect 19064 16609 19073 16643
rect 19073 16609 19107 16643
rect 19107 16609 19116 16643
rect 19064 16600 19116 16609
rect 20812 16668 20864 16720
rect 26148 16736 26200 16788
rect 26976 16779 27028 16788
rect 26976 16745 26985 16779
rect 26985 16745 27019 16779
rect 27019 16745 27028 16779
rect 26976 16736 27028 16745
rect 28908 16736 28960 16788
rect 19892 16600 19944 16652
rect 20536 16600 20588 16652
rect 22008 16643 22060 16652
rect 22008 16609 22017 16643
rect 22017 16609 22051 16643
rect 22051 16609 22060 16643
rect 22008 16600 22060 16609
rect 22192 16643 22244 16652
rect 22192 16609 22201 16643
rect 22201 16609 22235 16643
rect 22235 16609 22244 16643
rect 22192 16600 22244 16609
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 23112 16643 23164 16652
rect 23112 16609 23121 16643
rect 23121 16609 23155 16643
rect 23155 16609 23164 16643
rect 23112 16600 23164 16609
rect 23572 16600 23624 16652
rect 23848 16600 23900 16652
rect 24676 16600 24728 16652
rect 25872 16643 25924 16652
rect 25872 16609 25881 16643
rect 25881 16609 25915 16643
rect 25915 16609 25924 16643
rect 25872 16600 25924 16609
rect 26148 16600 26200 16652
rect 28448 16600 28500 16652
rect 28908 16643 28960 16652
rect 28908 16609 28917 16643
rect 28917 16609 28951 16643
rect 28951 16609 28960 16643
rect 28908 16600 28960 16609
rect 29276 16668 29328 16720
rect 29460 16668 29512 16720
rect 30196 16736 30248 16788
rect 30564 16736 30616 16788
rect 30840 16736 30892 16788
rect 31024 16736 31076 16788
rect 30472 16668 30524 16720
rect 11796 16575 11848 16584
rect 9956 16464 10008 16516
rect 10692 16464 10744 16516
rect 2504 16396 2556 16448
rect 3700 16396 3752 16448
rect 4068 16396 4120 16448
rect 8852 16439 8904 16448
rect 8852 16405 8861 16439
rect 8861 16405 8895 16439
rect 8895 16405 8904 16439
rect 8852 16396 8904 16405
rect 10508 16439 10560 16448
rect 10508 16405 10517 16439
rect 10517 16405 10551 16439
rect 10551 16405 10560 16439
rect 10508 16396 10560 16405
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 12808 16532 12860 16584
rect 13084 16532 13136 16584
rect 14188 16532 14240 16584
rect 14372 16532 14424 16584
rect 15292 16532 15344 16584
rect 15844 16532 15896 16584
rect 18144 16532 18196 16584
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 12808 16396 12860 16448
rect 13268 16396 13320 16448
rect 16304 16396 16356 16448
rect 18236 16464 18288 16516
rect 19156 16464 19208 16516
rect 23204 16532 23256 16584
rect 24308 16575 24360 16584
rect 24308 16541 24317 16575
rect 24317 16541 24351 16575
rect 24351 16541 24360 16575
rect 24308 16532 24360 16541
rect 27252 16532 27304 16584
rect 28816 16532 28868 16584
rect 22928 16507 22980 16516
rect 22928 16473 22937 16507
rect 22937 16473 22971 16507
rect 22971 16473 22980 16507
rect 22928 16464 22980 16473
rect 24492 16464 24544 16516
rect 28080 16464 28132 16516
rect 22836 16396 22888 16448
rect 27344 16396 27396 16448
rect 29644 16600 29696 16652
rect 30012 16600 30064 16652
rect 30288 16600 30340 16652
rect 31392 16600 31444 16652
rect 29092 16575 29144 16584
rect 29092 16541 29101 16575
rect 29101 16541 29135 16575
rect 29135 16541 29144 16575
rect 29092 16532 29144 16541
rect 29276 16532 29328 16584
rect 29828 16575 29880 16584
rect 29828 16541 29837 16575
rect 29837 16541 29871 16575
rect 29871 16541 29880 16575
rect 29828 16532 29880 16541
rect 29184 16464 29236 16516
rect 6102 16294 6154 16346
rect 6166 16294 6218 16346
rect 6230 16294 6282 16346
rect 6294 16294 6346 16346
rect 6358 16294 6410 16346
rect 16405 16294 16457 16346
rect 16469 16294 16521 16346
rect 16533 16294 16585 16346
rect 16597 16294 16649 16346
rect 16661 16294 16713 16346
rect 26709 16294 26761 16346
rect 26773 16294 26825 16346
rect 26837 16294 26889 16346
rect 26901 16294 26953 16346
rect 26965 16294 27017 16346
rect 2044 16192 2096 16244
rect 4252 16192 4304 16244
rect 4896 16192 4948 16244
rect 5172 16192 5224 16244
rect 7012 16192 7064 16244
rect 8300 16192 8352 16244
rect 8760 16192 8812 16244
rect 1952 16056 2004 16108
rect 2596 16056 2648 16108
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 5448 16056 5500 16108
rect 4252 16031 4304 16040
rect 4252 15997 4261 16031
rect 4261 15997 4295 16031
rect 4295 15997 4304 16031
rect 4252 15988 4304 15997
rect 4620 15988 4672 16040
rect 5264 15988 5316 16040
rect 3148 15963 3200 15972
rect 3148 15929 3157 15963
rect 3157 15929 3191 15963
rect 3191 15929 3200 15963
rect 3148 15920 3200 15929
rect 4988 15920 5040 15972
rect 1308 15852 1360 15904
rect 4068 15852 4120 15904
rect 5540 15852 5592 15904
rect 9312 16124 9364 16176
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 7196 16056 7248 16108
rect 8208 16056 8260 16108
rect 6460 16031 6512 16040
rect 6460 15997 6469 16031
rect 6469 15997 6503 16031
rect 6503 15997 6512 16031
rect 6736 16031 6788 16040
rect 6460 15988 6512 15997
rect 6736 15997 6745 16031
rect 6745 15997 6779 16031
rect 6779 15997 6788 16031
rect 6736 15988 6788 15997
rect 7656 16031 7708 16040
rect 7656 15997 7665 16031
rect 7665 15997 7699 16031
rect 7699 15997 7708 16031
rect 7656 15988 7708 15997
rect 8392 16031 8444 16040
rect 6828 15920 6880 15972
rect 7288 15920 7340 15972
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 8852 15988 8904 16040
rect 10232 16056 10284 16108
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10048 16031 10100 16040
rect 10048 15997 10057 16031
rect 10057 15997 10091 16031
rect 10091 15997 10100 16031
rect 10048 15988 10100 15997
rect 11060 15988 11112 16040
rect 12072 16192 12124 16244
rect 13084 16192 13136 16244
rect 14372 16192 14424 16244
rect 15200 16192 15252 16244
rect 15476 16192 15528 16244
rect 17316 16192 17368 16244
rect 18052 16192 18104 16244
rect 18788 16192 18840 16244
rect 19156 16192 19208 16244
rect 20812 16192 20864 16244
rect 21456 16192 21508 16244
rect 23480 16192 23532 16244
rect 24676 16235 24728 16244
rect 24676 16201 24685 16235
rect 24685 16201 24719 16235
rect 24719 16201 24728 16235
rect 24676 16192 24728 16201
rect 27436 16192 27488 16244
rect 28632 16192 28684 16244
rect 29460 16192 29512 16244
rect 30104 16235 30156 16244
rect 30104 16201 30113 16235
rect 30113 16201 30147 16235
rect 30147 16201 30156 16235
rect 30104 16192 30156 16201
rect 11336 16124 11388 16176
rect 11796 16056 11848 16108
rect 16396 16124 16448 16176
rect 16764 16124 16816 16176
rect 11428 15988 11480 16040
rect 7564 15852 7616 15904
rect 12072 15988 12124 16040
rect 16120 16056 16172 16108
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 16856 16056 16908 16108
rect 17316 16056 17368 16108
rect 18144 16056 18196 16108
rect 18328 16056 18380 16108
rect 18880 16056 18932 16108
rect 19340 16056 19392 16108
rect 19892 16056 19944 16108
rect 12624 15920 12676 15972
rect 13268 15920 13320 15972
rect 13912 15988 13964 16040
rect 14832 15988 14884 16040
rect 14924 15920 14976 15972
rect 15384 15920 15436 15972
rect 16212 15988 16264 16040
rect 16948 15988 17000 16040
rect 17408 15988 17460 16040
rect 17592 15988 17644 16040
rect 17868 16031 17920 16040
rect 17868 15997 17877 16031
rect 17877 15997 17911 16031
rect 17911 15997 17920 16031
rect 17868 15988 17920 15997
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 18604 15988 18656 16040
rect 16672 15920 16724 15972
rect 16856 15963 16908 15972
rect 16856 15929 16865 15963
rect 16865 15929 16899 15963
rect 16899 15929 16908 15963
rect 16856 15920 16908 15929
rect 20168 15988 20220 16040
rect 22100 15988 22152 16040
rect 12900 15852 12952 15904
rect 13360 15852 13412 15904
rect 15108 15852 15160 15904
rect 16212 15852 16264 15904
rect 18052 15852 18104 15904
rect 22468 15895 22520 15904
rect 22468 15861 22477 15895
rect 22477 15861 22511 15895
rect 22511 15861 22520 15895
rect 22468 15852 22520 15861
rect 25228 16099 25280 16108
rect 25228 16065 25237 16099
rect 25237 16065 25271 16099
rect 25271 16065 25280 16099
rect 25228 16056 25280 16065
rect 30012 16056 30064 16108
rect 24308 15988 24360 16040
rect 26056 15988 26108 16040
rect 23480 15920 23532 15972
rect 23756 15920 23808 15972
rect 25780 15920 25832 15972
rect 26608 15895 26660 15904
rect 26608 15861 26617 15895
rect 26617 15861 26651 15895
rect 26651 15861 26660 15895
rect 26608 15852 26660 15861
rect 27712 15920 27764 15972
rect 29184 15920 29236 15972
rect 27528 15852 27580 15904
rect 30932 15852 30984 15904
rect 11253 15750 11305 15802
rect 11317 15750 11369 15802
rect 11381 15750 11433 15802
rect 11445 15750 11497 15802
rect 11509 15750 11561 15802
rect 21557 15750 21609 15802
rect 21621 15750 21673 15802
rect 21685 15750 21737 15802
rect 21749 15750 21801 15802
rect 21813 15750 21865 15802
rect 2964 15648 3016 15700
rect 4712 15648 4764 15700
rect 8392 15648 8444 15700
rect 9680 15648 9732 15700
rect 10692 15691 10744 15700
rect 10692 15657 10701 15691
rect 10701 15657 10735 15691
rect 10735 15657 10744 15691
rect 10692 15648 10744 15657
rect 15384 15691 15436 15700
rect 1492 15512 1544 15564
rect 2688 15580 2740 15632
rect 3700 15580 3752 15632
rect 2504 15555 2556 15564
rect 2504 15521 2538 15555
rect 2538 15521 2556 15555
rect 2504 15512 2556 15521
rect 3792 15512 3844 15564
rect 5264 15555 5316 15564
rect 5264 15521 5273 15555
rect 5273 15521 5307 15555
rect 5307 15521 5316 15555
rect 5264 15512 5316 15521
rect 8484 15580 8536 15632
rect 9588 15623 9640 15632
rect 9588 15589 9622 15623
rect 9622 15589 9640 15623
rect 9588 15580 9640 15589
rect 7380 15512 7432 15564
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 4988 15444 5040 15496
rect 5632 15444 5684 15496
rect 7564 15444 7616 15496
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 11888 15580 11940 15632
rect 13268 15580 13320 15632
rect 14096 15580 14148 15632
rect 3884 15376 3936 15428
rect 8300 15444 8352 15496
rect 8852 15487 8904 15496
rect 8852 15453 8861 15487
rect 8861 15453 8895 15487
rect 8895 15453 8904 15487
rect 8852 15444 8904 15453
rect 12072 15512 12124 15564
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 14648 15555 14700 15564
rect 14648 15521 14657 15555
rect 14657 15521 14691 15555
rect 14691 15521 14700 15555
rect 14648 15512 14700 15521
rect 15108 15580 15160 15632
rect 15384 15657 15393 15691
rect 15393 15657 15427 15691
rect 15427 15657 15436 15691
rect 15384 15648 15436 15657
rect 15568 15648 15620 15700
rect 16396 15648 16448 15700
rect 15200 15555 15252 15564
rect 9220 15444 9272 15496
rect 1492 15308 1544 15360
rect 4344 15308 4396 15360
rect 4712 15308 4764 15360
rect 5816 15308 5868 15360
rect 7288 15308 7340 15360
rect 14740 15376 14792 15428
rect 15200 15521 15209 15555
rect 15209 15521 15243 15555
rect 15243 15521 15252 15555
rect 15200 15512 15252 15521
rect 15292 15444 15344 15496
rect 15476 15376 15528 15428
rect 15936 15512 15988 15564
rect 16672 15512 16724 15564
rect 17960 15512 18012 15564
rect 18144 15555 18196 15564
rect 18144 15521 18153 15555
rect 18153 15521 18187 15555
rect 18187 15521 18196 15555
rect 18144 15512 18196 15521
rect 18236 15512 18288 15564
rect 18972 15555 19024 15564
rect 18972 15521 18981 15555
rect 18981 15521 19015 15555
rect 19015 15521 19024 15555
rect 19248 15555 19300 15564
rect 18972 15512 19024 15521
rect 19248 15521 19257 15555
rect 19257 15521 19291 15555
rect 19291 15521 19300 15555
rect 19248 15512 19300 15521
rect 19524 15512 19576 15564
rect 19064 15487 19116 15496
rect 19064 15453 19073 15487
rect 19073 15453 19107 15487
rect 19107 15453 19116 15487
rect 19064 15444 19116 15453
rect 19800 15444 19852 15496
rect 22100 15691 22152 15700
rect 22100 15657 22109 15691
rect 22109 15657 22143 15691
rect 22143 15657 22152 15691
rect 23572 15691 23624 15700
rect 22100 15648 22152 15657
rect 23572 15657 23581 15691
rect 23581 15657 23615 15691
rect 23615 15657 23624 15691
rect 23572 15648 23624 15657
rect 24952 15648 25004 15700
rect 27712 15691 27764 15700
rect 27712 15657 27721 15691
rect 27721 15657 27755 15691
rect 27755 15657 27764 15691
rect 27712 15648 27764 15657
rect 30564 15648 30616 15700
rect 31024 15691 31076 15700
rect 31024 15657 31049 15691
rect 31049 15657 31076 15691
rect 31024 15648 31076 15657
rect 22284 15623 22336 15632
rect 22284 15589 22311 15623
rect 22311 15589 22336 15623
rect 22284 15580 22336 15589
rect 22376 15580 22428 15632
rect 20628 15555 20680 15564
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 28172 15623 28224 15632
rect 23112 15555 23164 15564
rect 22468 15444 22520 15496
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 23940 15512 23992 15564
rect 24308 15512 24360 15564
rect 26516 15512 26568 15564
rect 28172 15589 28181 15623
rect 28181 15589 28215 15623
rect 28215 15589 28224 15623
rect 28172 15580 28224 15589
rect 30932 15580 30984 15632
rect 23664 15444 23716 15496
rect 24768 15487 24820 15496
rect 24768 15453 24777 15487
rect 24777 15453 24811 15487
rect 24811 15453 24820 15487
rect 24768 15444 24820 15453
rect 26608 15444 26660 15496
rect 27436 15512 27488 15564
rect 27252 15487 27304 15496
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 9588 15308 9640 15360
rect 12164 15308 12216 15360
rect 13544 15308 13596 15360
rect 14004 15308 14056 15360
rect 15108 15308 15160 15360
rect 15384 15308 15436 15360
rect 17592 15376 17644 15428
rect 18972 15376 19024 15428
rect 20260 15419 20312 15428
rect 20260 15385 20269 15419
rect 20269 15385 20303 15419
rect 20303 15385 20312 15419
rect 20260 15376 20312 15385
rect 24676 15376 24728 15428
rect 29184 15512 29236 15564
rect 29276 15555 29328 15564
rect 29276 15521 29285 15555
rect 29285 15521 29319 15555
rect 29319 15521 29328 15555
rect 29276 15512 29328 15521
rect 29552 15487 29604 15496
rect 29552 15453 29561 15487
rect 29561 15453 29595 15487
rect 29595 15453 29604 15487
rect 29552 15444 29604 15453
rect 28356 15376 28408 15428
rect 16856 15308 16908 15360
rect 19984 15308 20036 15360
rect 20536 15308 20588 15360
rect 22468 15308 22520 15360
rect 23940 15308 23992 15360
rect 24860 15308 24912 15360
rect 30840 15308 30892 15360
rect 31208 15351 31260 15360
rect 31208 15317 31217 15351
rect 31217 15317 31251 15351
rect 31251 15317 31260 15351
rect 31208 15308 31260 15317
rect 6102 15206 6154 15258
rect 6166 15206 6218 15258
rect 6230 15206 6282 15258
rect 6294 15206 6346 15258
rect 6358 15206 6410 15258
rect 16405 15206 16457 15258
rect 16469 15206 16521 15258
rect 16533 15206 16585 15258
rect 16597 15206 16649 15258
rect 16661 15206 16713 15258
rect 26709 15206 26761 15258
rect 26773 15206 26825 15258
rect 26837 15206 26889 15258
rect 26901 15206 26953 15258
rect 26965 15206 27017 15258
rect 1676 15104 1728 15156
rect 4528 15104 4580 15156
rect 4712 15104 4764 15156
rect 6000 15036 6052 15088
rect 5540 15011 5592 15020
rect 5540 14977 5549 15011
rect 5549 14977 5583 15011
rect 5583 14977 5592 15011
rect 5540 14968 5592 14977
rect 6736 15036 6788 15088
rect 7840 15104 7892 15156
rect 8852 15104 8904 15156
rect 10324 15104 10376 15156
rect 11704 15104 11756 15156
rect 12900 15104 12952 15156
rect 13452 15147 13504 15156
rect 13452 15113 13461 15147
rect 13461 15113 13495 15147
rect 13495 15113 13504 15147
rect 13452 15104 13504 15113
rect 14464 15104 14516 15156
rect 15200 15104 15252 15156
rect 15660 15147 15712 15156
rect 15660 15113 15669 15147
rect 15669 15113 15703 15147
rect 15703 15113 15712 15147
rect 15660 15104 15712 15113
rect 10048 15036 10100 15088
rect 16212 15036 16264 15088
rect 18144 15104 18196 15156
rect 18328 15036 18380 15088
rect 18604 15104 18656 15156
rect 19616 15104 19668 15156
rect 19248 15036 19300 15088
rect 19340 15036 19392 15088
rect 19984 15104 20036 15156
rect 20168 15104 20220 15156
rect 20628 15104 20680 15156
rect 22928 15104 22980 15156
rect 23756 15104 23808 15156
rect 24308 15104 24360 15156
rect 24860 15104 24912 15156
rect 25780 15147 25832 15156
rect 25780 15113 25789 15147
rect 25789 15113 25823 15147
rect 25823 15113 25832 15147
rect 25780 15104 25832 15113
rect 27068 15104 27120 15156
rect 28356 15147 28408 15156
rect 20352 15036 20404 15088
rect 23664 15036 23716 15088
rect 24584 15036 24636 15088
rect 24952 15036 25004 15088
rect 28356 15113 28365 15147
rect 28365 15113 28399 15147
rect 28399 15113 28408 15147
rect 28356 15104 28408 15113
rect 30012 15104 30064 15156
rect 7288 15011 7340 15020
rect 2228 14900 2280 14952
rect 4804 14943 4856 14952
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 5816 14943 5868 14952
rect 5816 14909 5825 14943
rect 5825 14909 5859 14943
rect 5859 14909 5868 14943
rect 5816 14900 5868 14909
rect 1768 14832 1820 14884
rect 3240 14832 3292 14884
rect 5264 14832 5316 14884
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 7748 14943 7800 14952
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 7748 14900 7800 14909
rect 8668 14968 8720 15020
rect 2412 14764 2464 14816
rect 2596 14764 2648 14816
rect 3792 14764 3844 14816
rect 4252 14807 4304 14816
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 7196 14832 7248 14884
rect 7564 14832 7616 14884
rect 8208 14900 8260 14952
rect 9772 14968 9824 15020
rect 9680 14900 9732 14952
rect 10140 14900 10192 14952
rect 11060 14900 11112 14952
rect 13544 14943 13596 14952
rect 8024 14764 8076 14816
rect 8760 14832 8812 14884
rect 9772 14832 9824 14884
rect 10784 14832 10836 14884
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 14464 14900 14516 14952
rect 17040 14900 17092 14952
rect 18144 14943 18196 14952
rect 15568 14832 15620 14884
rect 15660 14832 15712 14884
rect 15936 14832 15988 14884
rect 13820 14764 13872 14816
rect 15752 14764 15804 14816
rect 16304 14764 16356 14816
rect 16764 14832 16816 14884
rect 18144 14909 18153 14943
rect 18153 14909 18187 14943
rect 18187 14909 18196 14943
rect 18144 14900 18196 14909
rect 18328 14900 18380 14952
rect 18420 14832 18472 14884
rect 18972 14900 19024 14952
rect 19340 14900 19392 14952
rect 20812 14968 20864 15020
rect 22836 14968 22888 15020
rect 19616 14832 19668 14884
rect 20168 14832 20220 14884
rect 21456 14875 21508 14884
rect 21456 14841 21490 14875
rect 21490 14841 21508 14875
rect 21456 14832 21508 14841
rect 18236 14764 18288 14816
rect 19892 14764 19944 14816
rect 19984 14764 20036 14816
rect 22468 14764 22520 14816
rect 22652 14764 22704 14816
rect 23112 14900 23164 14952
rect 23756 14900 23808 14952
rect 24032 14900 24084 14952
rect 24676 14968 24728 15020
rect 26608 14968 26660 15020
rect 26148 14943 26200 14952
rect 26148 14909 26157 14943
rect 26157 14909 26191 14943
rect 26191 14909 26200 14943
rect 26148 14900 26200 14909
rect 24768 14832 24820 14884
rect 24860 14764 24912 14816
rect 25964 14764 26016 14816
rect 26332 14943 26384 14952
rect 26332 14909 26341 14943
rect 26341 14909 26375 14943
rect 26375 14909 26384 14943
rect 26332 14900 26384 14909
rect 26516 14943 26568 14952
rect 26516 14909 26525 14943
rect 26525 14909 26559 14943
rect 26559 14909 26568 14943
rect 26516 14900 26568 14909
rect 28724 15036 28776 15088
rect 29736 14900 29788 14952
rect 30288 14832 30340 14884
rect 30380 14832 30432 14884
rect 30564 14764 30616 14816
rect 11253 14662 11305 14714
rect 11317 14662 11369 14714
rect 11381 14662 11433 14714
rect 11445 14662 11497 14714
rect 11509 14662 11561 14714
rect 21557 14662 21609 14714
rect 21621 14662 21673 14714
rect 21685 14662 21737 14714
rect 21749 14662 21801 14714
rect 21813 14662 21865 14714
rect 2596 14560 2648 14612
rect 2780 14560 2832 14612
rect 3240 14560 3292 14612
rect 2136 14492 2188 14544
rect 2872 14492 2924 14544
rect 5632 14560 5684 14612
rect 7656 14603 7708 14612
rect 7656 14569 7665 14603
rect 7665 14569 7699 14603
rect 7699 14569 7708 14603
rect 7656 14560 7708 14569
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 10140 14603 10192 14612
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 10600 14603 10652 14612
rect 10600 14569 10609 14603
rect 10609 14569 10643 14603
rect 10643 14569 10652 14603
rect 10600 14560 10652 14569
rect 12256 14560 12308 14612
rect 12624 14560 12676 14612
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 15752 14560 15804 14612
rect 19064 14560 19116 14612
rect 19248 14560 19300 14612
rect 2780 14424 2832 14476
rect 4160 14492 4212 14544
rect 4252 14467 4304 14476
rect 2412 14356 2464 14408
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 5080 14492 5132 14544
rect 4988 14467 5040 14476
rect 4988 14433 4997 14467
rect 4997 14433 5031 14467
rect 5031 14433 5040 14467
rect 4988 14424 5040 14433
rect 5264 14424 5316 14476
rect 6000 14492 6052 14544
rect 6644 14424 6696 14476
rect 3884 14356 3936 14408
rect 4068 14356 4120 14408
rect 4344 14356 4396 14408
rect 5080 14356 5132 14408
rect 5356 14356 5408 14408
rect 6460 14356 6512 14408
rect 7012 14424 7064 14476
rect 7564 14467 7616 14476
rect 7564 14433 7573 14467
rect 7573 14433 7607 14467
rect 7607 14433 7616 14467
rect 7564 14424 7616 14433
rect 7840 14492 7892 14544
rect 8116 14424 8168 14476
rect 8484 14424 8536 14476
rect 12072 14492 12124 14544
rect 14372 14492 14424 14544
rect 15200 14492 15252 14544
rect 16856 14492 16908 14544
rect 18052 14535 18104 14544
rect 18052 14501 18086 14535
rect 18086 14501 18104 14535
rect 18052 14492 18104 14501
rect 13360 14467 13412 14476
rect 13360 14433 13394 14467
rect 13394 14433 13412 14467
rect 7380 14356 7432 14408
rect 8208 14356 8260 14408
rect 5816 14288 5868 14340
rect 4252 14220 4304 14272
rect 4528 14220 4580 14272
rect 5540 14220 5592 14272
rect 5632 14220 5684 14272
rect 6736 14288 6788 14340
rect 7104 14288 7156 14340
rect 8760 14288 8812 14340
rect 6460 14220 6512 14272
rect 7932 14220 7984 14272
rect 13360 14424 13412 14433
rect 14648 14424 14700 14476
rect 15108 14467 15160 14476
rect 15108 14433 15117 14467
rect 15117 14433 15151 14467
rect 15151 14433 15160 14467
rect 15108 14424 15160 14433
rect 15292 14467 15344 14476
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 15476 14467 15528 14476
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 19984 14560 20036 14612
rect 15476 14424 15528 14433
rect 19524 14424 19576 14476
rect 20812 14492 20864 14544
rect 19892 14424 19944 14476
rect 22468 14560 22520 14612
rect 24032 14603 24084 14612
rect 23480 14492 23532 14544
rect 24032 14569 24041 14603
rect 24041 14569 24075 14603
rect 24075 14569 24084 14603
rect 24032 14560 24084 14569
rect 24676 14560 24728 14612
rect 24860 14560 24912 14612
rect 28448 14560 28500 14612
rect 28724 14560 28776 14612
rect 30380 14603 30432 14612
rect 30380 14569 30389 14603
rect 30389 14569 30423 14603
rect 30423 14569 30432 14603
rect 30380 14560 30432 14569
rect 31484 14560 31536 14612
rect 25136 14492 25188 14544
rect 26148 14492 26200 14544
rect 15384 14356 15436 14408
rect 16764 14356 16816 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 23388 14424 23440 14476
rect 24584 14424 24636 14476
rect 24952 14424 25004 14476
rect 25320 14424 25372 14476
rect 25596 14424 25648 14476
rect 24768 14399 24820 14408
rect 14096 14288 14148 14340
rect 17408 14288 17460 14340
rect 12256 14220 12308 14272
rect 14004 14220 14056 14272
rect 14924 14220 14976 14272
rect 16856 14220 16908 14272
rect 17132 14220 17184 14272
rect 17960 14220 18012 14272
rect 18052 14220 18104 14272
rect 19524 14288 19576 14340
rect 19064 14220 19116 14272
rect 21180 14220 21232 14272
rect 21640 14220 21692 14272
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 25136 14356 25188 14408
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 26332 14424 26384 14476
rect 27160 14424 27212 14476
rect 28632 14467 28684 14476
rect 28632 14433 28641 14467
rect 28641 14433 28675 14467
rect 28675 14433 28684 14467
rect 28632 14424 28684 14433
rect 29552 14492 29604 14544
rect 26148 14356 26200 14408
rect 28172 14356 28224 14408
rect 22928 14220 22980 14272
rect 23296 14220 23348 14272
rect 24860 14220 24912 14272
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 25596 14220 25648 14272
rect 26516 14288 26568 14340
rect 28448 14288 28500 14340
rect 29644 14467 29696 14476
rect 29644 14433 29653 14467
rect 29653 14433 29687 14467
rect 29687 14433 29696 14467
rect 29644 14424 29696 14433
rect 29828 14467 29880 14476
rect 29828 14433 29837 14467
rect 29837 14433 29871 14467
rect 29871 14433 29880 14467
rect 29828 14424 29880 14433
rect 30012 14492 30064 14544
rect 30472 14424 30524 14476
rect 31116 14467 31168 14476
rect 31116 14433 31125 14467
rect 31125 14433 31159 14467
rect 31159 14433 31168 14467
rect 31116 14424 31168 14433
rect 30104 14356 30156 14408
rect 30748 14356 30800 14408
rect 31208 14356 31260 14408
rect 26424 14263 26476 14272
rect 26424 14229 26433 14263
rect 26433 14229 26467 14263
rect 26467 14229 26476 14263
rect 26424 14220 26476 14229
rect 27068 14263 27120 14272
rect 27068 14229 27077 14263
rect 27077 14229 27111 14263
rect 27111 14229 27120 14263
rect 27068 14220 27120 14229
rect 29184 14263 29236 14272
rect 29184 14229 29193 14263
rect 29193 14229 29227 14263
rect 29227 14229 29236 14263
rect 29184 14220 29236 14229
rect 29920 14220 29972 14272
rect 6102 14118 6154 14170
rect 6166 14118 6218 14170
rect 6230 14118 6282 14170
rect 6294 14118 6346 14170
rect 6358 14118 6410 14170
rect 16405 14118 16457 14170
rect 16469 14118 16521 14170
rect 16533 14118 16585 14170
rect 16597 14118 16649 14170
rect 16661 14118 16713 14170
rect 26709 14118 26761 14170
rect 26773 14118 26825 14170
rect 26837 14118 26889 14170
rect 26901 14118 26953 14170
rect 26965 14118 27017 14170
rect 1768 14016 1820 14068
rect 2044 14016 2096 14068
rect 2412 14016 2464 14068
rect 2136 13948 2188 14000
rect 2964 13948 3016 14000
rect 3884 13948 3936 14000
rect 3332 13880 3384 13932
rect 2228 13812 2280 13864
rect 1400 13744 1452 13796
rect 2780 13812 2832 13864
rect 3884 13812 3936 13864
rect 4896 14016 4948 14068
rect 6736 14016 6788 14068
rect 8116 14016 8168 14068
rect 8208 14016 8260 14068
rect 4528 13948 4580 14000
rect 7104 13948 7156 14000
rect 7932 13948 7984 14000
rect 8024 13948 8076 14000
rect 10600 14016 10652 14068
rect 13360 14016 13412 14068
rect 14372 14016 14424 14068
rect 16120 14016 16172 14068
rect 16856 14016 16908 14068
rect 19708 14016 19760 14068
rect 20904 14059 20956 14068
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 21272 14016 21324 14068
rect 21456 14016 21508 14068
rect 21916 14016 21968 14068
rect 23020 14016 23072 14068
rect 23388 14059 23440 14068
rect 23388 14025 23397 14059
rect 23397 14025 23431 14059
rect 23431 14025 23440 14059
rect 23388 14016 23440 14025
rect 16580 13948 16632 14000
rect 21640 13991 21692 14000
rect 5632 13880 5684 13932
rect 10692 13880 10744 13932
rect 12900 13880 12952 13932
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 2412 13676 2464 13728
rect 3884 13676 3936 13728
rect 4068 13676 4120 13728
rect 4160 13676 4212 13728
rect 5448 13812 5500 13864
rect 6460 13812 6512 13864
rect 6644 13812 6696 13864
rect 6920 13812 6972 13864
rect 7104 13812 7156 13864
rect 7564 13812 7616 13864
rect 8760 13812 8812 13864
rect 9588 13855 9640 13864
rect 9588 13821 9597 13855
rect 9597 13821 9631 13855
rect 9631 13821 9640 13855
rect 9588 13812 9640 13821
rect 4804 13744 4856 13796
rect 5080 13744 5132 13796
rect 5264 13787 5316 13796
rect 5264 13753 5273 13787
rect 5273 13753 5307 13787
rect 5307 13753 5316 13787
rect 5264 13744 5316 13753
rect 8668 13744 8720 13796
rect 9864 13787 9916 13796
rect 9864 13753 9898 13787
rect 9898 13753 9916 13787
rect 11060 13812 11112 13864
rect 12992 13855 13044 13864
rect 12992 13821 13001 13855
rect 13001 13821 13035 13855
rect 13035 13821 13044 13855
rect 12992 13812 13044 13821
rect 14004 13880 14056 13932
rect 14648 13880 14700 13932
rect 15108 13880 15160 13932
rect 14096 13812 14148 13864
rect 15200 13812 15252 13864
rect 16396 13880 16448 13932
rect 15752 13812 15804 13864
rect 16672 13880 16724 13932
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 21640 13957 21649 13991
rect 21649 13957 21683 13991
rect 21683 13957 21692 13991
rect 21640 13948 21692 13957
rect 22100 13948 22152 14000
rect 25688 14016 25740 14068
rect 27160 14059 27212 14068
rect 18328 13880 18380 13932
rect 19524 13923 19576 13932
rect 19524 13889 19533 13923
rect 19533 13889 19567 13923
rect 19567 13889 19576 13923
rect 19524 13880 19576 13889
rect 24768 13948 24820 14000
rect 24860 13948 24912 14000
rect 27160 14025 27169 14059
rect 27169 14025 27203 14059
rect 27203 14025 27212 14059
rect 27160 14016 27212 14025
rect 27528 14016 27580 14068
rect 30748 14059 30800 14068
rect 30748 14025 30757 14059
rect 30757 14025 30791 14059
rect 30791 14025 30800 14059
rect 30748 14016 30800 14025
rect 28540 13948 28592 14000
rect 29828 13948 29880 14000
rect 30196 13948 30248 14000
rect 30840 13991 30892 14000
rect 30840 13957 30849 13991
rect 30849 13957 30883 13991
rect 30883 13957 30892 13991
rect 30840 13948 30892 13957
rect 9864 13744 9916 13753
rect 13268 13744 13320 13796
rect 14648 13744 14700 13796
rect 16488 13744 16540 13796
rect 17960 13855 18012 13864
rect 17960 13821 17969 13855
rect 17969 13821 18003 13855
rect 18003 13821 18012 13855
rect 17960 13812 18012 13821
rect 18052 13812 18104 13864
rect 21824 13855 21876 13864
rect 17224 13744 17276 13796
rect 18420 13744 18472 13796
rect 19984 13744 20036 13796
rect 21456 13744 21508 13796
rect 21824 13821 21833 13855
rect 21833 13821 21867 13855
rect 21867 13821 21876 13855
rect 21824 13812 21876 13821
rect 22652 13855 22704 13864
rect 22652 13821 22661 13855
rect 22661 13821 22695 13855
rect 22695 13821 22704 13855
rect 22652 13812 22704 13821
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 22928 13855 22980 13864
rect 22928 13821 22937 13855
rect 22937 13821 22971 13855
rect 22971 13821 22980 13855
rect 22928 13812 22980 13821
rect 23112 13812 23164 13864
rect 25136 13880 25188 13932
rect 22560 13744 22612 13796
rect 24952 13855 25004 13864
rect 24952 13821 24961 13855
rect 24961 13821 24995 13855
rect 24995 13821 25004 13855
rect 24952 13812 25004 13821
rect 25596 13812 25648 13864
rect 25872 13812 25924 13864
rect 26424 13812 26476 13864
rect 29000 13880 29052 13932
rect 30932 13880 30984 13932
rect 28172 13812 28224 13864
rect 27252 13744 27304 13796
rect 28448 13855 28500 13864
rect 28448 13821 28457 13855
rect 28457 13821 28491 13855
rect 28491 13821 28500 13855
rect 28448 13812 28500 13821
rect 28724 13812 28776 13864
rect 30380 13812 30432 13864
rect 30472 13812 30524 13864
rect 30656 13812 30708 13864
rect 6000 13676 6052 13728
rect 9956 13676 10008 13728
rect 10416 13676 10468 13728
rect 12716 13676 12768 13728
rect 13452 13676 13504 13728
rect 18236 13676 18288 13728
rect 20536 13676 20588 13728
rect 24768 13676 24820 13728
rect 25136 13719 25188 13728
rect 25136 13685 25145 13719
rect 25145 13685 25179 13719
rect 25179 13685 25188 13719
rect 25136 13676 25188 13685
rect 25688 13676 25740 13728
rect 27436 13676 27488 13728
rect 27896 13719 27948 13728
rect 27896 13685 27905 13719
rect 27905 13685 27939 13719
rect 27939 13685 27948 13719
rect 27896 13676 27948 13685
rect 11253 13574 11305 13626
rect 11317 13574 11369 13626
rect 11381 13574 11433 13626
rect 11445 13574 11497 13626
rect 11509 13574 11561 13626
rect 21557 13574 21609 13626
rect 21621 13574 21673 13626
rect 21685 13574 21737 13626
rect 21749 13574 21801 13626
rect 21813 13574 21865 13626
rect 1400 13515 1452 13524
rect 1400 13481 1409 13515
rect 1409 13481 1443 13515
rect 1443 13481 1452 13515
rect 1400 13472 1452 13481
rect 1676 13404 1728 13456
rect 2412 13404 2464 13456
rect 2688 13336 2740 13388
rect 4068 13472 4120 13524
rect 4252 13472 4304 13524
rect 5264 13472 5316 13524
rect 5724 13472 5776 13524
rect 5816 13515 5868 13524
rect 5816 13481 5825 13515
rect 5825 13481 5859 13515
rect 5859 13481 5868 13515
rect 5816 13472 5868 13481
rect 7748 13472 7800 13524
rect 9864 13472 9916 13524
rect 10324 13472 10376 13524
rect 13912 13472 13964 13524
rect 15476 13472 15528 13524
rect 16580 13472 16632 13524
rect 3884 13404 3936 13456
rect 4252 13336 4304 13388
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5080 13336 5132 13345
rect 6644 13404 6696 13456
rect 6828 13404 6880 13456
rect 6736 13379 6788 13388
rect 6736 13345 6745 13379
rect 6745 13345 6779 13379
rect 6779 13345 6788 13379
rect 6736 13336 6788 13345
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 8116 13336 8168 13388
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 14648 13404 14700 13456
rect 15660 13404 15712 13456
rect 10692 13336 10744 13388
rect 11612 13336 11664 13388
rect 13084 13336 13136 13388
rect 13544 13336 13596 13388
rect 1400 13268 1452 13320
rect 3332 13268 3384 13320
rect 3884 13268 3936 13320
rect 4712 13268 4764 13320
rect 5172 13268 5224 13320
rect 6920 13311 6972 13320
rect 6920 13277 6929 13311
rect 6929 13277 6963 13311
rect 6963 13277 6972 13311
rect 6920 13268 6972 13277
rect 1860 13132 1912 13184
rect 2136 13132 2188 13184
rect 4068 13200 4120 13252
rect 5448 13200 5500 13252
rect 6552 13200 6604 13252
rect 10600 13268 10652 13320
rect 11060 13268 11112 13320
rect 11152 13200 11204 13252
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4528 13132 4580 13141
rect 5172 13132 5224 13184
rect 5356 13132 5408 13184
rect 5724 13132 5776 13184
rect 5908 13132 5960 13184
rect 7288 13175 7340 13184
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 12900 13243 12952 13252
rect 12900 13209 12909 13243
rect 12909 13209 12943 13243
rect 12943 13209 12952 13243
rect 14832 13336 14884 13388
rect 15292 13336 15344 13388
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 16488 13404 16540 13456
rect 16948 13404 17000 13456
rect 16396 13336 16448 13388
rect 17592 13404 17644 13456
rect 17236 13381 17288 13388
rect 17236 13347 17245 13381
rect 17245 13347 17279 13381
rect 17279 13347 17288 13381
rect 17236 13336 17288 13347
rect 18144 13472 18196 13524
rect 19616 13472 19668 13524
rect 21180 13472 21232 13524
rect 22284 13472 22336 13524
rect 23112 13472 23164 13524
rect 18788 13404 18840 13456
rect 20168 13404 20220 13456
rect 21364 13404 21416 13456
rect 21548 13404 21600 13456
rect 21824 13404 21876 13456
rect 19524 13336 19576 13388
rect 19708 13336 19760 13388
rect 20720 13336 20772 13388
rect 22100 13336 22152 13388
rect 22376 13336 22428 13388
rect 12900 13200 12952 13209
rect 16120 13200 16172 13252
rect 16396 13200 16448 13252
rect 22468 13268 22520 13320
rect 11888 13132 11940 13184
rect 14188 13175 14240 13184
rect 14188 13141 14197 13175
rect 14197 13141 14231 13175
rect 14231 13141 14240 13175
rect 14188 13132 14240 13141
rect 15108 13132 15160 13184
rect 17408 13200 17460 13252
rect 18052 13200 18104 13252
rect 19340 13200 19392 13252
rect 23756 13472 23808 13524
rect 24952 13472 25004 13524
rect 23664 13404 23716 13456
rect 25136 13379 25188 13388
rect 30380 13472 30432 13524
rect 30564 13472 30616 13524
rect 25964 13404 26016 13456
rect 25136 13345 25154 13379
rect 25154 13345 25188 13379
rect 25136 13336 25188 13345
rect 27068 13336 27120 13388
rect 29184 13404 29236 13456
rect 29736 13379 29788 13388
rect 29736 13345 29745 13379
rect 29745 13345 29779 13379
rect 29779 13345 29788 13379
rect 29736 13336 29788 13345
rect 31208 13336 31260 13388
rect 26608 13268 26660 13320
rect 30840 13311 30892 13320
rect 30840 13277 30849 13311
rect 30849 13277 30883 13311
rect 30883 13277 30892 13311
rect 30840 13268 30892 13277
rect 16764 13132 16816 13184
rect 18144 13132 18196 13184
rect 20720 13132 20772 13184
rect 21456 13132 21508 13184
rect 21548 13132 21600 13184
rect 22284 13132 22336 13184
rect 22928 13132 22980 13184
rect 24768 13132 24820 13184
rect 25964 13175 26016 13184
rect 25964 13141 25973 13175
rect 25973 13141 26007 13175
rect 26007 13141 26016 13175
rect 25964 13132 26016 13141
rect 27068 13175 27120 13184
rect 27068 13141 27077 13175
rect 27077 13141 27111 13175
rect 27111 13141 27120 13175
rect 27068 13132 27120 13141
rect 28448 13132 28500 13184
rect 30288 13200 30340 13252
rect 30104 13132 30156 13184
rect 30748 13175 30800 13184
rect 30748 13141 30757 13175
rect 30757 13141 30791 13175
rect 30791 13141 30800 13175
rect 30748 13132 30800 13141
rect 6102 13030 6154 13082
rect 6166 13030 6218 13082
rect 6230 13030 6282 13082
rect 6294 13030 6346 13082
rect 6358 13030 6410 13082
rect 16405 13030 16457 13082
rect 16469 13030 16521 13082
rect 16533 13030 16585 13082
rect 16597 13030 16649 13082
rect 16661 13030 16713 13082
rect 26709 13030 26761 13082
rect 26773 13030 26825 13082
rect 26837 13030 26889 13082
rect 26901 13030 26953 13082
rect 26965 13030 27017 13082
rect 2780 12928 2832 12980
rect 3884 12928 3936 12980
rect 4988 12928 5040 12980
rect 5724 12928 5776 12980
rect 10324 12971 10376 12980
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 11612 12928 11664 12980
rect 2872 12860 2924 12912
rect 4252 12860 4304 12912
rect 6920 12860 6972 12912
rect 2688 12724 2740 12776
rect 4068 12724 4120 12776
rect 4252 12724 4304 12776
rect 4988 12792 5040 12844
rect 6552 12792 6604 12844
rect 12532 12860 12584 12912
rect 5080 12767 5132 12776
rect 5080 12733 5089 12767
rect 5089 12733 5123 12767
rect 5123 12733 5132 12767
rect 5080 12724 5132 12733
rect 6460 12724 6512 12776
rect 6644 12767 6696 12776
rect 6644 12733 6653 12767
rect 6653 12733 6687 12767
rect 6687 12733 6696 12767
rect 6644 12724 6696 12733
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 7196 12767 7248 12776
rect 1952 12656 2004 12708
rect 2596 12656 2648 12708
rect 3884 12656 3936 12708
rect 5540 12656 5592 12708
rect 5724 12656 5776 12708
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 7840 12767 7892 12776
rect 7840 12733 7849 12767
rect 7849 12733 7883 12767
rect 7883 12733 7892 12767
rect 7840 12724 7892 12733
rect 9588 12724 9640 12776
rect 10692 12724 10744 12776
rect 10876 12724 10928 12776
rect 7104 12656 7156 12708
rect 7656 12656 7708 12708
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 12900 12792 12952 12844
rect 15292 12860 15344 12912
rect 15384 12792 15436 12844
rect 11060 12724 11112 12733
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 14188 12724 14240 12776
rect 12716 12699 12768 12708
rect 12716 12665 12725 12699
rect 12725 12665 12759 12699
rect 12759 12665 12768 12699
rect 12716 12656 12768 12665
rect 13268 12656 13320 12708
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 15108 12724 15160 12776
rect 15476 12656 15528 12708
rect 16120 12928 16172 12980
rect 17776 12928 17828 12980
rect 18052 12928 18104 12980
rect 19984 12971 20036 12980
rect 19984 12937 19993 12971
rect 19993 12937 20027 12971
rect 20027 12937 20036 12971
rect 19984 12928 20036 12937
rect 16764 12767 16816 12776
rect 16764 12733 16782 12767
rect 16782 12733 16816 12767
rect 16764 12724 16816 12733
rect 16948 12724 17000 12776
rect 19524 12835 19576 12844
rect 19524 12801 19533 12835
rect 19533 12801 19567 12835
rect 19567 12801 19576 12835
rect 19524 12792 19576 12801
rect 20812 12860 20864 12912
rect 21272 12860 21324 12912
rect 22744 12928 22796 12980
rect 23664 12971 23716 12980
rect 23664 12937 23673 12971
rect 23673 12937 23707 12971
rect 23707 12937 23716 12971
rect 23664 12928 23716 12937
rect 24216 12928 24268 12980
rect 29000 12971 29052 12980
rect 22560 12860 22612 12912
rect 29000 12937 29009 12971
rect 29009 12937 29043 12971
rect 29043 12937 29052 12971
rect 29000 12928 29052 12937
rect 30288 12928 30340 12980
rect 22744 12792 22796 12844
rect 17224 12724 17276 12776
rect 17408 12724 17460 12776
rect 18144 12724 18196 12776
rect 19156 12724 19208 12776
rect 17960 12656 18012 12708
rect 19616 12767 19668 12776
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 20812 12724 20864 12776
rect 5080 12588 5132 12640
rect 7472 12588 7524 12640
rect 7932 12631 7984 12640
rect 7932 12597 7941 12631
rect 7941 12597 7975 12631
rect 7975 12597 7984 12631
rect 7932 12588 7984 12597
rect 9588 12588 9640 12640
rect 9772 12588 9824 12640
rect 10324 12588 10376 12640
rect 14372 12588 14424 12640
rect 14648 12588 14700 12640
rect 18052 12588 18104 12640
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 19708 12656 19760 12708
rect 21916 12724 21968 12776
rect 22468 12724 22520 12776
rect 22652 12724 22704 12776
rect 29092 12860 29144 12912
rect 25136 12792 25188 12844
rect 25504 12792 25556 12844
rect 24492 12767 24544 12776
rect 22192 12656 22244 12708
rect 22376 12656 22428 12708
rect 22928 12656 22980 12708
rect 24492 12733 24501 12767
rect 24501 12733 24535 12767
rect 24535 12733 24544 12767
rect 24492 12724 24544 12733
rect 25688 12724 25740 12776
rect 27252 12792 27304 12844
rect 30012 12835 30064 12844
rect 30012 12801 30021 12835
rect 30021 12801 30055 12835
rect 30055 12801 30064 12835
rect 30012 12792 30064 12801
rect 27068 12767 27120 12776
rect 27068 12733 27077 12767
rect 27077 12733 27111 12767
rect 27111 12733 27120 12767
rect 27068 12724 27120 12733
rect 27344 12724 27396 12776
rect 25412 12656 25464 12708
rect 25872 12656 25924 12708
rect 26056 12656 26108 12708
rect 29552 12724 29604 12776
rect 29644 12767 29696 12776
rect 29644 12733 29653 12767
rect 29653 12733 29687 12767
rect 29687 12733 29696 12767
rect 29644 12724 29696 12733
rect 27896 12699 27948 12708
rect 27896 12665 27930 12699
rect 27930 12665 27948 12699
rect 27896 12656 27948 12665
rect 29920 12767 29972 12776
rect 29920 12733 29929 12767
rect 29929 12733 29963 12767
rect 29963 12733 29972 12767
rect 30196 12767 30248 12776
rect 29920 12724 29972 12733
rect 30196 12733 30205 12767
rect 30205 12733 30239 12767
rect 30239 12733 30248 12767
rect 30196 12724 30248 12733
rect 30380 12724 30432 12776
rect 30840 12724 30892 12776
rect 20720 12588 20772 12640
rect 21180 12631 21232 12640
rect 21180 12597 21189 12631
rect 21189 12597 21223 12631
rect 21223 12597 21232 12631
rect 21180 12588 21232 12597
rect 21916 12631 21968 12640
rect 21916 12597 21941 12631
rect 21941 12597 21968 12631
rect 21916 12588 21968 12597
rect 25688 12588 25740 12640
rect 27528 12588 27580 12640
rect 30196 12588 30248 12640
rect 30840 12631 30892 12640
rect 30840 12597 30849 12631
rect 30849 12597 30883 12631
rect 30883 12597 30892 12631
rect 30840 12588 30892 12597
rect 31024 12631 31076 12640
rect 31024 12597 31041 12631
rect 31041 12597 31076 12631
rect 31024 12588 31076 12597
rect 11253 12486 11305 12538
rect 11317 12486 11369 12538
rect 11381 12486 11433 12538
rect 11445 12486 11497 12538
rect 11509 12486 11561 12538
rect 21557 12486 21609 12538
rect 21621 12486 21673 12538
rect 21685 12486 21737 12538
rect 21749 12486 21801 12538
rect 21813 12486 21865 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 1768 12384 1820 12436
rect 3608 12384 3660 12436
rect 3792 12427 3844 12436
rect 3792 12393 3801 12427
rect 3801 12393 3835 12427
rect 3835 12393 3844 12427
rect 3792 12384 3844 12393
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 2688 12248 2740 12300
rect 4160 12316 4212 12368
rect 5264 12316 5316 12368
rect 4528 12248 4580 12300
rect 5080 12248 5132 12300
rect 5356 12291 5408 12300
rect 5356 12257 5365 12291
rect 5365 12257 5399 12291
rect 5399 12257 5408 12291
rect 5356 12248 5408 12257
rect 5632 12248 5684 12300
rect 7932 12316 7984 12368
rect 6644 12248 6696 12300
rect 7196 12248 7248 12300
rect 8760 12248 8812 12300
rect 3976 12180 4028 12232
rect 5264 12180 5316 12232
rect 5816 12180 5868 12232
rect 7380 12180 7432 12232
rect 10048 12384 10100 12436
rect 10692 12384 10744 12436
rect 11796 12384 11848 12436
rect 12348 12384 12400 12436
rect 13268 12427 13320 12436
rect 13268 12393 13277 12427
rect 13277 12393 13311 12427
rect 13311 12393 13320 12427
rect 13268 12384 13320 12393
rect 15476 12427 15528 12436
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 15936 12427 15988 12436
rect 15936 12393 15945 12427
rect 15945 12393 15979 12427
rect 15979 12393 15988 12427
rect 15936 12384 15988 12393
rect 10324 12316 10376 12368
rect 12440 12316 12492 12368
rect 13360 12316 13412 12368
rect 14372 12359 14424 12368
rect 14372 12325 14406 12359
rect 14406 12325 14424 12359
rect 14372 12316 14424 12325
rect 17408 12316 17460 12368
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 12716 12291 12768 12300
rect 12716 12257 12725 12291
rect 12725 12257 12759 12291
rect 12759 12257 12768 12291
rect 12716 12248 12768 12257
rect 14004 12248 14056 12300
rect 18144 12384 18196 12436
rect 19432 12384 19484 12436
rect 17960 12316 18012 12368
rect 10324 12180 10376 12232
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 10692 12180 10744 12232
rect 11152 12180 11204 12232
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 15476 12180 15528 12232
rect 16028 12180 16080 12232
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 18420 12316 18472 12368
rect 18696 12316 18748 12368
rect 19156 12248 19208 12300
rect 20076 12316 20128 12368
rect 21916 12384 21968 12436
rect 23296 12384 23348 12436
rect 24492 12384 24544 12436
rect 25320 12384 25372 12436
rect 25412 12384 25464 12436
rect 25872 12384 25924 12436
rect 27344 12427 27396 12436
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 24584 12316 24636 12368
rect 25228 12316 25280 12368
rect 18420 12180 18472 12232
rect 19340 12180 19392 12232
rect 19432 12180 19484 12232
rect 13912 12112 13964 12164
rect 15936 12112 15988 12164
rect 19984 12180 20036 12232
rect 20812 12180 20864 12232
rect 20168 12112 20220 12164
rect 22100 12248 22152 12300
rect 22744 12291 22796 12300
rect 22744 12257 22753 12291
rect 22753 12257 22787 12291
rect 22787 12257 22796 12291
rect 23664 12291 23716 12300
rect 22744 12248 22796 12257
rect 23664 12257 23673 12291
rect 23673 12257 23707 12291
rect 23707 12257 23716 12291
rect 23664 12248 23716 12257
rect 26056 12291 26108 12300
rect 26056 12257 26065 12291
rect 26065 12257 26099 12291
rect 26099 12257 26108 12291
rect 26056 12248 26108 12257
rect 27344 12393 27353 12427
rect 27353 12393 27387 12427
rect 27387 12393 27396 12427
rect 27344 12384 27396 12393
rect 30288 12384 30340 12436
rect 30380 12384 30432 12436
rect 26608 12316 26660 12368
rect 27712 12316 27764 12368
rect 30196 12359 30248 12368
rect 30196 12325 30230 12359
rect 30230 12325 30248 12359
rect 30196 12316 30248 12325
rect 28448 12248 28500 12300
rect 29736 12248 29788 12300
rect 21364 12180 21416 12232
rect 21548 12180 21600 12232
rect 22928 12223 22980 12232
rect 22928 12189 22937 12223
rect 22937 12189 22971 12223
rect 22971 12189 22980 12223
rect 22928 12180 22980 12189
rect 24768 12180 24820 12232
rect 4160 12044 4212 12096
rect 4436 12044 4488 12096
rect 9220 12044 9272 12096
rect 9404 12044 9456 12096
rect 11704 12044 11756 12096
rect 12256 12044 12308 12096
rect 12900 12044 12952 12096
rect 16028 12044 16080 12096
rect 17408 12044 17460 12096
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 19892 12044 19944 12096
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 21824 12112 21876 12164
rect 24400 12044 24452 12096
rect 28632 12180 28684 12232
rect 29552 12180 29604 12232
rect 28356 12112 28408 12164
rect 29644 12112 29696 12164
rect 27160 12087 27212 12096
rect 27160 12053 27169 12087
rect 27169 12053 27203 12087
rect 27203 12053 27212 12087
rect 27160 12044 27212 12053
rect 27896 12044 27948 12096
rect 6102 11942 6154 11994
rect 6166 11942 6218 11994
rect 6230 11942 6282 11994
rect 6294 11942 6346 11994
rect 6358 11942 6410 11994
rect 16405 11942 16457 11994
rect 16469 11942 16521 11994
rect 16533 11942 16585 11994
rect 16597 11942 16649 11994
rect 16661 11942 16713 11994
rect 26709 11942 26761 11994
rect 26773 11942 26825 11994
rect 26837 11942 26889 11994
rect 26901 11942 26953 11994
rect 26965 11942 27017 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 2780 11772 2832 11824
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 2872 11704 2924 11756
rect 3332 11704 3384 11756
rect 2320 11636 2372 11688
rect 2964 11636 3016 11688
rect 9496 11840 9548 11892
rect 9588 11883 9640 11892
rect 9588 11849 9597 11883
rect 9597 11849 9631 11883
rect 9631 11849 9640 11883
rect 13360 11883 13412 11892
rect 9588 11840 9640 11849
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 14556 11840 14608 11892
rect 15844 11840 15896 11892
rect 16120 11840 16172 11892
rect 5448 11815 5500 11824
rect 5448 11781 5457 11815
rect 5457 11781 5491 11815
rect 5491 11781 5500 11815
rect 5448 11772 5500 11781
rect 5540 11772 5592 11824
rect 10232 11772 10284 11824
rect 10508 11772 10560 11824
rect 13912 11772 13964 11824
rect 18604 11772 18656 11824
rect 6092 11704 6144 11756
rect 7012 11747 7064 11756
rect 4436 11636 4488 11688
rect 2044 11568 2096 11620
rect 3884 11568 3936 11620
rect 5448 11568 5500 11620
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 10416 11704 10468 11756
rect 15200 11704 15252 11756
rect 7288 11679 7340 11688
rect 7288 11645 7322 11679
rect 7322 11645 7340 11679
rect 9772 11679 9824 11688
rect 7288 11636 7340 11645
rect 9772 11645 9781 11679
rect 9781 11645 9815 11679
rect 9815 11645 9824 11679
rect 9772 11636 9824 11645
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 10324 11679 10376 11688
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 11796 11636 11848 11688
rect 11980 11679 12032 11688
rect 11980 11645 11989 11679
rect 11989 11645 12023 11679
rect 12023 11645 12032 11679
rect 19340 11704 19392 11756
rect 19616 11840 19668 11892
rect 19708 11772 19760 11824
rect 20628 11840 20680 11892
rect 21548 11840 21600 11892
rect 11980 11636 12032 11645
rect 2504 11500 2556 11552
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 7656 11500 7708 11552
rect 8484 11500 8536 11552
rect 10232 11568 10284 11620
rect 12256 11611 12308 11620
rect 12256 11577 12290 11611
rect 12290 11577 12308 11611
rect 12256 11568 12308 11577
rect 10600 11500 10652 11552
rect 11796 11500 11848 11552
rect 15016 11543 15068 11552
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 15752 11611 15804 11620
rect 15752 11577 15761 11611
rect 15761 11577 15795 11611
rect 15795 11577 15804 11611
rect 17132 11636 17184 11688
rect 17868 11636 17920 11688
rect 19156 11636 19208 11688
rect 19432 11679 19484 11688
rect 19432 11645 19441 11679
rect 19441 11645 19475 11679
rect 19475 11645 19484 11679
rect 19432 11636 19484 11645
rect 21272 11772 21324 11824
rect 22100 11883 22152 11892
rect 22100 11849 22109 11883
rect 22109 11849 22143 11883
rect 22143 11849 22152 11883
rect 24400 11883 24452 11892
rect 22100 11840 22152 11849
rect 24400 11849 24409 11883
rect 24409 11849 24443 11883
rect 24443 11849 24452 11883
rect 24400 11840 24452 11849
rect 24492 11840 24544 11892
rect 25412 11840 25464 11892
rect 20628 11704 20680 11756
rect 22192 11704 22244 11756
rect 25964 11772 26016 11824
rect 25320 11704 25372 11756
rect 25780 11704 25832 11756
rect 15752 11568 15804 11577
rect 16856 11568 16908 11620
rect 18236 11568 18288 11620
rect 16028 11500 16080 11552
rect 16948 11500 17000 11552
rect 17684 11500 17736 11552
rect 18420 11500 18472 11552
rect 22468 11636 22520 11688
rect 22836 11636 22888 11688
rect 24952 11679 25004 11688
rect 24952 11645 24961 11679
rect 24961 11645 24995 11679
rect 24995 11645 25004 11679
rect 24952 11636 25004 11645
rect 25688 11679 25740 11688
rect 25688 11645 25697 11679
rect 25697 11645 25731 11679
rect 25731 11645 25740 11679
rect 25688 11636 25740 11645
rect 25872 11679 25924 11688
rect 25872 11645 25881 11679
rect 25881 11645 25915 11679
rect 25915 11645 25924 11679
rect 25872 11636 25924 11645
rect 29828 11840 29880 11892
rect 30748 11840 30800 11892
rect 19800 11500 19852 11552
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 22928 11568 22980 11620
rect 26516 11636 26568 11688
rect 27160 11679 27212 11688
rect 27160 11645 27169 11679
rect 27169 11645 27203 11679
rect 27203 11645 27212 11679
rect 27160 11636 27212 11645
rect 27344 11636 27396 11688
rect 28724 11704 28776 11756
rect 29828 11747 29880 11756
rect 27896 11636 27948 11688
rect 28356 11636 28408 11688
rect 28448 11679 28500 11688
rect 28448 11645 28457 11679
rect 28457 11645 28491 11679
rect 28491 11645 28500 11679
rect 29828 11713 29837 11747
rect 29837 11713 29871 11747
rect 29871 11713 29880 11747
rect 29828 11704 29880 11713
rect 30012 11704 30064 11756
rect 30840 11747 30892 11756
rect 30840 11713 30849 11747
rect 30849 11713 30883 11747
rect 30883 11713 30892 11747
rect 30840 11704 30892 11713
rect 28448 11636 28500 11645
rect 27528 11568 27580 11620
rect 29736 11679 29788 11688
rect 29736 11645 29745 11679
rect 29745 11645 29779 11679
rect 29779 11645 29788 11679
rect 29736 11636 29788 11645
rect 30932 11636 30984 11688
rect 31116 11679 31168 11688
rect 31116 11645 31125 11679
rect 31125 11645 31159 11679
rect 31159 11645 31168 11679
rect 31116 11636 31168 11645
rect 21916 11543 21968 11552
rect 21916 11509 21925 11543
rect 21925 11509 21959 11543
rect 21959 11509 21968 11543
rect 21916 11500 21968 11509
rect 24308 11500 24360 11552
rect 26608 11500 26660 11552
rect 27068 11543 27120 11552
rect 27068 11509 27077 11543
rect 27077 11509 27111 11543
rect 27111 11509 27120 11543
rect 27068 11500 27120 11509
rect 27620 11543 27672 11552
rect 27620 11509 27629 11543
rect 27629 11509 27663 11543
rect 27663 11509 27672 11543
rect 27620 11500 27672 11509
rect 29644 11500 29696 11552
rect 30288 11543 30340 11552
rect 30288 11509 30297 11543
rect 30297 11509 30331 11543
rect 30331 11509 30340 11543
rect 30288 11500 30340 11509
rect 31116 11500 31168 11552
rect 11253 11398 11305 11450
rect 11317 11398 11369 11450
rect 11381 11398 11433 11450
rect 11445 11398 11497 11450
rect 11509 11398 11561 11450
rect 21557 11398 21609 11450
rect 21621 11398 21673 11450
rect 21685 11398 21737 11450
rect 21749 11398 21801 11450
rect 21813 11398 21865 11450
rect 2964 11296 3016 11348
rect 3332 11296 3384 11348
rect 4068 11296 4120 11348
rect 4620 11296 4672 11348
rect 4712 11296 4764 11348
rect 5080 11296 5132 11348
rect 5356 11296 5408 11348
rect 5816 11296 5868 11348
rect 6000 11296 6052 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 10048 11296 10100 11348
rect 12256 11296 12308 11348
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 1584 11160 1636 11212
rect 1768 11160 1820 11212
rect 2872 11228 2924 11280
rect 2320 11203 2372 11212
rect 2320 11169 2329 11203
rect 2329 11169 2363 11203
rect 2363 11169 2372 11203
rect 2320 11160 2372 11169
rect 2780 11160 2832 11212
rect 3884 11228 3936 11280
rect 4344 11228 4396 11280
rect 3240 11160 3292 11212
rect 6460 11228 6512 11280
rect 6736 11271 6788 11280
rect 6736 11237 6745 11271
rect 6745 11237 6779 11271
rect 6779 11237 6788 11271
rect 6736 11228 6788 11237
rect 7472 11228 7524 11280
rect 1860 11092 1912 11144
rect 1768 11067 1820 11076
rect 1768 11033 1777 11067
rect 1777 11033 1811 11067
rect 1811 11033 1820 11067
rect 1768 11024 1820 11033
rect 2872 11092 2924 11144
rect 3608 11092 3660 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 4804 11092 4856 11144
rect 5356 11160 5408 11212
rect 4344 11024 4396 11076
rect 4896 11024 4948 11076
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 3884 10956 3936 11008
rect 6460 11092 6512 11144
rect 6092 11024 6144 11076
rect 7012 11160 7064 11212
rect 9220 11203 9272 11212
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 16028 11296 16080 11348
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 16948 11271 17000 11280
rect 11796 11160 11848 11212
rect 12072 11160 12124 11212
rect 16948 11237 16957 11271
rect 16957 11237 16991 11271
rect 16991 11237 17000 11271
rect 16948 11228 17000 11237
rect 14556 11160 14608 11212
rect 14924 11160 14976 11212
rect 15936 11160 15988 11212
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 10692 11092 10744 11144
rect 14004 11092 14056 11144
rect 19064 11296 19116 11348
rect 20628 11296 20680 11348
rect 24124 11296 24176 11348
rect 24308 11339 24360 11348
rect 24308 11305 24317 11339
rect 24317 11305 24351 11339
rect 24351 11305 24360 11339
rect 24308 11296 24360 11305
rect 25872 11339 25924 11348
rect 25872 11305 25881 11339
rect 25881 11305 25915 11339
rect 25915 11305 25924 11339
rect 25872 11296 25924 11305
rect 27160 11339 27212 11348
rect 27160 11305 27169 11339
rect 27169 11305 27203 11339
rect 27203 11305 27212 11339
rect 27160 11296 27212 11305
rect 28448 11296 28500 11348
rect 29000 11296 29052 11348
rect 30656 11296 30708 11348
rect 17408 11092 17460 11144
rect 19984 11228 20036 11280
rect 23480 11228 23532 11280
rect 21272 11160 21324 11212
rect 22100 11203 22152 11212
rect 22100 11169 22109 11203
rect 22109 11169 22143 11203
rect 22143 11169 22152 11203
rect 22100 11160 22152 11169
rect 23204 11203 23256 11212
rect 23204 11169 23238 11203
rect 23238 11169 23256 11203
rect 24768 11203 24820 11212
rect 23204 11160 23256 11169
rect 24768 11169 24777 11203
rect 24777 11169 24811 11203
rect 24811 11169 24820 11203
rect 24768 11160 24820 11169
rect 25412 11203 25464 11212
rect 25412 11169 25421 11203
rect 25421 11169 25455 11203
rect 25455 11169 25464 11203
rect 25412 11160 25464 11169
rect 25780 11160 25832 11212
rect 25964 11160 26016 11212
rect 27344 11203 27396 11212
rect 27344 11169 27353 11203
rect 27353 11169 27387 11203
rect 27387 11169 27396 11203
rect 27344 11160 27396 11169
rect 27896 11228 27948 11280
rect 28908 11228 28960 11280
rect 27620 11203 27672 11212
rect 27620 11169 27629 11203
rect 27629 11169 27663 11203
rect 27663 11169 27672 11203
rect 27620 11160 27672 11169
rect 19156 11092 19208 11144
rect 22744 11092 22796 11144
rect 27528 11135 27580 11144
rect 27528 11101 27537 11135
rect 27537 11101 27571 11135
rect 27571 11101 27580 11135
rect 27528 11092 27580 11101
rect 25688 11024 25740 11076
rect 30472 11160 30524 11212
rect 31116 11203 31168 11212
rect 31116 11169 31125 11203
rect 31125 11169 31159 11203
rect 31159 11169 31168 11203
rect 31116 11160 31168 11169
rect 5908 10956 5960 11008
rect 6000 10956 6052 11008
rect 14188 10956 14240 11008
rect 15844 10956 15896 11008
rect 17408 10956 17460 11008
rect 18144 10956 18196 11008
rect 24952 10956 25004 11008
rect 25136 10956 25188 11008
rect 28908 10956 28960 11008
rect 29552 10999 29604 11008
rect 29552 10965 29561 10999
rect 29561 10965 29595 10999
rect 29595 10965 29604 10999
rect 29552 10956 29604 10965
rect 6102 10854 6154 10906
rect 6166 10854 6218 10906
rect 6230 10854 6282 10906
rect 6294 10854 6346 10906
rect 6358 10854 6410 10906
rect 16405 10854 16457 10906
rect 16469 10854 16521 10906
rect 16533 10854 16585 10906
rect 16597 10854 16649 10906
rect 16661 10854 16713 10906
rect 26709 10854 26761 10906
rect 26773 10854 26825 10906
rect 26837 10854 26889 10906
rect 26901 10854 26953 10906
rect 26965 10854 27017 10906
rect 2688 10752 2740 10804
rect 3608 10752 3660 10804
rect 3976 10795 4028 10804
rect 3976 10761 3985 10795
rect 3985 10761 4019 10795
rect 4019 10761 4028 10795
rect 3976 10752 4028 10761
rect 5816 10752 5868 10804
rect 2872 10616 2924 10668
rect 3148 10616 3200 10668
rect 3976 10616 4028 10668
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4620 10548 4672 10600
rect 5908 10684 5960 10736
rect 5816 10616 5868 10668
rect 5724 10591 5776 10600
rect 4436 10480 4488 10532
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 5724 10548 5776 10557
rect 6920 10616 6972 10668
rect 6184 10548 6236 10600
rect 6552 10548 6604 10600
rect 6828 10548 6880 10600
rect 10232 10752 10284 10804
rect 10784 10752 10836 10804
rect 13728 10752 13780 10804
rect 18696 10752 18748 10804
rect 9956 10684 10008 10736
rect 10416 10684 10468 10736
rect 17500 10684 17552 10736
rect 18236 10684 18288 10736
rect 19800 10752 19852 10804
rect 20444 10752 20496 10804
rect 20996 10752 21048 10804
rect 21916 10752 21968 10804
rect 24492 10795 24544 10804
rect 24492 10761 24501 10795
rect 24501 10761 24535 10795
rect 24535 10761 24544 10795
rect 24492 10752 24544 10761
rect 27988 10752 28040 10804
rect 29736 10752 29788 10804
rect 21088 10684 21140 10736
rect 21364 10684 21416 10736
rect 10140 10616 10192 10668
rect 8852 10548 8904 10600
rect 9680 10548 9732 10600
rect 10416 10548 10468 10600
rect 11704 10591 11756 10600
rect 11704 10557 11722 10591
rect 11722 10557 11756 10591
rect 11704 10548 11756 10557
rect 11888 10548 11940 10600
rect 17132 10616 17184 10668
rect 19616 10616 19668 10668
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 22008 10616 22060 10668
rect 25504 10616 25556 10668
rect 9312 10480 9364 10532
rect 12532 10548 12584 10600
rect 13912 10548 13964 10600
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 14740 10548 14792 10600
rect 17960 10591 18012 10600
rect 17960 10557 17969 10591
rect 17969 10557 18003 10591
rect 18003 10557 18012 10591
rect 17960 10548 18012 10557
rect 18144 10591 18196 10600
rect 18144 10557 18153 10591
rect 18153 10557 18187 10591
rect 18187 10557 18196 10591
rect 18144 10548 18196 10557
rect 18420 10548 18472 10600
rect 19340 10548 19392 10600
rect 12808 10480 12860 10532
rect 13360 10480 13412 10532
rect 14188 10480 14240 10532
rect 14372 10523 14424 10532
rect 14372 10489 14406 10523
rect 14406 10489 14424 10523
rect 14372 10480 14424 10489
rect 14556 10480 14608 10532
rect 5080 10412 5132 10464
rect 5908 10412 5960 10464
rect 6460 10455 6512 10464
rect 6460 10421 6469 10455
rect 6469 10421 6503 10455
rect 6503 10421 6512 10455
rect 6460 10412 6512 10421
rect 6736 10412 6788 10464
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7656 10455 7708 10464
rect 7656 10421 7665 10455
rect 7665 10421 7699 10455
rect 7699 10421 7708 10455
rect 7656 10412 7708 10421
rect 12992 10412 13044 10464
rect 15108 10412 15160 10464
rect 16764 10480 16816 10532
rect 19800 10480 19852 10532
rect 20352 10523 20404 10532
rect 20352 10489 20386 10523
rect 20386 10489 20404 10523
rect 22192 10548 22244 10600
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 22468 10548 22520 10557
rect 22560 10591 22612 10600
rect 22560 10557 22569 10591
rect 22569 10557 22603 10591
rect 22603 10557 22612 10591
rect 23112 10591 23164 10600
rect 22560 10548 22612 10557
rect 23112 10557 23121 10591
rect 23121 10557 23155 10591
rect 23155 10557 23164 10591
rect 23112 10548 23164 10557
rect 23480 10548 23532 10600
rect 24584 10548 24636 10600
rect 20352 10480 20404 10489
rect 22744 10480 22796 10532
rect 24032 10480 24084 10532
rect 25964 10523 26016 10532
rect 25964 10489 25973 10523
rect 25973 10489 26007 10523
rect 26007 10489 26016 10523
rect 25964 10480 26016 10489
rect 26516 10616 26568 10668
rect 26608 10591 26660 10600
rect 26608 10557 26617 10591
rect 26617 10557 26651 10591
rect 26651 10557 26660 10591
rect 26608 10548 26660 10557
rect 27436 10548 27488 10600
rect 29552 10591 29604 10600
rect 29552 10557 29561 10591
rect 29561 10557 29595 10591
rect 29595 10557 29604 10591
rect 29552 10548 29604 10557
rect 29644 10548 29696 10600
rect 28172 10480 28224 10532
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 22376 10412 22428 10464
rect 23388 10412 23440 10464
rect 25688 10412 25740 10464
rect 26148 10455 26200 10464
rect 26148 10421 26157 10455
rect 26157 10421 26191 10455
rect 26191 10421 26200 10455
rect 26148 10412 26200 10421
rect 28724 10412 28776 10464
rect 11253 10310 11305 10362
rect 11317 10310 11369 10362
rect 11381 10310 11433 10362
rect 11445 10310 11497 10362
rect 11509 10310 11561 10362
rect 21557 10310 21609 10362
rect 21621 10310 21673 10362
rect 21685 10310 21737 10362
rect 21749 10310 21801 10362
rect 21813 10310 21865 10362
rect 2044 10208 2096 10260
rect 2688 10208 2740 10260
rect 5356 10208 5408 10260
rect 6828 10208 6880 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 10232 10208 10284 10260
rect 2964 10140 3016 10192
rect 3148 10072 3200 10124
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 6460 10140 6512 10192
rect 7656 10140 7708 10192
rect 4712 10072 4764 10124
rect 5356 10115 5408 10124
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 5356 10072 5408 10081
rect 5448 10072 5500 10124
rect 10416 10208 10468 10260
rect 14372 10208 14424 10260
rect 17500 10208 17552 10260
rect 18052 10208 18104 10260
rect 19432 10251 19484 10260
rect 11888 10140 11940 10192
rect 12624 10140 12676 10192
rect 3792 10004 3844 10013
rect 2136 9868 2188 9920
rect 4712 9868 4764 9920
rect 7656 10004 7708 10056
rect 12716 10072 12768 10124
rect 13084 10072 13136 10124
rect 13728 10115 13780 10124
rect 13728 10081 13737 10115
rect 13737 10081 13771 10115
rect 13771 10081 13780 10115
rect 13728 10072 13780 10081
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 14004 10072 14056 10124
rect 14556 10072 14608 10124
rect 14832 10072 14884 10124
rect 19156 10140 19208 10192
rect 19432 10217 19441 10251
rect 19441 10217 19475 10251
rect 19475 10217 19484 10251
rect 19432 10208 19484 10217
rect 20352 10208 20404 10260
rect 21916 10208 21968 10260
rect 22284 10208 22336 10260
rect 23204 10251 23256 10260
rect 23204 10217 23213 10251
rect 23213 10217 23247 10251
rect 23247 10217 23256 10251
rect 23204 10208 23256 10217
rect 18696 10072 18748 10124
rect 19892 10072 19944 10124
rect 20812 10140 20864 10192
rect 30748 10208 30800 10260
rect 30932 10251 30984 10260
rect 30932 10217 30941 10251
rect 30941 10217 30975 10251
rect 30975 10217 30984 10251
rect 30932 10208 30984 10217
rect 24584 10140 24636 10192
rect 21456 10072 21508 10124
rect 21732 10072 21784 10124
rect 22284 10115 22336 10124
rect 22284 10081 22293 10115
rect 22293 10081 22327 10115
rect 22327 10081 22336 10115
rect 22284 10072 22336 10081
rect 22376 10072 22428 10124
rect 23388 10115 23440 10124
rect 23388 10081 23397 10115
rect 23397 10081 23431 10115
rect 23431 10081 23440 10115
rect 23388 10072 23440 10081
rect 24032 10115 24084 10124
rect 24032 10081 24041 10115
rect 24041 10081 24075 10115
rect 24075 10081 24084 10115
rect 24032 10072 24084 10081
rect 14372 10004 14424 10056
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 16028 10004 16080 10056
rect 17592 10004 17644 10056
rect 23020 10004 23072 10056
rect 14096 9936 14148 9988
rect 5632 9868 5684 9920
rect 7840 9868 7892 9920
rect 11152 9868 11204 9920
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 12624 9868 12676 9920
rect 12808 9868 12860 9920
rect 22100 9979 22152 9988
rect 22100 9945 22109 9979
rect 22109 9945 22143 9979
rect 22143 9945 22152 9979
rect 25320 10004 25372 10056
rect 29276 10140 29328 10192
rect 30288 10140 30340 10192
rect 25964 10072 26016 10124
rect 27344 10072 27396 10124
rect 29000 10004 29052 10056
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 22100 9936 22152 9945
rect 15752 9868 15804 9920
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 16856 9868 16908 9920
rect 21824 9911 21876 9920
rect 21824 9877 21833 9911
rect 21833 9877 21867 9911
rect 21867 9877 21876 9911
rect 21824 9868 21876 9877
rect 25044 9911 25096 9920
rect 25044 9877 25053 9911
rect 25053 9877 25087 9911
rect 25087 9877 25096 9911
rect 25044 9868 25096 9877
rect 26608 9936 26660 9988
rect 26424 9868 26476 9920
rect 27620 9868 27672 9920
rect 6102 9766 6154 9818
rect 6166 9766 6218 9818
rect 6230 9766 6282 9818
rect 6294 9766 6346 9818
rect 6358 9766 6410 9818
rect 16405 9766 16457 9818
rect 16469 9766 16521 9818
rect 16533 9766 16585 9818
rect 16597 9766 16649 9818
rect 16661 9766 16713 9818
rect 26709 9766 26761 9818
rect 26773 9766 26825 9818
rect 26837 9766 26889 9818
rect 26901 9766 26953 9818
rect 26965 9766 27017 9818
rect 3332 9664 3384 9716
rect 3884 9664 3936 9716
rect 4620 9664 4672 9716
rect 7012 9664 7064 9716
rect 14832 9707 14884 9716
rect 14832 9673 14841 9707
rect 14841 9673 14875 9707
rect 14875 9673 14884 9707
rect 14832 9664 14884 9673
rect 22100 9664 22152 9716
rect 23572 9707 23624 9716
rect 23572 9673 23581 9707
rect 23581 9673 23615 9707
rect 23615 9673 23624 9707
rect 23572 9664 23624 9673
rect 24492 9664 24544 9716
rect 27252 9664 27304 9716
rect 30012 9664 30064 9716
rect 4528 9596 4580 9648
rect 4988 9596 5040 9648
rect 6000 9596 6052 9648
rect 7380 9639 7432 9648
rect 7380 9605 7389 9639
rect 7389 9605 7423 9639
rect 7423 9605 7432 9639
rect 7380 9596 7432 9605
rect 10324 9596 10376 9648
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 2504 9503 2556 9512
rect 2504 9469 2522 9503
rect 2522 9469 2556 9503
rect 2504 9460 2556 9469
rect 3792 9460 3844 9512
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 6828 9528 6880 9580
rect 8392 9528 8444 9580
rect 12716 9528 12768 9580
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 5632 9460 5684 9512
rect 9128 9460 9180 9512
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 13176 9596 13228 9648
rect 15016 9596 15068 9648
rect 15568 9596 15620 9648
rect 16764 9639 16816 9648
rect 16764 9605 16773 9639
rect 16773 9605 16807 9639
rect 16807 9605 16816 9639
rect 16764 9596 16816 9605
rect 17960 9639 18012 9648
rect 17960 9605 17969 9639
rect 17969 9605 18003 9639
rect 18003 9605 18012 9639
rect 17960 9596 18012 9605
rect 19340 9596 19392 9648
rect 22192 9639 22244 9648
rect 22192 9605 22201 9639
rect 22201 9605 22235 9639
rect 22235 9605 22244 9639
rect 22192 9596 22244 9605
rect 30104 9639 30156 9648
rect 30104 9605 30113 9639
rect 30113 9605 30147 9639
rect 30147 9605 30156 9639
rect 30104 9596 30156 9605
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 12900 9460 12952 9512
rect 4896 9392 4948 9444
rect 2228 9324 2280 9376
rect 5632 9324 5684 9376
rect 6552 9392 6604 9444
rect 7380 9392 7432 9444
rect 6368 9324 6420 9376
rect 10968 9324 11020 9376
rect 11612 9324 11664 9376
rect 14004 9324 14056 9376
rect 15200 9469 15209 9490
rect 15209 9469 15243 9490
rect 15243 9469 15252 9490
rect 15200 9438 15252 9469
rect 16120 9528 16172 9580
rect 15660 9460 15712 9512
rect 16028 9503 16080 9512
rect 16028 9469 16037 9503
rect 16037 9469 16071 9503
rect 16071 9469 16080 9503
rect 16028 9460 16080 9469
rect 15292 9392 15344 9444
rect 17500 9460 17552 9512
rect 17132 9392 17184 9444
rect 19892 9460 19944 9512
rect 21824 9528 21876 9580
rect 20444 9460 20496 9512
rect 22008 9528 22060 9580
rect 22560 9460 22612 9512
rect 24032 9460 24084 9512
rect 24584 9460 24636 9512
rect 25320 9503 25372 9512
rect 25320 9469 25329 9503
rect 25329 9469 25363 9503
rect 25363 9469 25372 9503
rect 25320 9460 25372 9469
rect 27436 9528 27488 9580
rect 25964 9460 26016 9512
rect 26516 9460 26568 9512
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 16120 9324 16172 9376
rect 16304 9324 16356 9376
rect 16948 9324 17000 9376
rect 17500 9324 17552 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 20260 9324 20312 9376
rect 24860 9392 24912 9444
rect 26240 9392 26292 9444
rect 26884 9392 26936 9444
rect 26700 9324 26752 9376
rect 27528 9460 27580 9512
rect 29000 9503 29052 9512
rect 29000 9469 29009 9503
rect 29009 9469 29043 9503
rect 29043 9469 29052 9503
rect 29000 9460 29052 9469
rect 27528 9324 27580 9376
rect 28816 9324 28868 9376
rect 11253 9222 11305 9274
rect 11317 9222 11369 9274
rect 11381 9222 11433 9274
rect 11445 9222 11497 9274
rect 11509 9222 11561 9274
rect 21557 9222 21609 9274
rect 21621 9222 21673 9274
rect 21685 9222 21737 9274
rect 21749 9222 21801 9274
rect 21813 9222 21865 9274
rect 1676 9120 1728 9172
rect 2412 9120 2464 9172
rect 4804 9120 4856 9172
rect 5356 9120 5408 9172
rect 11704 9120 11756 9172
rect 16304 9120 16356 9172
rect 17316 9120 17368 9172
rect 17592 9120 17644 9172
rect 22100 9120 22152 9172
rect 22652 9120 22704 9172
rect 23480 9120 23532 9172
rect 2044 8984 2096 9036
rect 2228 8984 2280 9036
rect 2780 8984 2832 9036
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 4896 8984 4948 9036
rect 5080 8984 5132 9036
rect 5816 8984 5868 9036
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 7196 9052 7248 9104
rect 9128 9052 9180 9104
rect 6828 8984 6880 9036
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 8944 8984 8996 9036
rect 2228 8780 2280 8832
rect 4528 8848 4580 8900
rect 5540 8916 5592 8968
rect 6460 8916 6512 8968
rect 4252 8823 4304 8832
rect 4252 8789 4261 8823
rect 4261 8789 4295 8823
rect 4295 8789 4304 8823
rect 4252 8780 4304 8789
rect 4712 8780 4764 8832
rect 9128 8848 9180 8900
rect 11796 9052 11848 9104
rect 13452 9052 13504 9104
rect 16212 9052 16264 9104
rect 21180 9052 21232 9104
rect 23848 9095 23900 9104
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 11612 8984 11664 9036
rect 12348 9027 12400 9036
rect 11244 8916 11296 8968
rect 11612 8848 11664 8900
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 12440 8916 12492 8968
rect 13636 8984 13688 9036
rect 14004 8984 14056 9036
rect 14188 9027 14240 9036
rect 14188 8993 14197 9027
rect 14197 8993 14231 9027
rect 14231 8993 14240 9027
rect 14188 8984 14240 8993
rect 13084 8916 13136 8968
rect 17224 8984 17276 9036
rect 17684 9027 17736 9036
rect 17684 8993 17693 9027
rect 17693 8993 17727 9027
rect 17727 8993 17736 9027
rect 17684 8984 17736 8993
rect 18144 8984 18196 9036
rect 20536 8984 20588 9036
rect 14280 8848 14332 8900
rect 15476 8848 15528 8900
rect 16212 8848 16264 8900
rect 17868 8916 17920 8968
rect 20260 8916 20312 8968
rect 22560 8984 22612 9036
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 17316 8848 17368 8900
rect 18328 8848 18380 8900
rect 18512 8848 18564 8900
rect 20076 8848 20128 8900
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 10692 8780 10744 8832
rect 12256 8780 12308 8832
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 15752 8780 15804 8832
rect 16856 8780 16908 8832
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 17960 8780 18012 8832
rect 19156 8780 19208 8832
rect 20444 8780 20496 8832
rect 21272 8891 21324 8900
rect 21272 8857 21281 8891
rect 21281 8857 21315 8891
rect 21315 8857 21324 8891
rect 22284 8916 22336 8968
rect 23572 8984 23624 9036
rect 23848 9061 23857 9095
rect 23857 9061 23891 9095
rect 23891 9061 23900 9095
rect 23848 9052 23900 9061
rect 24768 9052 24820 9104
rect 27620 9120 27672 9172
rect 28540 9120 28592 9172
rect 25688 9052 25740 9104
rect 25872 9027 25924 9036
rect 25872 8993 25881 9027
rect 25881 8993 25915 9027
rect 25915 8993 25924 9027
rect 25872 8984 25924 8993
rect 26148 9027 26200 9036
rect 26148 8993 26157 9027
rect 26157 8993 26191 9027
rect 26191 8993 26200 9027
rect 26148 8984 26200 8993
rect 29092 9120 29144 9172
rect 26424 9027 26476 9036
rect 26424 8993 26433 9027
rect 26433 8993 26467 9027
rect 26467 8993 26476 9027
rect 26424 8984 26476 8993
rect 26516 8984 26568 9036
rect 27528 9027 27580 9036
rect 27528 8993 27537 9027
rect 27537 8993 27571 9027
rect 27571 8993 27580 9027
rect 27528 8984 27580 8993
rect 27896 9027 27948 9036
rect 27896 8993 27905 9027
rect 27905 8993 27939 9027
rect 27939 8993 27948 9027
rect 27896 8984 27948 8993
rect 29368 8984 29420 9036
rect 30380 8984 30432 9036
rect 21272 8848 21324 8857
rect 21640 8780 21692 8832
rect 21824 8823 21876 8832
rect 21824 8789 21833 8823
rect 21833 8789 21867 8823
rect 21867 8789 21876 8823
rect 21824 8780 21876 8789
rect 22468 8848 22520 8900
rect 23388 8916 23440 8968
rect 25044 8916 25096 8968
rect 26056 8959 26108 8968
rect 26056 8925 26065 8959
rect 26065 8925 26099 8959
rect 26099 8925 26108 8959
rect 26056 8916 26108 8925
rect 27436 8916 27488 8968
rect 23572 8848 23624 8900
rect 22376 8780 22428 8832
rect 23204 8780 23256 8832
rect 23480 8780 23532 8832
rect 23940 8780 23992 8832
rect 25136 8780 25188 8832
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 26424 8848 26476 8900
rect 26700 8848 26752 8900
rect 27068 8848 27120 8900
rect 29368 8848 29420 8900
rect 29092 8780 29144 8832
rect 30840 8823 30892 8832
rect 30840 8789 30849 8823
rect 30849 8789 30883 8823
rect 30883 8789 30892 8823
rect 30840 8780 30892 8789
rect 6102 8678 6154 8730
rect 6166 8678 6218 8730
rect 6230 8678 6282 8730
rect 6294 8678 6346 8730
rect 6358 8678 6410 8730
rect 16405 8678 16457 8730
rect 16469 8678 16521 8730
rect 16533 8678 16585 8730
rect 16597 8678 16649 8730
rect 16661 8678 16713 8730
rect 26709 8678 26761 8730
rect 26773 8678 26825 8730
rect 26837 8678 26889 8730
rect 26901 8678 26953 8730
rect 26965 8678 27017 8730
rect 5816 8576 5868 8628
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 10140 8576 10192 8628
rect 2136 8508 2188 8560
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 2688 8440 2740 8492
rect 5080 8508 5132 8560
rect 6828 8508 6880 8560
rect 10232 8508 10284 8560
rect 2228 8415 2280 8424
rect 1584 8304 1636 8356
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 2780 8372 2832 8424
rect 3792 8372 3844 8424
rect 3240 8304 3292 8356
rect 10968 8440 11020 8492
rect 4252 8415 4304 8424
rect 4252 8381 4286 8415
rect 4286 8381 4304 8415
rect 4252 8372 4304 8381
rect 5908 8372 5960 8424
rect 7104 8372 7156 8424
rect 7748 8372 7800 8424
rect 10876 8372 10928 8424
rect 11060 8415 11112 8424
rect 11060 8381 11069 8415
rect 11069 8381 11103 8415
rect 11103 8381 11112 8415
rect 11060 8372 11112 8381
rect 11152 8372 11204 8424
rect 12624 8576 12676 8628
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 14096 8619 14148 8628
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 14832 8576 14884 8628
rect 15568 8576 15620 8628
rect 18788 8576 18840 8628
rect 19524 8576 19576 8628
rect 20996 8576 21048 8628
rect 12072 8440 12124 8492
rect 13084 8508 13136 8560
rect 16948 8508 17000 8560
rect 17132 8508 17184 8560
rect 17776 8508 17828 8560
rect 18236 8508 18288 8560
rect 19340 8508 19392 8560
rect 12256 8415 12308 8424
rect 5356 8304 5408 8356
rect 1400 8236 1452 8288
rect 2228 8236 2280 8288
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 6000 8236 6052 8288
rect 9588 8304 9640 8356
rect 10692 8304 10744 8356
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 13636 8440 13688 8492
rect 13176 8372 13228 8424
rect 13544 8372 13596 8424
rect 18328 8440 18380 8492
rect 19156 8440 19208 8492
rect 21640 8576 21692 8628
rect 23572 8576 23624 8628
rect 24768 8619 24820 8628
rect 24768 8585 24777 8619
rect 24777 8585 24811 8619
rect 24811 8585 24820 8619
rect 24768 8576 24820 8585
rect 27344 8619 27396 8628
rect 27344 8585 27353 8619
rect 27353 8585 27387 8619
rect 27387 8585 27396 8619
rect 27344 8576 27396 8585
rect 28080 8576 28132 8628
rect 29460 8576 29512 8628
rect 21456 8508 21508 8560
rect 21916 8508 21968 8560
rect 23388 8508 23440 8560
rect 24952 8508 25004 8560
rect 25872 8508 25924 8560
rect 28172 8508 28224 8560
rect 15752 8372 15804 8424
rect 16212 8372 16264 8424
rect 17776 8415 17828 8424
rect 14372 8304 14424 8356
rect 14924 8304 14976 8356
rect 17040 8304 17092 8356
rect 17316 8347 17368 8356
rect 17316 8313 17325 8347
rect 17325 8313 17359 8347
rect 17359 8313 17368 8347
rect 17316 8304 17368 8313
rect 17776 8381 17785 8415
rect 17785 8381 17819 8415
rect 17819 8381 17828 8415
rect 17776 8372 17828 8381
rect 17960 8415 18012 8424
rect 17960 8381 17969 8415
rect 17969 8381 18003 8415
rect 18003 8381 18012 8415
rect 17960 8372 18012 8381
rect 18052 8304 18104 8356
rect 21824 8372 21876 8424
rect 26700 8440 26752 8492
rect 22376 8415 22428 8424
rect 11704 8236 11756 8288
rect 16948 8279 17000 8288
rect 16948 8245 16957 8279
rect 16957 8245 16991 8279
rect 16991 8245 17000 8279
rect 16948 8236 17000 8245
rect 17960 8236 18012 8288
rect 18144 8236 18196 8288
rect 18512 8236 18564 8288
rect 19248 8236 19300 8288
rect 21364 8304 21416 8356
rect 22100 8304 22152 8356
rect 22376 8381 22385 8415
rect 22385 8381 22419 8415
rect 22419 8381 22428 8415
rect 22376 8372 22428 8381
rect 23940 8372 23992 8424
rect 25964 8415 26016 8424
rect 25964 8381 25973 8415
rect 25973 8381 26007 8415
rect 26007 8381 26016 8415
rect 25964 8372 26016 8381
rect 26424 8372 26476 8424
rect 26516 8372 26568 8424
rect 22652 8347 22704 8356
rect 22652 8313 22686 8347
rect 22686 8313 22704 8347
rect 22652 8304 22704 8313
rect 24768 8304 24820 8356
rect 26332 8304 26384 8356
rect 27068 8372 27120 8424
rect 28908 8440 28960 8492
rect 30932 8440 30984 8492
rect 27528 8372 27580 8424
rect 27436 8304 27488 8356
rect 20720 8236 20772 8288
rect 21088 8236 21140 8288
rect 21272 8236 21324 8288
rect 30380 8304 30432 8356
rect 11253 8134 11305 8186
rect 11317 8134 11369 8186
rect 11381 8134 11433 8186
rect 11445 8134 11497 8186
rect 11509 8134 11561 8186
rect 21557 8134 21609 8186
rect 21621 8134 21673 8186
rect 21685 8134 21737 8186
rect 21749 8134 21801 8186
rect 21813 8134 21865 8186
rect 2412 8032 2464 8084
rect 1676 7964 1728 8016
rect 9588 8075 9640 8084
rect 6736 7964 6788 8016
rect 2228 7942 2280 7951
rect 2228 7908 2237 7942
rect 2237 7908 2271 7942
rect 2271 7908 2280 7942
rect 2228 7899 2280 7908
rect 2688 7896 2740 7948
rect 3240 7939 3292 7948
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 2964 7828 3016 7880
rect 3148 7828 3200 7880
rect 4804 7896 4856 7948
rect 5816 7896 5868 7948
rect 6828 7896 6880 7948
rect 8392 7939 8444 7948
rect 3516 7871 3568 7880
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 4712 7828 4764 7880
rect 4988 7828 5040 7880
rect 5540 7828 5592 7880
rect 5908 7828 5960 7880
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 8852 7939 8904 7948
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 9128 7964 9180 8016
rect 9312 7964 9364 8016
rect 9588 8041 9597 8075
rect 9597 8041 9631 8075
rect 9631 8041 9640 8075
rect 9588 8032 9640 8041
rect 11060 8032 11112 8084
rect 11704 8032 11756 8084
rect 10048 7896 10100 7948
rect 9312 7828 9364 7880
rect 2688 7760 2740 7812
rect 5356 7760 5408 7812
rect 1676 7692 1728 7744
rect 1952 7692 2004 7744
rect 2780 7692 2832 7744
rect 3976 7692 4028 7744
rect 6552 7760 6604 7812
rect 6644 7760 6696 7812
rect 8300 7760 8352 7812
rect 10324 7828 10376 7880
rect 11612 7896 11664 7948
rect 12256 7964 12308 8016
rect 13452 7964 13504 8016
rect 13636 7964 13688 8016
rect 12348 7896 12400 7948
rect 12532 7896 12584 7948
rect 13728 7939 13780 7948
rect 13728 7905 13737 7939
rect 13737 7905 13771 7939
rect 13771 7905 13780 7939
rect 13728 7896 13780 7905
rect 15016 7896 15068 7948
rect 13176 7828 13228 7880
rect 15752 7828 15804 7880
rect 13912 7760 13964 7812
rect 5540 7692 5592 7744
rect 6920 7692 6972 7744
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 10232 7735 10284 7744
rect 10232 7701 10241 7735
rect 10241 7701 10275 7735
rect 10275 7701 10284 7735
rect 10232 7692 10284 7701
rect 10600 7692 10652 7744
rect 10784 7692 10836 7744
rect 12716 7692 12768 7744
rect 13820 7692 13872 7744
rect 16120 7692 16172 7744
rect 17592 7964 17644 8016
rect 16764 7896 16816 7948
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 16672 7760 16724 7812
rect 17224 7760 17276 7812
rect 18144 7964 18196 8016
rect 19524 7964 19576 8016
rect 21272 7964 21324 8016
rect 22652 8032 22704 8084
rect 24492 8032 24544 8084
rect 25964 8032 26016 8084
rect 23480 8007 23532 8016
rect 19708 7896 19760 7948
rect 18880 7828 18932 7880
rect 19156 7871 19208 7880
rect 19156 7837 19165 7871
rect 19165 7837 19199 7871
rect 19199 7837 19208 7871
rect 19156 7828 19208 7837
rect 20352 7828 20404 7880
rect 22100 7896 22152 7948
rect 22284 7871 22336 7880
rect 18512 7760 18564 7812
rect 20536 7803 20588 7812
rect 20536 7769 20545 7803
rect 20545 7769 20579 7803
rect 20579 7769 20588 7803
rect 20536 7760 20588 7769
rect 21272 7760 21324 7812
rect 22008 7760 22060 7812
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 22468 7896 22520 7948
rect 23480 7973 23514 8007
rect 23514 7973 23532 8007
rect 23480 7964 23532 7973
rect 25504 7964 25556 8016
rect 22836 7828 22888 7880
rect 22652 7760 22704 7812
rect 18420 7692 18472 7744
rect 19800 7692 19852 7744
rect 22928 7692 22980 7744
rect 24676 7896 24728 7948
rect 25596 7939 25648 7948
rect 25596 7905 25605 7939
rect 25605 7905 25639 7939
rect 25639 7905 25648 7939
rect 25596 7896 25648 7905
rect 26516 7896 26568 7948
rect 27896 8032 27948 8084
rect 28356 8032 28408 8084
rect 30748 8032 30800 8084
rect 27436 7964 27488 8016
rect 29368 8007 29420 8016
rect 29368 7973 29386 8007
rect 29386 7973 29420 8007
rect 29368 7964 29420 7973
rect 27620 7939 27672 7948
rect 27620 7905 27629 7939
rect 27629 7905 27663 7939
rect 27663 7905 27672 7939
rect 27620 7896 27672 7905
rect 27160 7828 27212 7880
rect 23940 7692 23992 7744
rect 24124 7692 24176 7744
rect 25044 7692 25096 7744
rect 26332 7692 26384 7744
rect 27804 7735 27856 7744
rect 27804 7701 27813 7735
rect 27813 7701 27847 7735
rect 27847 7701 27856 7735
rect 27804 7692 27856 7701
rect 29000 7692 29052 7744
rect 6102 7590 6154 7642
rect 6166 7590 6218 7642
rect 6230 7590 6282 7642
rect 6294 7590 6346 7642
rect 6358 7590 6410 7642
rect 16405 7590 16457 7642
rect 16469 7590 16521 7642
rect 16533 7590 16585 7642
rect 16597 7590 16649 7642
rect 16661 7590 16713 7642
rect 26709 7590 26761 7642
rect 26773 7590 26825 7642
rect 26837 7590 26889 7642
rect 26901 7590 26953 7642
rect 26965 7590 27017 7642
rect 3516 7488 3568 7540
rect 3976 7531 4028 7540
rect 3976 7497 3985 7531
rect 3985 7497 4019 7531
rect 4019 7497 4028 7531
rect 3976 7488 4028 7497
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 5448 7488 5500 7540
rect 3148 7463 3200 7472
rect 3148 7429 3157 7463
rect 3157 7429 3191 7463
rect 3191 7429 3200 7463
rect 3148 7420 3200 7429
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2320 7352 2372 7404
rect 3056 7352 3108 7404
rect 6000 7420 6052 7472
rect 6552 7488 6604 7540
rect 7288 7488 7340 7540
rect 8944 7531 8996 7540
rect 8944 7497 8953 7531
rect 8953 7497 8987 7531
rect 8987 7497 8996 7531
rect 8944 7488 8996 7497
rect 10232 7488 10284 7540
rect 10784 7488 10836 7540
rect 13084 7488 13136 7540
rect 13728 7488 13780 7540
rect 6644 7420 6696 7472
rect 8852 7420 8904 7472
rect 9588 7420 9640 7472
rect 5356 7395 5408 7404
rect 1400 7284 1452 7336
rect 2412 7284 2464 7336
rect 2688 7284 2740 7336
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 3516 7284 3568 7336
rect 5080 7284 5132 7336
rect 2780 7216 2832 7268
rect 3976 7259 4028 7268
rect 1676 7148 1728 7200
rect 3976 7225 4003 7259
rect 4003 7225 4028 7259
rect 3976 7216 4028 7225
rect 4252 7216 4304 7268
rect 8392 7352 8444 7404
rect 5724 7284 5776 7336
rect 6092 7284 6144 7336
rect 6644 7259 6696 7268
rect 6644 7225 6653 7259
rect 6653 7225 6687 7259
rect 6687 7225 6696 7259
rect 6644 7216 6696 7225
rect 6920 7284 6972 7336
rect 7012 7284 7064 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 9220 7216 9272 7268
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 14004 7420 14056 7472
rect 14372 7488 14424 7540
rect 14924 7531 14976 7540
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 15108 7488 15160 7540
rect 16764 7531 16816 7540
rect 16764 7497 16773 7531
rect 16773 7497 16807 7531
rect 16807 7497 16816 7531
rect 16764 7488 16816 7497
rect 17132 7488 17184 7540
rect 10692 7352 10744 7404
rect 16856 7420 16908 7472
rect 17776 7463 17828 7472
rect 17776 7429 17785 7463
rect 17785 7429 17819 7463
rect 17819 7429 17828 7463
rect 18236 7488 18288 7540
rect 19892 7488 19944 7540
rect 22100 7488 22152 7540
rect 23112 7488 23164 7540
rect 24768 7531 24820 7540
rect 24768 7497 24777 7531
rect 24777 7497 24811 7531
rect 24811 7497 24820 7531
rect 24768 7488 24820 7497
rect 17776 7420 17828 7429
rect 9496 7284 9548 7293
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11060 7284 11112 7336
rect 9956 7216 10008 7268
rect 11796 7284 11848 7336
rect 12256 7284 12308 7336
rect 12532 7284 12584 7336
rect 13084 7284 13136 7336
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 16396 7352 16448 7404
rect 14832 7284 14884 7336
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 15660 7327 15712 7336
rect 13912 7216 13964 7268
rect 15660 7293 15669 7327
rect 15669 7293 15703 7327
rect 15703 7293 15712 7327
rect 15660 7284 15712 7293
rect 16948 7352 17000 7404
rect 17132 7352 17184 7404
rect 16764 7284 16816 7336
rect 18420 7420 18472 7472
rect 22560 7420 22612 7472
rect 25504 7463 25556 7472
rect 25504 7429 25513 7463
rect 25513 7429 25547 7463
rect 25547 7429 25556 7463
rect 25504 7420 25556 7429
rect 29276 7488 29328 7540
rect 30012 7488 30064 7540
rect 30840 7420 30892 7472
rect 17408 7284 17460 7336
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 18696 7352 18748 7404
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 24492 7352 24544 7404
rect 26332 7395 26384 7404
rect 18512 7284 18564 7336
rect 19432 7327 19484 7336
rect 16948 7216 17000 7268
rect 19432 7293 19441 7327
rect 19441 7293 19475 7327
rect 19475 7293 19484 7327
rect 19432 7284 19484 7293
rect 4896 7148 4948 7200
rect 5172 7148 5224 7200
rect 5724 7148 5776 7200
rect 7104 7148 7156 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 11704 7148 11756 7200
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 13636 7148 13688 7200
rect 15108 7148 15160 7200
rect 16120 7148 16172 7200
rect 17408 7148 17460 7200
rect 17500 7148 17552 7200
rect 20444 7284 20496 7336
rect 22376 7284 22428 7336
rect 20168 7216 20220 7268
rect 20812 7216 20864 7268
rect 22008 7216 22060 7268
rect 24860 7284 24912 7336
rect 26332 7361 26341 7395
rect 26341 7361 26375 7395
rect 26375 7361 26384 7395
rect 26332 7352 26384 7361
rect 26516 7352 26568 7404
rect 25688 7327 25740 7336
rect 25688 7293 25697 7327
rect 25697 7293 25731 7327
rect 25731 7293 25740 7327
rect 25688 7284 25740 7293
rect 25964 7284 26016 7336
rect 27068 7284 27120 7336
rect 27804 7284 27856 7336
rect 29000 7327 29052 7336
rect 29000 7293 29009 7327
rect 29009 7293 29043 7327
rect 29043 7293 29052 7327
rect 29000 7284 29052 7293
rect 31116 7327 31168 7336
rect 31116 7293 31125 7327
rect 31125 7293 31159 7327
rect 31159 7293 31168 7327
rect 31116 7284 31168 7293
rect 25780 7216 25832 7268
rect 23756 7191 23808 7200
rect 23756 7157 23765 7191
rect 23765 7157 23799 7191
rect 23799 7157 23808 7191
rect 23756 7148 23808 7157
rect 25136 7148 25188 7200
rect 27620 7191 27672 7200
rect 27620 7157 27629 7191
rect 27629 7157 27663 7191
rect 27663 7157 27672 7191
rect 27620 7148 27672 7157
rect 11253 7046 11305 7098
rect 11317 7046 11369 7098
rect 11381 7046 11433 7098
rect 11445 7046 11497 7098
rect 11509 7046 11561 7098
rect 21557 7046 21609 7098
rect 21621 7046 21673 7098
rect 21685 7046 21737 7098
rect 21749 7046 21801 7098
rect 21813 7046 21865 7098
rect 1584 6808 1636 6860
rect 1952 6944 2004 6996
rect 3516 6987 3568 6996
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 5356 6944 5408 6996
rect 2412 6876 2464 6928
rect 3976 6876 4028 6928
rect 4068 6876 4120 6928
rect 5724 6944 5776 6996
rect 5816 6944 5868 6996
rect 8024 6944 8076 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 15660 6944 15712 6996
rect 17224 6987 17276 6996
rect 17224 6953 17233 6987
rect 17233 6953 17267 6987
rect 17267 6953 17276 6987
rect 17224 6944 17276 6953
rect 18144 6944 18196 6996
rect 22008 6987 22060 6996
rect 22008 6953 22017 6987
rect 22017 6953 22051 6987
rect 22051 6953 22060 6987
rect 22008 6944 22060 6953
rect 22928 6944 22980 6996
rect 28356 6944 28408 6996
rect 31116 6944 31168 6996
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 2688 6808 2740 6860
rect 2964 6808 3016 6860
rect 3332 6808 3384 6860
rect 3608 6808 3660 6860
rect 4160 6808 4212 6860
rect 2504 6740 2556 6792
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3148 6740 3200 6792
rect 5264 6808 5316 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 5448 6808 5500 6817
rect 5172 6740 5224 6792
rect 2964 6672 3016 6724
rect 4436 6672 4488 6724
rect 5724 6808 5776 6860
rect 10692 6876 10744 6928
rect 8392 6808 8444 6860
rect 9864 6808 9916 6860
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 11704 6851 11756 6860
rect 11704 6817 11713 6851
rect 11713 6817 11747 6851
rect 11747 6817 11756 6851
rect 11704 6808 11756 6817
rect 11796 6808 11848 6860
rect 12716 6876 12768 6928
rect 14740 6876 14792 6928
rect 12256 6851 12308 6860
rect 12256 6817 12265 6851
rect 12265 6817 12299 6851
rect 12299 6817 12308 6851
rect 12256 6808 12308 6817
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 14004 6851 14056 6860
rect 12440 6808 12492 6817
rect 14004 6817 14022 6851
rect 14022 6817 14056 6851
rect 14004 6808 14056 6817
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 15108 6808 15160 6860
rect 15384 6851 15436 6860
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 15660 6808 15712 6860
rect 15936 6876 15988 6928
rect 23756 6876 23808 6928
rect 24860 6876 24912 6928
rect 15844 6808 15896 6860
rect 16856 6851 16908 6860
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 17040 6851 17092 6860
rect 17040 6817 17049 6851
rect 17049 6817 17083 6851
rect 17083 6817 17092 6851
rect 17040 6808 17092 6817
rect 11060 6740 11112 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 16120 6740 16172 6792
rect 17868 6740 17920 6792
rect 18144 6808 18196 6860
rect 19340 6851 19392 6860
rect 19340 6817 19349 6851
rect 19349 6817 19383 6851
rect 19383 6817 19392 6851
rect 19340 6808 19392 6817
rect 19708 6808 19760 6860
rect 18512 6740 18564 6792
rect 5816 6672 5868 6724
rect 6092 6672 6144 6724
rect 7748 6672 7800 6724
rect 16304 6672 16356 6724
rect 17592 6672 17644 6724
rect 22100 6808 22152 6860
rect 22284 6808 22336 6860
rect 22652 6808 22704 6860
rect 23480 6808 23532 6860
rect 24952 6808 25004 6860
rect 25136 6851 25188 6860
rect 25136 6817 25145 6851
rect 25145 6817 25179 6851
rect 25179 6817 25188 6851
rect 25136 6808 25188 6817
rect 2504 6604 2556 6656
rect 6000 6604 6052 6656
rect 9680 6604 9732 6656
rect 10140 6604 10192 6656
rect 12532 6604 12584 6656
rect 13544 6604 13596 6656
rect 15568 6604 15620 6656
rect 21088 6672 21140 6724
rect 23848 6740 23900 6792
rect 24860 6740 24912 6792
rect 20720 6647 20772 6656
rect 20720 6613 20729 6647
rect 20729 6613 20763 6647
rect 20763 6613 20772 6647
rect 20720 6604 20772 6613
rect 22468 6672 22520 6724
rect 22928 6672 22980 6724
rect 25596 6851 25648 6860
rect 25596 6817 25605 6851
rect 25605 6817 25639 6851
rect 25639 6817 25648 6851
rect 25596 6808 25648 6817
rect 25780 6851 25832 6860
rect 25780 6817 25789 6851
rect 25789 6817 25823 6851
rect 25823 6817 25832 6851
rect 25780 6808 25832 6817
rect 26516 6808 26568 6860
rect 27620 6808 27672 6860
rect 28448 6808 28500 6860
rect 29092 6808 29144 6860
rect 29276 6808 29328 6860
rect 31300 6808 31352 6860
rect 25504 6783 25556 6792
rect 25504 6749 25513 6783
rect 25513 6749 25547 6783
rect 25547 6749 25556 6783
rect 25504 6740 25556 6749
rect 27436 6783 27488 6792
rect 27436 6749 27445 6783
rect 27445 6749 27479 6783
rect 27479 6749 27488 6783
rect 27436 6740 27488 6749
rect 27528 6783 27580 6792
rect 27528 6749 27537 6783
rect 27537 6749 27571 6783
rect 27571 6749 27580 6783
rect 27528 6740 27580 6749
rect 28724 6740 28776 6792
rect 30748 6740 30800 6792
rect 25412 6715 25464 6724
rect 25412 6681 25421 6715
rect 25421 6681 25455 6715
rect 25455 6681 25464 6715
rect 25412 6672 25464 6681
rect 23664 6604 23716 6656
rect 24400 6604 24452 6656
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 27896 6647 27948 6656
rect 27896 6613 27905 6647
rect 27905 6613 27939 6647
rect 27939 6613 27948 6647
rect 27896 6604 27948 6613
rect 28356 6647 28408 6656
rect 28356 6613 28365 6647
rect 28365 6613 28399 6647
rect 28399 6613 28408 6647
rect 28356 6604 28408 6613
rect 28632 6604 28684 6656
rect 6102 6502 6154 6554
rect 6166 6502 6218 6554
rect 6230 6502 6282 6554
rect 6294 6502 6346 6554
rect 6358 6502 6410 6554
rect 16405 6502 16457 6554
rect 16469 6502 16521 6554
rect 16533 6502 16585 6554
rect 16597 6502 16649 6554
rect 16661 6502 16713 6554
rect 26709 6502 26761 6554
rect 26773 6502 26825 6554
rect 26837 6502 26889 6554
rect 26901 6502 26953 6554
rect 26965 6502 27017 6554
rect 2688 6400 2740 6452
rect 3056 6400 3108 6452
rect 4804 6400 4856 6452
rect 5080 6400 5132 6452
rect 1952 6332 2004 6384
rect 4068 6332 4120 6384
rect 5724 6264 5776 6316
rect 9220 6400 9272 6452
rect 10416 6400 10468 6452
rect 11612 6400 11664 6452
rect 11888 6400 11940 6452
rect 12256 6400 12308 6452
rect 14004 6400 14056 6452
rect 14556 6400 14608 6452
rect 5908 6375 5960 6384
rect 5908 6341 5917 6375
rect 5917 6341 5951 6375
rect 5951 6341 5960 6375
rect 5908 6332 5960 6341
rect 7564 6264 7616 6316
rect 10232 6332 10284 6384
rect 8668 6264 8720 6316
rect 4436 6196 4488 6248
rect 5080 6196 5132 6248
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 6000 6196 6052 6248
rect 7196 6196 7248 6248
rect 8852 6196 8904 6248
rect 10600 6264 10652 6316
rect 1676 6128 1728 6180
rect 2964 6128 3016 6180
rect 5632 6128 5684 6180
rect 8760 6128 8812 6180
rect 9220 6205 9223 6226
rect 9223 6205 9257 6226
rect 9257 6205 9272 6226
rect 9220 6174 9272 6205
rect 9496 6239 9548 6248
rect 9496 6205 9516 6239
rect 9516 6205 9548 6239
rect 9496 6196 9548 6205
rect 9864 6196 9916 6248
rect 10140 6239 10192 6248
rect 10140 6205 10149 6239
rect 10149 6205 10183 6239
rect 10183 6205 10192 6239
rect 10140 6196 10192 6205
rect 9404 6128 9456 6180
rect 10048 6128 10100 6180
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 12348 6264 12400 6316
rect 10416 6196 10468 6205
rect 12716 6239 12768 6248
rect 12716 6205 12725 6239
rect 12725 6205 12759 6239
rect 12759 6205 12768 6239
rect 12716 6196 12768 6205
rect 12808 6196 12860 6248
rect 13544 6196 13596 6248
rect 14372 6196 14424 6248
rect 16120 6400 16172 6452
rect 16856 6400 16908 6452
rect 17040 6400 17092 6452
rect 17316 6332 17368 6384
rect 12624 6128 12676 6180
rect 13452 6128 13504 6180
rect 16856 6196 16908 6248
rect 17592 6400 17644 6452
rect 21272 6400 21324 6452
rect 21916 6400 21968 6452
rect 23112 6400 23164 6452
rect 27068 6443 27120 6452
rect 27068 6409 27077 6443
rect 27077 6409 27111 6443
rect 27111 6409 27120 6443
rect 27068 6400 27120 6409
rect 20260 6332 20312 6384
rect 23664 6332 23716 6384
rect 28356 6400 28408 6452
rect 28724 6400 28776 6452
rect 29276 6400 29328 6452
rect 30104 6443 30156 6452
rect 30104 6409 30113 6443
rect 30113 6409 30147 6443
rect 30147 6409 30156 6443
rect 30104 6400 30156 6409
rect 31024 6400 31076 6452
rect 31576 6400 31628 6452
rect 27344 6332 27396 6384
rect 27528 6332 27580 6384
rect 19892 6307 19944 6316
rect 19892 6273 19901 6307
rect 19901 6273 19935 6307
rect 19935 6273 19944 6307
rect 19892 6264 19944 6273
rect 20904 6264 20956 6316
rect 21916 6264 21968 6316
rect 22284 6264 22336 6316
rect 22836 6307 22888 6316
rect 22836 6273 22845 6307
rect 22845 6273 22879 6307
rect 22879 6273 22888 6307
rect 22836 6264 22888 6273
rect 23756 6307 23808 6316
rect 23756 6273 23765 6307
rect 23765 6273 23799 6307
rect 23799 6273 23808 6307
rect 23756 6264 23808 6273
rect 26424 6264 26476 6316
rect 27160 6264 27212 6316
rect 19248 6196 19300 6248
rect 16764 6128 16816 6180
rect 17776 6128 17828 6180
rect 19064 6128 19116 6180
rect 19800 6239 19852 6248
rect 19800 6205 19809 6239
rect 19809 6205 19843 6239
rect 19843 6205 19852 6239
rect 19800 6196 19852 6205
rect 21088 6196 21140 6248
rect 22008 6196 22060 6248
rect 22560 6239 22612 6248
rect 22560 6205 22569 6239
rect 22569 6205 22603 6239
rect 22603 6205 22612 6239
rect 22560 6196 22612 6205
rect 22928 6239 22980 6248
rect 4528 6060 4580 6112
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 8024 6060 8076 6112
rect 15292 6103 15344 6112
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 16672 6060 16724 6112
rect 20904 6128 20956 6180
rect 22468 6128 22520 6180
rect 22928 6205 22937 6239
rect 22937 6205 22971 6239
rect 22971 6205 22980 6239
rect 22928 6196 22980 6205
rect 23848 6196 23900 6248
rect 24584 6196 24636 6248
rect 23480 6128 23532 6180
rect 24768 6128 24820 6180
rect 26148 6128 26200 6180
rect 26332 6239 26384 6248
rect 26332 6205 26341 6239
rect 26341 6205 26375 6239
rect 26375 6205 26384 6239
rect 26608 6239 26660 6248
rect 26332 6196 26384 6205
rect 26608 6205 26617 6239
rect 26617 6205 26651 6239
rect 26651 6205 26660 6239
rect 26608 6196 26660 6205
rect 27528 6196 27580 6248
rect 27896 6239 27948 6248
rect 27896 6205 27930 6239
rect 27930 6205 27948 6239
rect 27896 6196 27948 6205
rect 28356 6128 28408 6180
rect 20168 6060 20220 6112
rect 23296 6103 23348 6112
rect 23296 6069 23305 6103
rect 23305 6069 23339 6103
rect 23339 6069 23348 6103
rect 23296 6060 23348 6069
rect 26424 6060 26476 6112
rect 28448 6060 28500 6112
rect 11253 5958 11305 6010
rect 11317 5958 11369 6010
rect 11381 5958 11433 6010
rect 11445 5958 11497 6010
rect 11509 5958 11561 6010
rect 21557 5958 21609 6010
rect 21621 5958 21673 6010
rect 21685 5958 21737 6010
rect 21749 5958 21801 6010
rect 21813 5958 21865 6010
rect 2412 5856 2464 5908
rect 2780 5856 2832 5908
rect 3240 5856 3292 5908
rect 5172 5899 5224 5908
rect 2228 5831 2280 5840
rect 2228 5797 2237 5831
rect 2237 5797 2271 5831
rect 2271 5797 2280 5831
rect 2228 5788 2280 5797
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 5448 5856 5500 5908
rect 7196 5899 7248 5908
rect 1584 5720 1636 5772
rect 2504 5720 2556 5772
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 4804 5788 4856 5840
rect 2136 5584 2188 5636
rect 3148 5584 3200 5636
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 4988 5720 5040 5772
rect 5356 5720 5408 5772
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 8760 5856 8812 5908
rect 9220 5856 9272 5908
rect 6736 5788 6788 5840
rect 8024 5831 8076 5840
rect 8024 5797 8058 5831
rect 8058 5797 8076 5831
rect 8024 5788 8076 5797
rect 8668 5788 8720 5840
rect 9864 5788 9916 5840
rect 12072 5856 12124 5908
rect 16672 5856 16724 5908
rect 16856 5856 16908 5908
rect 17408 5856 17460 5908
rect 17868 5856 17920 5908
rect 19064 5899 19116 5908
rect 19064 5865 19073 5899
rect 19073 5865 19107 5899
rect 19107 5865 19116 5899
rect 19064 5856 19116 5865
rect 21916 5856 21968 5908
rect 23848 5856 23900 5908
rect 24492 5899 24544 5908
rect 24492 5865 24501 5899
rect 24501 5865 24535 5899
rect 24535 5865 24544 5899
rect 24492 5856 24544 5865
rect 25412 5856 25464 5908
rect 7104 5763 7156 5772
rect 4620 5652 4672 5704
rect 5356 5584 5408 5636
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 6000 5652 6052 5704
rect 6920 5652 6972 5704
rect 9128 5652 9180 5704
rect 9956 5720 10008 5772
rect 10048 5652 10100 5704
rect 4068 5516 4120 5568
rect 5172 5516 5224 5568
rect 7012 5584 7064 5636
rect 10692 5720 10744 5772
rect 11152 5720 11204 5772
rect 11244 5720 11296 5772
rect 15292 5788 15344 5840
rect 14004 5763 14056 5772
rect 14004 5729 14022 5763
rect 14022 5729 14056 5763
rect 14004 5720 14056 5729
rect 15476 5763 15528 5772
rect 11060 5652 11112 5704
rect 12348 5652 12400 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 15476 5720 15528 5729
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 15844 5720 15896 5772
rect 17316 5720 17368 5772
rect 17776 5763 17828 5772
rect 17776 5729 17785 5763
rect 17785 5729 17819 5763
rect 17819 5729 17828 5763
rect 17776 5720 17828 5729
rect 23296 5788 23348 5840
rect 24400 5788 24452 5840
rect 19616 5720 19668 5772
rect 21088 5763 21140 5772
rect 21088 5729 21097 5763
rect 21097 5729 21131 5763
rect 21131 5729 21140 5763
rect 21088 5720 21140 5729
rect 23940 5720 23992 5772
rect 24676 5763 24728 5772
rect 24676 5729 24685 5763
rect 24685 5729 24719 5763
rect 24719 5729 24728 5763
rect 24676 5720 24728 5729
rect 24768 5720 24820 5772
rect 25228 5763 25280 5772
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 26516 5856 26568 5908
rect 26608 5856 26660 5908
rect 28356 5899 28408 5908
rect 28356 5865 28365 5899
rect 28365 5865 28399 5899
rect 28399 5865 28408 5899
rect 28356 5856 28408 5865
rect 29276 5856 29328 5908
rect 30564 5899 30616 5908
rect 30564 5865 30573 5899
rect 30573 5865 30607 5899
rect 30607 5865 30616 5899
rect 30564 5856 30616 5865
rect 31116 5899 31168 5908
rect 31116 5865 31125 5899
rect 31125 5865 31159 5899
rect 31159 5865 31168 5899
rect 31116 5856 31168 5865
rect 26056 5763 26108 5772
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 10232 5516 10284 5568
rect 10968 5516 11020 5568
rect 12808 5516 12860 5568
rect 15660 5584 15712 5636
rect 14556 5516 14608 5568
rect 15016 5559 15068 5568
rect 15016 5525 15025 5559
rect 15025 5525 15059 5559
rect 15059 5525 15068 5559
rect 15016 5516 15068 5525
rect 17408 5652 17460 5704
rect 18604 5652 18656 5704
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 21456 5652 21508 5704
rect 22284 5652 22336 5704
rect 26056 5729 26065 5763
rect 26065 5729 26099 5763
rect 26099 5729 26108 5763
rect 26056 5720 26108 5729
rect 26157 5695 26209 5704
rect 26157 5661 26163 5695
rect 26163 5661 26197 5695
rect 26197 5661 26209 5695
rect 26157 5652 26209 5661
rect 26424 5763 26476 5772
rect 26424 5729 26433 5763
rect 26433 5729 26467 5763
rect 26467 5729 26476 5763
rect 26424 5720 26476 5729
rect 26608 5720 26660 5772
rect 27620 5763 27672 5772
rect 27620 5729 27629 5763
rect 27629 5729 27663 5763
rect 27663 5729 27672 5763
rect 27620 5720 27672 5729
rect 28448 5763 28500 5772
rect 28448 5729 28457 5763
rect 28457 5729 28491 5763
rect 28491 5729 28500 5763
rect 28448 5720 28500 5729
rect 27252 5652 27304 5704
rect 17960 5584 18012 5636
rect 18052 5516 18104 5568
rect 20996 5559 21048 5568
rect 20996 5525 21005 5559
rect 21005 5525 21039 5559
rect 21039 5525 21048 5559
rect 20996 5516 21048 5525
rect 25228 5516 25280 5568
rect 30104 5516 30156 5568
rect 6102 5414 6154 5466
rect 6166 5414 6218 5466
rect 6230 5414 6282 5466
rect 6294 5414 6346 5466
rect 6358 5414 6410 5466
rect 16405 5414 16457 5466
rect 16469 5414 16521 5466
rect 16533 5414 16585 5466
rect 16597 5414 16649 5466
rect 16661 5414 16713 5466
rect 26709 5414 26761 5466
rect 26773 5414 26825 5466
rect 26837 5414 26889 5466
rect 26901 5414 26953 5466
rect 26965 5414 27017 5466
rect 2964 5312 3016 5364
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 9588 5312 9640 5364
rect 11980 5312 12032 5364
rect 17684 5312 17736 5364
rect 18236 5312 18288 5364
rect 18696 5355 18748 5364
rect 18696 5321 18705 5355
rect 18705 5321 18739 5355
rect 18739 5321 18748 5355
rect 18696 5312 18748 5321
rect 10784 5244 10836 5296
rect 11060 5244 11112 5296
rect 11244 5244 11296 5296
rect 7748 5176 7800 5228
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 3792 5151 3844 5160
rect 1676 5108 1728 5117
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 4068 5151 4120 5160
rect 4068 5117 4102 5151
rect 4102 5117 4120 5151
rect 4068 5108 4120 5117
rect 5724 5108 5776 5160
rect 1768 5040 1820 5092
rect 4160 5040 4212 5092
rect 5632 5040 5684 5092
rect 6000 5040 6052 5092
rect 2320 4972 2372 5024
rect 2688 4972 2740 5024
rect 5356 4972 5408 5024
rect 6828 5108 6880 5160
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 9404 5108 9456 5160
rect 10600 5176 10652 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 12716 5244 12768 5296
rect 10968 5176 11020 5185
rect 12348 5176 12400 5228
rect 14372 5244 14424 5296
rect 17132 5244 17184 5296
rect 7104 5040 7156 5092
rect 10692 5108 10744 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 10968 5040 11020 5092
rect 11612 5040 11664 5092
rect 12256 5040 12308 5092
rect 6920 4972 6972 5024
rect 11888 4972 11940 5024
rect 17224 5176 17276 5228
rect 18052 5176 18104 5228
rect 18604 5244 18656 5296
rect 20720 5244 20772 5296
rect 24952 5312 25004 5364
rect 27068 5312 27120 5364
rect 27804 5312 27856 5364
rect 28724 5355 28776 5364
rect 28724 5321 28733 5355
rect 28733 5321 28767 5355
rect 28767 5321 28776 5355
rect 28724 5312 28776 5321
rect 30012 5312 30064 5364
rect 30656 5355 30708 5364
rect 30656 5321 30665 5355
rect 30665 5321 30699 5355
rect 30699 5321 30708 5355
rect 30656 5312 30708 5321
rect 31116 5312 31168 5364
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 14280 5108 14332 5160
rect 15752 5108 15804 5160
rect 15016 5040 15068 5092
rect 13084 4972 13136 5024
rect 14372 4972 14424 5024
rect 15660 4972 15712 5024
rect 17408 5108 17460 5160
rect 17960 5151 18012 5160
rect 17960 5117 17969 5151
rect 17969 5117 18003 5151
rect 18003 5117 18012 5151
rect 17960 5108 18012 5117
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 20996 5176 21048 5228
rect 22376 5176 22428 5228
rect 24584 5244 24636 5296
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 22928 5176 22980 5228
rect 24492 5176 24544 5228
rect 26056 5244 26108 5296
rect 27436 5244 27488 5296
rect 30288 5244 30340 5296
rect 26884 5176 26936 5228
rect 18052 5040 18104 5092
rect 18604 5108 18656 5160
rect 19800 5108 19852 5160
rect 23480 5108 23532 5160
rect 24860 5151 24912 5160
rect 24860 5117 24869 5151
rect 24869 5117 24903 5151
rect 24903 5117 24912 5151
rect 24860 5108 24912 5117
rect 25136 5151 25188 5160
rect 21824 5083 21876 5092
rect 21824 5049 21842 5083
rect 21842 5049 21876 5083
rect 21824 5040 21876 5049
rect 23664 5040 23716 5092
rect 25136 5117 25145 5151
rect 25145 5117 25179 5151
rect 25179 5117 25188 5151
rect 25136 5108 25188 5117
rect 26056 5151 26108 5160
rect 16764 4972 16816 5024
rect 16856 4972 16908 5024
rect 18880 4972 18932 5024
rect 20720 5015 20772 5024
rect 20720 4981 20729 5015
rect 20729 4981 20763 5015
rect 20763 4981 20772 5015
rect 20720 4972 20772 4981
rect 24308 4972 24360 5024
rect 26056 5117 26065 5151
rect 26065 5117 26099 5151
rect 26099 5117 26108 5151
rect 26056 5108 26108 5117
rect 26240 5108 26292 5160
rect 27068 5108 27120 5160
rect 27436 5108 27488 5160
rect 27620 5108 27672 5160
rect 31300 5108 31352 5160
rect 26332 4972 26384 5024
rect 27252 5040 27304 5092
rect 27436 4972 27488 5024
rect 27712 5015 27764 5024
rect 27712 4981 27721 5015
rect 27721 4981 27755 5015
rect 27755 4981 27764 5015
rect 27712 4972 27764 4981
rect 11253 4870 11305 4922
rect 11317 4870 11369 4922
rect 11381 4870 11433 4922
rect 11445 4870 11497 4922
rect 11509 4870 11561 4922
rect 21557 4870 21609 4922
rect 21621 4870 21673 4922
rect 21685 4870 21737 4922
rect 21749 4870 21801 4922
rect 21813 4870 21865 4922
rect 2136 4768 2188 4820
rect 2688 4768 2740 4820
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 3700 4811 3752 4820
rect 3700 4777 3709 4811
rect 3709 4777 3743 4811
rect 3743 4777 3752 4811
rect 3700 4768 3752 4777
rect 4620 4768 4672 4820
rect 7104 4811 7156 4820
rect 3240 4700 3292 4752
rect 3148 4632 3200 4684
rect 3884 4632 3936 4684
rect 4436 4632 4488 4684
rect 4712 4632 4764 4684
rect 5080 4632 5132 4684
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 9128 4768 9180 4820
rect 14004 4768 14056 4820
rect 15568 4768 15620 4820
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 7748 4632 7800 4684
rect 9128 4632 9180 4684
rect 11060 4632 11112 4684
rect 12532 4700 12584 4752
rect 13176 4700 13228 4752
rect 5264 4564 5316 4616
rect 5632 4564 5684 4616
rect 6460 4496 6512 4548
rect 10232 4564 10284 4616
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 12808 4632 12860 4684
rect 13084 4675 13136 4684
rect 12440 4564 12492 4616
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 15200 4700 15252 4752
rect 18604 4700 18656 4752
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 15476 4675 15528 4684
rect 15476 4641 15494 4675
rect 15494 4641 15528 4675
rect 15476 4632 15528 4641
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 17500 4675 17552 4684
rect 17500 4641 17509 4675
rect 17509 4641 17543 4675
rect 17543 4641 17552 4675
rect 17500 4632 17552 4641
rect 19248 4768 19300 4820
rect 19616 4768 19668 4820
rect 21916 4768 21968 4820
rect 23480 4768 23532 4820
rect 26516 4768 26568 4820
rect 27620 4811 27672 4820
rect 19064 4700 19116 4752
rect 18880 4675 18932 4684
rect 18880 4641 18889 4675
rect 18889 4641 18923 4675
rect 18923 4641 18932 4675
rect 18880 4632 18932 4641
rect 20444 4700 20496 4752
rect 22192 4700 22244 4752
rect 12256 4496 12308 4548
rect 12348 4496 12400 4548
rect 16304 4564 16356 4616
rect 17408 4564 17460 4616
rect 19064 4607 19116 4616
rect 19064 4573 19073 4607
rect 19073 4573 19107 4607
rect 19107 4573 19116 4607
rect 19064 4564 19116 4573
rect 20168 4675 20220 4684
rect 20168 4641 20202 4675
rect 20202 4641 20220 4675
rect 20168 4632 20220 4641
rect 20720 4632 20772 4684
rect 23940 4700 23992 4752
rect 22560 4675 22612 4684
rect 22560 4641 22569 4675
rect 22569 4641 22603 4675
rect 22603 4641 22612 4675
rect 22560 4632 22612 4641
rect 24308 4632 24360 4684
rect 26056 4700 26108 4752
rect 26884 4700 26936 4752
rect 24768 4632 24820 4684
rect 25044 4632 25096 4684
rect 26148 4675 26200 4684
rect 26148 4641 26157 4675
rect 26157 4641 26191 4675
rect 26191 4641 26200 4675
rect 26148 4632 26200 4641
rect 27620 4777 27629 4811
rect 27629 4777 27663 4811
rect 27663 4777 27672 4811
rect 27620 4768 27672 4777
rect 30012 4768 30064 4820
rect 30564 4768 30616 4820
rect 31024 4811 31076 4820
rect 31024 4777 31033 4811
rect 31033 4777 31067 4811
rect 31067 4777 31076 4811
rect 31024 4768 31076 4777
rect 27712 4700 27764 4752
rect 30472 4743 30524 4752
rect 30472 4709 30481 4743
rect 30481 4709 30515 4743
rect 30515 4709 30524 4743
rect 30472 4700 30524 4709
rect 31208 4700 31260 4752
rect 29000 4675 29052 4684
rect 19800 4564 19852 4616
rect 22192 4607 22244 4616
rect 17960 4539 18012 4548
rect 17960 4505 17969 4539
rect 17969 4505 18003 4539
rect 18003 4505 18012 4539
rect 17960 4496 18012 4505
rect 22192 4573 22201 4607
rect 22201 4573 22235 4607
rect 22235 4573 22244 4607
rect 22192 4564 22244 4573
rect 22836 4564 22888 4616
rect 25136 4607 25188 4616
rect 25136 4573 25145 4607
rect 25145 4573 25179 4607
rect 25179 4573 25188 4607
rect 25136 4564 25188 4573
rect 25964 4564 26016 4616
rect 29000 4641 29009 4675
rect 29009 4641 29043 4675
rect 29043 4641 29052 4675
rect 29000 4632 29052 4641
rect 5540 4428 5592 4480
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 19892 4428 19944 4480
rect 27988 4496 28040 4548
rect 21088 4428 21140 4480
rect 26424 4428 26476 4480
rect 28356 4428 28408 4480
rect 6102 4326 6154 4378
rect 6166 4326 6218 4378
rect 6230 4326 6282 4378
rect 6294 4326 6346 4378
rect 6358 4326 6410 4378
rect 16405 4326 16457 4378
rect 16469 4326 16521 4378
rect 16533 4326 16585 4378
rect 16597 4326 16649 4378
rect 16661 4326 16713 4378
rect 26709 4326 26761 4378
rect 26773 4326 26825 4378
rect 26837 4326 26889 4378
rect 26901 4326 26953 4378
rect 26965 4326 27017 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 2872 4224 2924 4276
rect 4436 4267 4488 4276
rect 4436 4233 4445 4267
rect 4445 4233 4479 4267
rect 4479 4233 4488 4267
rect 4436 4224 4488 4233
rect 6920 4224 6972 4276
rect 12348 4224 12400 4276
rect 1860 4088 1912 4140
rect 4344 4156 4396 4208
rect 7748 4156 7800 4208
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 9404 4088 9456 4140
rect 10232 4088 10284 4140
rect 5540 4063 5592 4072
rect 5540 4029 5558 4063
rect 5558 4029 5592 4063
rect 5540 4020 5592 4029
rect 7932 4020 7984 4072
rect 8576 4020 8628 4072
rect 9220 4020 9272 4072
rect 4896 3952 4948 4004
rect 10048 4020 10100 4072
rect 10692 4156 10744 4208
rect 12808 4224 12860 4276
rect 13820 4224 13872 4276
rect 15476 4267 15528 4276
rect 15476 4233 15485 4267
rect 15485 4233 15519 4267
rect 15519 4233 15528 4267
rect 15476 4224 15528 4233
rect 12624 4156 12676 4208
rect 14096 4156 14148 4208
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 12256 4063 12308 4072
rect 12256 4029 12265 4063
rect 12265 4029 12299 4063
rect 12299 4029 12308 4063
rect 12256 4020 12308 4029
rect 13636 4088 13688 4140
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 9956 3952 10008 4004
rect 7288 3884 7340 3936
rect 10324 3952 10376 4004
rect 12532 3952 12584 4004
rect 10140 3884 10192 3936
rect 10600 3884 10652 3936
rect 13176 4020 13228 4072
rect 14096 4063 14148 4072
rect 14096 4029 14105 4063
rect 14105 4029 14139 4063
rect 14139 4029 14148 4063
rect 14096 4020 14148 4029
rect 14556 4088 14608 4140
rect 15384 4088 15436 4140
rect 17960 4224 18012 4276
rect 18144 4224 18196 4276
rect 22376 4224 22428 4276
rect 27436 4224 27488 4276
rect 17224 4156 17276 4208
rect 16764 4088 16816 4140
rect 17592 4088 17644 4140
rect 18236 4156 18288 4208
rect 19248 4156 19300 4208
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 18328 4088 18380 4140
rect 24676 4088 24728 4140
rect 27160 4088 27212 4140
rect 27528 4131 27580 4140
rect 14280 3952 14332 4004
rect 15568 4020 15620 4072
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 16304 4020 16356 4072
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 17040 3952 17092 4004
rect 12900 3884 12952 3936
rect 16120 3884 16172 3936
rect 17684 4063 17736 4072
rect 17684 4029 17693 4063
rect 17693 4029 17727 4063
rect 17727 4029 17736 4063
rect 17684 4020 17736 4029
rect 18236 4063 18288 4072
rect 18236 4029 18245 4063
rect 18245 4029 18279 4063
rect 18279 4029 18288 4063
rect 18236 4020 18288 4029
rect 19708 4020 19760 4072
rect 21180 4063 21232 4072
rect 21180 4029 21189 4063
rect 21189 4029 21223 4063
rect 21223 4029 21232 4063
rect 21180 4020 21232 4029
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 24584 4063 24636 4072
rect 24584 4029 24593 4063
rect 24593 4029 24627 4063
rect 24627 4029 24636 4063
rect 24584 4020 24636 4029
rect 26056 4020 26108 4072
rect 27528 4097 27537 4131
rect 27537 4097 27571 4131
rect 27571 4097 27580 4131
rect 27528 4088 27580 4097
rect 28724 4088 28776 4140
rect 30656 4088 30708 4140
rect 30932 4131 30984 4140
rect 30932 4097 30941 4131
rect 30941 4097 30975 4131
rect 30975 4097 30984 4131
rect 30932 4088 30984 4097
rect 27988 4020 28040 4072
rect 28356 4063 28408 4072
rect 28356 4029 28365 4063
rect 28365 4029 28399 4063
rect 28399 4029 28408 4063
rect 28356 4020 28408 4029
rect 29552 4020 29604 4072
rect 30380 4020 30432 4072
rect 30564 4020 30616 4072
rect 19340 3952 19392 4004
rect 29000 3952 29052 4004
rect 17500 3884 17552 3936
rect 11253 3782 11305 3834
rect 11317 3782 11369 3834
rect 11381 3782 11433 3834
rect 11445 3782 11497 3834
rect 11509 3782 11561 3834
rect 21557 3782 21609 3834
rect 21621 3782 21673 3834
rect 21685 3782 21737 3834
rect 21749 3782 21801 3834
rect 21813 3782 21865 3834
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 4160 3680 4212 3732
rect 6736 3680 6788 3732
rect 7104 3680 7156 3732
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 11060 3680 11112 3732
rect 15200 3680 15252 3732
rect 17684 3723 17736 3732
rect 5816 3612 5868 3664
rect 7380 3612 7432 3664
rect 8484 3612 8536 3664
rect 9772 3612 9824 3664
rect 10876 3612 10928 3664
rect 7472 3476 7524 3528
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10692 3544 10744 3596
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 14188 3612 14240 3664
rect 14372 3612 14424 3664
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 18696 3680 18748 3732
rect 19248 3680 19300 3732
rect 23572 3680 23624 3732
rect 24584 3680 24636 3732
rect 24676 3680 24728 3732
rect 16948 3612 17000 3664
rect 12072 3544 12124 3553
rect 16764 3544 16816 3596
rect 19248 3544 19300 3596
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 19800 3587 19852 3596
rect 19800 3553 19809 3587
rect 19809 3553 19843 3587
rect 19843 3553 19852 3587
rect 19800 3544 19852 3553
rect 22836 3544 22888 3596
rect 25228 3612 25280 3664
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 17592 3476 17644 3528
rect 18328 3476 18380 3528
rect 19064 3476 19116 3528
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 20720 3476 20772 3528
rect 21916 3476 21968 3528
rect 24584 3587 24636 3596
rect 24584 3553 24593 3587
rect 24593 3553 24627 3587
rect 24627 3553 24636 3587
rect 24584 3544 24636 3553
rect 24676 3544 24728 3596
rect 25136 3587 25188 3596
rect 25136 3553 25145 3587
rect 25145 3553 25179 3587
rect 25179 3553 25188 3587
rect 25136 3544 25188 3553
rect 25688 3544 25740 3596
rect 26240 3680 26292 3732
rect 27252 3680 27304 3732
rect 27804 3680 27856 3732
rect 28264 3680 28316 3732
rect 30380 3680 30432 3732
rect 30564 3723 30616 3732
rect 30564 3689 30573 3723
rect 30573 3689 30607 3723
rect 30607 3689 30616 3723
rect 30564 3680 30616 3689
rect 30472 3612 30524 3664
rect 27528 3544 27580 3596
rect 27804 3544 27856 3596
rect 28356 3544 28408 3596
rect 28816 3544 28868 3596
rect 30288 3544 30340 3596
rect 24492 3476 24544 3528
rect 24768 3519 24820 3528
rect 24768 3485 24777 3519
rect 24777 3485 24811 3519
rect 24811 3485 24820 3519
rect 24768 3476 24820 3485
rect 25044 3476 25096 3528
rect 18512 3408 18564 3460
rect 21088 3408 21140 3460
rect 8576 3340 8628 3392
rect 10324 3340 10376 3392
rect 11796 3340 11848 3392
rect 17868 3340 17920 3392
rect 24308 3340 24360 3392
rect 25044 3340 25096 3392
rect 25872 3340 25924 3392
rect 26608 3340 26660 3392
rect 6102 3238 6154 3290
rect 6166 3238 6218 3290
rect 6230 3238 6282 3290
rect 6294 3238 6346 3290
rect 6358 3238 6410 3290
rect 16405 3238 16457 3290
rect 16469 3238 16521 3290
rect 16533 3238 16585 3290
rect 16597 3238 16649 3290
rect 16661 3238 16713 3290
rect 26709 3238 26761 3290
rect 26773 3238 26825 3290
rect 26837 3238 26889 3290
rect 26901 3238 26953 3290
rect 26965 3238 27017 3290
rect 2872 3136 2924 3188
rect 4160 3136 4212 3188
rect 5448 3136 5500 3188
rect 7288 3179 7340 3188
rect 7288 3145 7297 3179
rect 7297 3145 7331 3179
rect 7331 3145 7340 3179
rect 7288 3136 7340 3145
rect 8484 3136 8536 3188
rect 9864 3136 9916 3188
rect 11152 3136 11204 3188
rect 12440 3136 12492 3188
rect 16028 3136 16080 3188
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 18236 3136 18288 3188
rect 19340 3179 19392 3188
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 24308 3136 24360 3188
rect 2780 3068 2832 3120
rect 9036 3068 9088 3120
rect 10048 3068 10100 3120
rect 5356 3000 5408 3052
rect 7472 3000 7524 3052
rect 10232 3068 10284 3120
rect 22192 3111 22244 3120
rect 22192 3077 22201 3111
rect 22201 3077 22235 3111
rect 22235 3077 22244 3111
rect 22192 3068 22244 3077
rect 9680 2932 9732 2984
rect 10600 3000 10652 3052
rect 13820 3000 13872 3052
rect 10048 2975 10100 2984
rect 10048 2941 10057 2975
rect 10057 2941 10091 2975
rect 10091 2941 10100 2975
rect 10048 2932 10100 2941
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 10784 2932 10836 2984
rect 6000 2864 6052 2916
rect 12716 2932 12768 2984
rect 17316 2975 17368 2984
rect 11980 2864 12032 2916
rect 16672 2864 16724 2916
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 18052 2864 18104 2916
rect 10600 2839 10652 2848
rect 10600 2805 10609 2839
rect 10609 2805 10643 2839
rect 10643 2805 10652 2839
rect 10600 2796 10652 2805
rect 10968 2796 11020 2848
rect 12716 2796 12768 2848
rect 19800 3000 19852 3052
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 24952 3068 25004 3120
rect 27804 3136 27856 3188
rect 28724 3136 28776 3188
rect 30104 3179 30156 3188
rect 30104 3145 30113 3179
rect 30113 3145 30147 3179
rect 30147 3145 30156 3179
rect 30104 3136 30156 3145
rect 31024 3179 31076 3188
rect 31024 3145 31033 3179
rect 31033 3145 31067 3179
rect 31067 3145 31076 3179
rect 31024 3136 31076 3145
rect 31300 3136 31352 3188
rect 26056 3043 26108 3052
rect 26056 3009 26065 3043
rect 26065 3009 26099 3043
rect 26099 3009 26108 3043
rect 26056 3000 26108 3009
rect 26240 3000 26292 3052
rect 28632 3043 28684 3052
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18512 2975 18564 2984
rect 18328 2932 18380 2941
rect 18512 2941 18521 2975
rect 18521 2941 18555 2975
rect 18555 2941 18564 2975
rect 18512 2932 18564 2941
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 19064 2932 19116 2984
rect 22100 2932 22152 2984
rect 22376 2932 22428 2984
rect 23388 2975 23440 2984
rect 23388 2941 23397 2975
rect 23397 2941 23431 2975
rect 23431 2941 23440 2975
rect 23388 2932 23440 2941
rect 23572 2932 23624 2984
rect 23756 2932 23808 2984
rect 25136 2975 25188 2984
rect 21364 2864 21416 2916
rect 21916 2864 21968 2916
rect 22836 2864 22888 2916
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 25964 2975 26016 2984
rect 19708 2796 19760 2848
rect 22192 2796 22244 2848
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 26608 2932 26660 2984
rect 27160 2932 27212 2984
rect 28632 3009 28641 3043
rect 28641 3009 28675 3043
rect 28675 3009 28684 3043
rect 28632 3000 28684 3009
rect 28540 2932 28592 2984
rect 28908 2932 28960 2984
rect 27344 2864 27396 2916
rect 29092 2932 29144 2984
rect 29184 2864 29236 2916
rect 26240 2796 26292 2848
rect 27068 2796 27120 2848
rect 28080 2796 28132 2848
rect 28172 2796 28224 2848
rect 28816 2796 28868 2848
rect 11253 2694 11305 2746
rect 11317 2694 11369 2746
rect 11381 2694 11433 2746
rect 11445 2694 11497 2746
rect 11509 2694 11561 2746
rect 21557 2694 21609 2746
rect 21621 2694 21673 2746
rect 21685 2694 21737 2746
rect 21749 2694 21801 2746
rect 21813 2694 21865 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 3148 2592 3200 2644
rect 3240 2635 3292 2644
rect 3240 2601 3249 2635
rect 3249 2601 3283 2635
rect 3283 2601 3292 2635
rect 4160 2635 4212 2644
rect 3240 2592 3292 2601
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 5448 2592 5500 2644
rect 7104 2592 7156 2644
rect 8576 2592 8628 2644
rect 9680 2592 9732 2644
rect 12716 2635 12768 2644
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 10324 2456 10376 2508
rect 12716 2601 12725 2635
rect 12725 2601 12759 2635
rect 12759 2601 12768 2635
rect 12716 2592 12768 2601
rect 14280 2592 14332 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 10692 2524 10744 2576
rect 10784 2499 10836 2508
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 13176 2524 13228 2576
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 11980 2456 12032 2508
rect 10232 2388 10284 2440
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 15936 2524 15988 2576
rect 15384 2456 15436 2508
rect 17224 2592 17276 2644
rect 17776 2524 17828 2576
rect 14740 2431 14792 2440
rect 14740 2397 14749 2431
rect 14749 2397 14783 2431
rect 14783 2397 14792 2431
rect 14740 2388 14792 2397
rect 16028 2388 16080 2440
rect 15936 2320 15988 2372
rect 17408 2499 17460 2508
rect 17408 2465 17413 2499
rect 17413 2465 17447 2499
rect 17447 2465 17460 2499
rect 17408 2456 17460 2465
rect 18052 2499 18104 2508
rect 18052 2465 18061 2499
rect 18061 2465 18095 2499
rect 18095 2465 18104 2499
rect 18052 2456 18104 2465
rect 18420 2499 18472 2508
rect 17960 2388 18012 2440
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 18696 2456 18748 2508
rect 19248 2499 19300 2508
rect 19248 2465 19257 2499
rect 19257 2465 19291 2499
rect 19291 2465 19300 2499
rect 19248 2456 19300 2465
rect 19800 2524 19852 2576
rect 19524 2456 19576 2508
rect 20260 2456 20312 2508
rect 22008 2592 22060 2644
rect 23664 2592 23716 2644
rect 24584 2592 24636 2644
rect 24860 2592 24912 2644
rect 26056 2592 26108 2644
rect 28540 2592 28592 2644
rect 29552 2635 29604 2644
rect 29552 2601 29561 2635
rect 29561 2601 29595 2635
rect 29595 2601 29604 2635
rect 29552 2592 29604 2601
rect 30932 2592 30984 2644
rect 22192 2524 22244 2576
rect 25044 2456 25096 2508
rect 26608 2524 26660 2576
rect 25228 2456 25280 2508
rect 27344 2456 27396 2508
rect 28080 2456 28132 2508
rect 28264 2499 28316 2508
rect 28264 2465 28273 2499
rect 28273 2465 28307 2499
rect 28307 2465 28316 2499
rect 28264 2456 28316 2465
rect 28816 2499 28868 2508
rect 28816 2465 28825 2499
rect 28825 2465 28859 2499
rect 28859 2465 28868 2499
rect 28816 2456 28868 2465
rect 18052 2320 18104 2372
rect 18880 2320 18932 2372
rect 10140 2252 10192 2304
rect 10692 2252 10744 2304
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 17040 2252 17092 2304
rect 18604 2295 18656 2304
rect 18604 2261 18613 2295
rect 18613 2261 18647 2295
rect 18647 2261 18656 2295
rect 18604 2252 18656 2261
rect 19616 2320 19668 2372
rect 21364 2388 21416 2440
rect 28632 2431 28684 2440
rect 19800 2295 19852 2304
rect 19800 2261 19809 2295
rect 19809 2261 19843 2295
rect 19843 2261 19852 2295
rect 19800 2252 19852 2261
rect 24768 2252 24820 2304
rect 25780 2252 25832 2304
rect 28632 2397 28641 2431
rect 28641 2397 28675 2431
rect 28675 2397 28684 2431
rect 28632 2388 28684 2397
rect 28264 2320 28316 2372
rect 29184 2320 29236 2372
rect 30104 2320 30156 2372
rect 27344 2252 27396 2304
rect 6102 2150 6154 2202
rect 6166 2150 6218 2202
rect 6230 2150 6282 2202
rect 6294 2150 6346 2202
rect 6358 2150 6410 2202
rect 16405 2150 16457 2202
rect 16469 2150 16521 2202
rect 16533 2150 16585 2202
rect 16597 2150 16649 2202
rect 16661 2150 16713 2202
rect 26709 2150 26761 2202
rect 26773 2150 26825 2202
rect 26837 2150 26889 2202
rect 26901 2150 26953 2202
rect 26965 2150 27017 2202
rect 1492 2091 1544 2100
rect 1492 2057 1501 2091
rect 1501 2057 1535 2091
rect 1535 2057 1544 2091
rect 1492 2048 1544 2057
rect 2136 2048 2188 2100
rect 3332 2048 3384 2100
rect 3424 2048 3476 2100
rect 6000 2091 6052 2100
rect 6000 2057 6009 2091
rect 6009 2057 6043 2091
rect 6043 2057 6052 2091
rect 9588 2091 9640 2100
rect 6000 2048 6052 2057
rect 9588 2057 9597 2091
rect 9597 2057 9631 2091
rect 9631 2057 9640 2091
rect 9588 2048 9640 2057
rect 2596 1980 2648 2032
rect 5448 1980 5500 2032
rect 8392 2023 8444 2032
rect 8392 1989 8401 2023
rect 8401 1989 8435 2023
rect 8435 1989 8444 2023
rect 8392 1980 8444 1989
rect 9128 1980 9180 2032
rect 12072 2048 12124 2100
rect 12992 2048 13044 2100
rect 13268 2091 13320 2100
rect 13268 2057 13277 2091
rect 13277 2057 13311 2091
rect 13311 2057 13320 2091
rect 13268 2048 13320 2057
rect 16856 2048 16908 2100
rect 10048 1980 10100 2032
rect 18788 2048 18840 2100
rect 19248 2048 19300 2100
rect 22836 2091 22888 2100
rect 22836 2057 22845 2091
rect 22845 2057 22879 2091
rect 22879 2057 22888 2091
rect 22836 2048 22888 2057
rect 23112 2048 23164 2100
rect 24676 2048 24728 2100
rect 24860 2048 24912 2100
rect 26332 2091 26384 2100
rect 13820 1912 13872 1964
rect 14740 1912 14792 1964
rect 26332 2057 26341 2091
rect 26341 2057 26375 2091
rect 26375 2057 26384 2091
rect 26332 2048 26384 2057
rect 28816 2048 28868 2100
rect 30012 2048 30064 2100
rect 26424 1912 26476 1964
rect 10876 1844 10928 1896
rect 14372 1887 14424 1896
rect 14372 1853 14381 1887
rect 14381 1853 14415 1887
rect 14415 1853 14424 1887
rect 14372 1844 14424 1853
rect 15752 1844 15804 1896
rect 18604 1844 18656 1896
rect 20260 1844 20312 1896
rect 25872 1844 25924 1896
rect 12256 1776 12308 1828
rect 20720 1819 20772 1828
rect 20720 1785 20738 1819
rect 20738 1785 20772 1819
rect 20720 1776 20772 1785
rect 22652 1776 22704 1828
rect 25688 1776 25740 1828
rect 27344 1819 27396 1828
rect 27344 1785 27378 1819
rect 27378 1785 27396 1819
rect 27344 1776 27396 1785
rect 27528 1776 27580 1828
rect 29000 1776 29052 1828
rect 30104 1819 30156 1828
rect 30104 1785 30113 1819
rect 30113 1785 30147 1819
rect 30147 1785 30156 1819
rect 30104 1776 30156 1785
rect 16212 1708 16264 1760
rect 16948 1708 17000 1760
rect 17316 1751 17368 1760
rect 17316 1717 17325 1751
rect 17325 1717 17359 1751
rect 17359 1717 17368 1751
rect 17316 1708 17368 1717
rect 18420 1708 18472 1760
rect 30932 1751 30984 1760
rect 30932 1717 30941 1751
rect 30941 1717 30975 1751
rect 30975 1717 30984 1751
rect 30932 1708 30984 1717
rect 11253 1606 11305 1658
rect 11317 1606 11369 1658
rect 11381 1606 11433 1658
rect 11445 1606 11497 1658
rect 11509 1606 11561 1658
rect 21557 1606 21609 1658
rect 21621 1606 21673 1658
rect 21685 1606 21737 1658
rect 21749 1606 21801 1658
rect 21813 1606 21865 1658
rect 8392 1504 8444 1556
rect 9128 1547 9180 1556
rect 9128 1513 9137 1547
rect 9137 1513 9171 1547
rect 9171 1513 9180 1547
rect 9128 1504 9180 1513
rect 9680 1504 9732 1556
rect 13360 1504 13412 1556
rect 14372 1504 14424 1556
rect 10600 1436 10652 1488
rect 1860 1411 1912 1420
rect 1860 1377 1869 1411
rect 1869 1377 1903 1411
rect 1903 1377 1912 1411
rect 1860 1368 1912 1377
rect 10876 1368 10928 1420
rect 2964 1300 3016 1352
rect 13820 1436 13872 1488
rect 14004 1368 14056 1420
rect 15936 1504 15988 1556
rect 18880 1547 18932 1556
rect 18880 1513 18889 1547
rect 18889 1513 18923 1547
rect 18923 1513 18932 1547
rect 18880 1504 18932 1513
rect 21456 1504 21508 1556
rect 29000 1547 29052 1556
rect 17316 1436 17368 1488
rect 19064 1436 19116 1488
rect 19800 1436 19852 1488
rect 29000 1513 29009 1547
rect 29009 1513 29043 1547
rect 29043 1513 29052 1547
rect 29000 1504 29052 1513
rect 30012 1547 30064 1556
rect 30012 1513 30021 1547
rect 30021 1513 30055 1547
rect 30055 1513 30064 1547
rect 30012 1504 30064 1513
rect 16764 1368 16816 1420
rect 17408 1368 17460 1420
rect 17500 1368 17552 1420
rect 22836 1368 22888 1420
rect 29092 1436 29144 1488
rect 13176 1343 13228 1352
rect 13176 1309 13185 1343
rect 13185 1309 13219 1343
rect 13219 1309 13228 1343
rect 13176 1300 13228 1309
rect 15384 1343 15436 1352
rect 15384 1309 15393 1343
rect 15393 1309 15427 1343
rect 15427 1309 15436 1343
rect 15384 1300 15436 1309
rect 7380 1232 7432 1284
rect 12164 1232 12216 1284
rect 16028 1300 16080 1352
rect 19156 1300 19208 1352
rect 20260 1343 20312 1352
rect 20260 1309 20269 1343
rect 20269 1309 20303 1343
rect 20303 1309 20312 1343
rect 20260 1300 20312 1309
rect 22652 1300 22704 1352
rect 17132 1232 17184 1284
rect 23388 1300 23440 1352
rect 24584 1368 24636 1420
rect 25136 1368 25188 1420
rect 25596 1368 25648 1420
rect 26424 1411 26476 1420
rect 26424 1377 26433 1411
rect 26433 1377 26467 1411
rect 26467 1377 26476 1411
rect 26424 1368 26476 1377
rect 28172 1411 28224 1420
rect 28172 1377 28190 1411
rect 28190 1377 28224 1411
rect 28172 1368 28224 1377
rect 30472 1368 30524 1420
rect 24768 1232 24820 1284
rect 10600 1164 10652 1216
rect 12992 1164 13044 1216
rect 25504 1164 25556 1216
rect 25688 1164 25740 1216
rect 26148 1164 26200 1216
rect 27528 1164 27580 1216
rect 6102 1062 6154 1114
rect 6166 1062 6218 1114
rect 6230 1062 6282 1114
rect 6294 1062 6346 1114
rect 6358 1062 6410 1114
rect 16405 1062 16457 1114
rect 16469 1062 16521 1114
rect 16533 1062 16585 1114
rect 16597 1062 16649 1114
rect 16661 1062 16713 1114
rect 26709 1062 26761 1114
rect 26773 1062 26825 1114
rect 26837 1062 26889 1114
rect 26901 1062 26953 1114
rect 26965 1062 27017 1114
rect 1860 960 1912 1012
rect 8392 1003 8444 1012
rect 8392 969 8401 1003
rect 8401 969 8435 1003
rect 8435 969 8444 1003
rect 8392 960 8444 969
rect 14464 960 14516 1012
rect 15844 960 15896 1012
rect 16120 960 16172 1012
rect 17500 1003 17552 1012
rect 17500 969 17509 1003
rect 17509 969 17543 1003
rect 17543 969 17552 1003
rect 17500 960 17552 969
rect 18512 960 18564 1012
rect 18972 960 19024 1012
rect 19432 1003 19484 1012
rect 19432 969 19441 1003
rect 19441 969 19475 1003
rect 19475 969 19484 1003
rect 19432 960 19484 969
rect 20812 960 20864 1012
rect 20904 960 20956 1012
rect 22284 960 22336 1012
rect 22744 960 22796 1012
rect 29000 960 29052 1012
rect 8300 892 8352 944
rect 11704 892 11756 944
rect 14004 892 14056 944
rect 20076 892 20128 944
rect 23020 935 23072 944
rect 23020 901 23029 935
rect 23029 901 23063 935
rect 23063 901 23072 935
rect 23020 892 23072 901
rect 23204 892 23256 944
rect 25596 892 25648 944
rect 25688 892 25740 944
rect 13176 867 13228 876
rect 13176 833 13185 867
rect 13185 833 13219 867
rect 13219 833 13228 867
rect 13176 824 13228 833
rect 16028 824 16080 876
rect 17224 824 17276 876
rect 25964 867 26016 876
rect 25964 833 25973 867
rect 25973 833 26007 867
rect 26007 833 26016 867
rect 25964 824 26016 833
rect 27160 824 27212 876
rect 12900 799 12952 808
rect 12900 765 12918 799
rect 12918 765 12952 799
rect 12900 756 12952 765
rect 13912 756 13964 808
rect 15936 799 15988 808
rect 15936 765 15945 799
rect 15945 765 15979 799
rect 15979 765 15988 799
rect 15936 756 15988 765
rect 16764 799 16816 808
rect 16764 765 16773 799
rect 16773 765 16807 799
rect 16807 765 16816 799
rect 16764 756 16816 765
rect 16948 799 17000 808
rect 16948 765 16957 799
rect 16957 765 16991 799
rect 16991 765 17000 799
rect 16948 756 17000 765
rect 17316 799 17368 808
rect 17316 765 17325 799
rect 17325 765 17359 799
rect 17359 765 17368 799
rect 17316 756 17368 765
rect 19432 756 19484 808
rect 24032 756 24084 808
rect 24952 799 25004 808
rect 24952 765 24961 799
rect 24961 765 24995 799
rect 24995 765 25004 799
rect 24952 756 25004 765
rect 25504 756 25556 808
rect 25780 756 25832 808
rect 26148 756 26200 808
rect 26240 799 26292 808
rect 26240 765 26249 799
rect 26249 765 26283 799
rect 26283 765 26292 799
rect 26240 756 26292 765
rect 26700 756 26752 808
rect 30932 756 30984 808
rect 9496 663 9548 672
rect 9496 629 9505 663
rect 9505 629 9539 663
rect 9539 629 9548 663
rect 9496 620 9548 629
rect 14648 620 14700 672
rect 20168 663 20220 672
rect 20168 629 20177 663
rect 20177 629 20211 663
rect 20211 629 20220 663
rect 20168 620 20220 629
rect 25688 620 25740 672
rect 26148 620 26200 672
rect 11253 518 11305 570
rect 11317 518 11369 570
rect 11381 518 11433 570
rect 11445 518 11497 570
rect 11509 518 11561 570
rect 21557 518 21609 570
rect 21621 518 21673 570
rect 21685 518 21737 570
rect 21749 518 21801 570
rect 21813 518 21865 570
rect 9496 416 9548 468
rect 23020 416 23072 468
rect 24952 416 25004 468
rect 26148 416 26200 468
rect 20168 348 20220 400
rect 26700 348 26752 400
<< metal2 >>
rect 8298 48160 8354 48960
rect 11253 48444 11561 48464
rect 11253 48442 11259 48444
rect 11315 48442 11339 48444
rect 11395 48442 11419 48444
rect 11475 48442 11499 48444
rect 11555 48442 11561 48444
rect 11315 48390 11317 48442
rect 11497 48390 11499 48442
rect 11253 48388 11259 48390
rect 11315 48388 11339 48390
rect 11395 48388 11419 48390
rect 11475 48388 11499 48390
rect 11555 48388 11561 48390
rect 11253 48368 11561 48388
rect 21557 48444 21865 48464
rect 21557 48442 21563 48444
rect 21619 48442 21643 48444
rect 21699 48442 21723 48444
rect 21779 48442 21803 48444
rect 21859 48442 21865 48444
rect 21619 48390 21621 48442
rect 21801 48390 21803 48442
rect 21557 48388 21563 48390
rect 21619 48388 21643 48390
rect 21699 48388 21723 48390
rect 21779 48388 21803 48390
rect 21859 48388 21865 48390
rect 21557 48368 21865 48388
rect 8484 48204 8536 48210
rect 8312 48074 8340 48160
rect 8484 48146 8536 48152
rect 15844 48204 15896 48210
rect 15844 48146 15896 48152
rect 24768 48204 24820 48210
rect 24858 48160 24914 48960
rect 31300 48204 31352 48210
rect 24768 48146 24820 48152
rect 8300 48068 8352 48074
rect 8300 48010 8352 48016
rect 5724 48000 5776 48006
rect 5724 47942 5776 47948
rect 1400 46028 1452 46034
rect 1400 45970 1452 45976
rect 1412 45626 1440 45970
rect 4988 45824 5040 45830
rect 4988 45766 5040 45772
rect 1400 45620 1452 45626
rect 1400 45562 1452 45568
rect 2688 44532 2740 44538
rect 2688 44474 2740 44480
rect 1860 44260 1912 44266
rect 1860 44202 1912 44208
rect 1872 43926 1900 44202
rect 1860 43920 1912 43926
rect 1860 43862 1912 43868
rect 2136 43648 2188 43654
rect 2136 43590 2188 43596
rect 1584 43104 1636 43110
rect 1584 43046 1636 43052
rect 1768 43104 1820 43110
rect 1768 43046 1820 43052
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1400 40588 1452 40594
rect 1400 40530 1452 40536
rect 1412 39846 1440 40530
rect 1400 39840 1452 39846
rect 1400 39782 1452 39788
rect 1400 39500 1452 39506
rect 1400 39442 1452 39448
rect 1412 38962 1440 39442
rect 1400 38956 1452 38962
rect 1400 38898 1452 38904
rect 1504 36394 1532 42502
rect 1412 36366 1532 36394
rect 1412 34066 1440 36366
rect 1596 36122 1624 43046
rect 1676 39840 1728 39846
rect 1676 39782 1728 39788
rect 1688 39506 1716 39782
rect 1676 39500 1728 39506
rect 1676 39442 1728 39448
rect 1780 38978 1808 43046
rect 2044 42560 2096 42566
rect 2044 42502 2096 42508
rect 1860 41472 1912 41478
rect 1860 41414 1912 41420
rect 1688 38950 1808 38978
rect 1688 36666 1716 38950
rect 1768 38820 1820 38826
rect 1768 38762 1820 38768
rect 1780 38554 1808 38762
rect 1768 38548 1820 38554
rect 1768 38490 1820 38496
rect 1768 38412 1820 38418
rect 1768 38354 1820 38360
rect 1780 36786 1808 38354
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1688 36638 1808 36666
rect 1676 36576 1728 36582
rect 1676 36518 1728 36524
rect 1688 36242 1716 36518
rect 1676 36236 1728 36242
rect 1676 36178 1728 36184
rect 1780 36122 1808 36638
rect 1504 36094 1624 36122
rect 1688 36094 1808 36122
rect 1400 34060 1452 34066
rect 1400 34002 1452 34008
rect 1400 33856 1452 33862
rect 1400 33798 1452 33804
rect 1308 31748 1360 31754
rect 1308 31690 1360 31696
rect 1216 29776 1268 29782
rect 1216 29718 1268 29724
rect 1228 28150 1256 29718
rect 1320 28218 1348 31690
rect 1412 29306 1440 33798
rect 1400 29300 1452 29306
rect 1400 29242 1452 29248
rect 1308 28212 1360 28218
rect 1308 28154 1360 28160
rect 1216 28144 1268 28150
rect 1216 28086 1268 28092
rect 1320 27334 1348 28154
rect 1504 28014 1532 36094
rect 1688 36020 1716 36094
rect 1872 36020 1900 41414
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1596 35992 1716 36020
rect 1780 35992 1900 36020
rect 1596 31686 1624 35992
rect 1676 34536 1728 34542
rect 1676 34478 1728 34484
rect 1688 33046 1716 34478
rect 1676 33040 1728 33046
rect 1676 32982 1728 32988
rect 1676 32768 1728 32774
rect 1676 32710 1728 32716
rect 1688 32434 1716 32710
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1676 32292 1728 32298
rect 1676 32234 1728 32240
rect 1688 31890 1716 32234
rect 1676 31884 1728 31890
rect 1676 31826 1728 31832
rect 1584 31680 1636 31686
rect 1584 31622 1636 31628
rect 1596 31278 1624 31622
rect 1584 31272 1636 31278
rect 1584 31214 1636 31220
rect 1780 30802 1808 35992
rect 1964 33912 1992 40326
rect 2056 37806 2084 42502
rect 2148 42158 2176 43590
rect 2320 42560 2372 42566
rect 2320 42502 2372 42508
rect 2136 42152 2188 42158
rect 2136 42094 2188 42100
rect 2228 39976 2280 39982
rect 2228 39918 2280 39924
rect 2136 39500 2188 39506
rect 2136 39442 2188 39448
rect 2148 38350 2176 39442
rect 2240 38758 2268 39918
rect 2228 38752 2280 38758
rect 2228 38694 2280 38700
rect 2240 38554 2268 38694
rect 2228 38548 2280 38554
rect 2228 38490 2280 38496
rect 2136 38344 2188 38350
rect 2136 38286 2188 38292
rect 2044 37800 2096 37806
rect 2044 37742 2096 37748
rect 2148 37618 2176 38286
rect 2056 37590 2176 37618
rect 2056 36786 2084 37590
rect 2136 37324 2188 37330
rect 2136 37266 2188 37272
rect 2044 36780 2096 36786
rect 2044 36722 2096 36728
rect 2148 36718 2176 37266
rect 2228 37120 2280 37126
rect 2228 37062 2280 37068
rect 2136 36712 2188 36718
rect 2136 36654 2188 36660
rect 2044 36644 2096 36650
rect 2044 36586 2096 36592
rect 2056 35170 2084 36586
rect 2148 36038 2176 36654
rect 2136 36032 2188 36038
rect 2136 35974 2188 35980
rect 2240 35290 2268 37062
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 2056 35142 2268 35170
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 2056 34542 2084 35022
rect 2240 34542 2268 35142
rect 2044 34536 2096 34542
rect 2228 34536 2280 34542
rect 2096 34496 2176 34524
rect 2044 34478 2096 34484
rect 1872 33884 1992 33912
rect 1768 30796 1820 30802
rect 1768 30738 1820 30744
rect 1676 30048 1728 30054
rect 1676 29990 1728 29996
rect 1584 29708 1636 29714
rect 1584 29650 1636 29656
rect 1596 29034 1624 29650
rect 1584 29028 1636 29034
rect 1584 28970 1636 28976
rect 1492 28008 1544 28014
rect 1492 27950 1544 27956
rect 1504 27674 1532 27950
rect 1492 27668 1544 27674
rect 1492 27610 1544 27616
rect 1596 27606 1624 28970
rect 1688 28558 1716 29990
rect 1780 29646 1808 30738
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1768 29300 1820 29306
rect 1768 29242 1820 29248
rect 1676 28552 1728 28558
rect 1676 28494 1728 28500
rect 1584 27600 1636 27606
rect 1584 27542 1636 27548
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1308 27328 1360 27334
rect 1308 27270 1360 27276
rect 1412 26042 1440 27406
rect 1676 27396 1728 27402
rect 1676 27338 1728 27344
rect 1688 27010 1716 27338
rect 1780 27130 1808 29242
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1688 26982 1808 27010
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22098 1440 23054
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1504 21026 1532 25094
rect 1584 23520 1636 23526
rect 1584 23462 1636 23468
rect 1228 20998 1532 21026
rect 1228 16794 1256 20998
rect 1400 20868 1452 20874
rect 1400 20810 1452 20816
rect 1308 20052 1360 20058
rect 1308 19994 1360 20000
rect 1216 16788 1268 16794
rect 1216 16730 1268 16736
rect 1320 15910 1348 19994
rect 1412 18952 1440 20810
rect 1596 20346 1624 23462
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 1688 21690 1716 22034
rect 1676 21684 1728 21690
rect 1676 21626 1728 21632
rect 1504 20318 1624 20346
rect 1504 20058 1532 20318
rect 1780 20262 1808 26982
rect 1872 26246 1900 33884
rect 2044 33448 2096 33454
rect 2044 33390 2096 33396
rect 1952 33312 2004 33318
rect 1952 33254 2004 33260
rect 1964 31822 1992 33254
rect 2056 33114 2084 33390
rect 2148 33318 2176 34496
rect 2228 34478 2280 34484
rect 2136 33312 2188 33318
rect 2136 33254 2188 33260
rect 2044 33108 2096 33114
rect 2044 33050 2096 33056
rect 2240 32978 2268 34478
rect 2228 32972 2280 32978
rect 2228 32914 2280 32920
rect 2044 32904 2096 32910
rect 2044 32846 2096 32852
rect 2056 32570 2084 32846
rect 2136 32836 2188 32842
rect 2136 32778 2188 32784
rect 2044 32564 2096 32570
rect 2044 32506 2096 32512
rect 2044 32428 2096 32434
rect 2044 32370 2096 32376
rect 1952 31816 2004 31822
rect 1952 31758 2004 31764
rect 2056 30870 2084 32370
rect 2148 30938 2176 32778
rect 2240 32502 2268 32914
rect 2228 32496 2280 32502
rect 2228 32438 2280 32444
rect 2228 32224 2280 32230
rect 2228 32166 2280 32172
rect 2240 31890 2268 32166
rect 2228 31884 2280 31890
rect 2228 31826 2280 31832
rect 2332 31754 2360 42502
rect 2700 41818 2728 44474
rect 2872 43104 2924 43110
rect 2872 43046 2924 43052
rect 2964 43104 3016 43110
rect 2964 43046 3016 43052
rect 4160 43104 4212 43110
rect 4160 43046 4212 43052
rect 2688 41812 2740 41818
rect 2688 41754 2740 41760
rect 2504 40928 2556 40934
rect 2504 40870 2556 40876
rect 2516 40050 2544 40870
rect 2884 40730 2912 43046
rect 2872 40724 2924 40730
rect 2872 40666 2924 40672
rect 2780 40656 2832 40662
rect 2780 40598 2832 40604
rect 2504 40044 2556 40050
rect 2504 39986 2556 39992
rect 2412 39976 2464 39982
rect 2412 39918 2464 39924
rect 2424 38418 2452 39918
rect 2516 38826 2544 39986
rect 2596 39840 2648 39846
rect 2596 39782 2648 39788
rect 2688 39840 2740 39846
rect 2688 39782 2740 39788
rect 2608 39386 2636 39782
rect 2700 39506 2728 39782
rect 2792 39574 2820 40598
rect 2780 39568 2832 39574
rect 2780 39510 2832 39516
rect 2688 39500 2740 39506
rect 2688 39442 2740 39448
rect 2608 39358 2728 39386
rect 2700 39302 2728 39358
rect 2688 39296 2740 39302
rect 2688 39238 2740 39244
rect 2504 38820 2556 38826
rect 2504 38762 2556 38768
rect 2516 38554 2544 38762
rect 2700 38654 2728 39238
rect 2700 38626 2912 38654
rect 2504 38548 2556 38554
rect 2504 38490 2556 38496
rect 2412 38412 2464 38418
rect 2412 38354 2464 38360
rect 2424 36718 2452 38354
rect 2516 37330 2544 38490
rect 2596 38344 2648 38350
rect 2596 38286 2648 38292
rect 2608 37670 2636 38286
rect 2596 37664 2648 37670
rect 2596 37606 2648 37612
rect 2504 37324 2556 37330
rect 2504 37266 2556 37272
rect 2412 36712 2464 36718
rect 2412 36654 2464 36660
rect 2424 35698 2452 36654
rect 2608 36122 2636 37606
rect 2884 36650 2912 38626
rect 2872 36644 2924 36650
rect 2872 36586 2924 36592
rect 2608 36094 2728 36122
rect 2412 35692 2464 35698
rect 2412 35634 2464 35640
rect 2412 34672 2464 34678
rect 2412 34614 2464 34620
rect 2424 33590 2452 34614
rect 2504 34400 2556 34406
rect 2504 34342 2556 34348
rect 2516 34134 2544 34342
rect 2504 34128 2556 34134
rect 2504 34070 2556 34076
rect 2412 33584 2464 33590
rect 2412 33526 2464 33532
rect 2424 32502 2452 33526
rect 2516 32570 2544 34070
rect 2596 33380 2648 33386
rect 2596 33322 2648 33328
rect 2504 32564 2556 32570
rect 2504 32506 2556 32512
rect 2412 32496 2464 32502
rect 2608 32450 2636 33322
rect 2412 32438 2464 32444
rect 2516 32422 2636 32450
rect 2516 31906 2544 32422
rect 2596 32360 2648 32366
rect 2596 32302 2648 32308
rect 2608 31958 2636 32302
rect 2240 31726 2360 31754
rect 2424 31878 2544 31906
rect 2596 31952 2648 31958
rect 2596 31894 2648 31900
rect 2136 30932 2188 30938
rect 2136 30874 2188 30880
rect 2044 30864 2096 30870
rect 2044 30806 2096 30812
rect 2056 30394 2084 30806
rect 2044 30388 2096 30394
rect 2044 30330 2096 30336
rect 1952 30184 2004 30190
rect 1952 30126 2004 30132
rect 1964 29714 1992 30126
rect 1952 29708 2004 29714
rect 2240 29696 2268 31726
rect 2320 31680 2372 31686
rect 2320 31622 2372 31628
rect 2332 31414 2360 31622
rect 2320 31408 2372 31414
rect 2320 31350 2372 31356
rect 2332 30734 2360 31350
rect 2424 30802 2452 31878
rect 2700 31804 2728 36094
rect 2780 36032 2832 36038
rect 2780 35974 2832 35980
rect 2792 35154 2820 35974
rect 2780 35148 2832 35154
rect 2780 35090 2832 35096
rect 2792 34474 2820 35090
rect 2884 35086 2912 36586
rect 2872 35080 2924 35086
rect 2872 35022 2924 35028
rect 2872 34944 2924 34950
rect 2872 34886 2924 34892
rect 2780 34468 2832 34474
rect 2780 34410 2832 34416
rect 2792 33930 2820 34410
rect 2780 33924 2832 33930
rect 2780 33866 2832 33872
rect 2884 33386 2912 34886
rect 2872 33380 2924 33386
rect 2792 33340 2872 33368
rect 2792 32230 2820 33340
rect 2872 33322 2924 33328
rect 2872 32972 2924 32978
rect 2872 32914 2924 32920
rect 2780 32224 2832 32230
rect 2780 32166 2832 32172
rect 2884 32026 2912 32914
rect 2872 32020 2924 32026
rect 2872 31962 2924 31968
rect 2608 31776 2728 31804
rect 2412 30796 2464 30802
rect 2412 30738 2464 30744
rect 2320 30728 2372 30734
rect 2320 30670 2372 30676
rect 2504 30184 2556 30190
rect 2504 30126 2556 30132
rect 1952 29650 2004 29656
rect 2237 29668 2268 29696
rect 2237 29594 2265 29668
rect 1952 29572 2004 29578
rect 2148 29566 2265 29594
rect 2004 29532 2084 29560
rect 1952 29514 2004 29520
rect 1952 28620 2004 28626
rect 1952 28562 2004 28568
rect 1964 27606 1992 28562
rect 1952 27600 2004 27606
rect 1952 27542 2004 27548
rect 2056 27538 2084 29532
rect 2044 27532 2096 27538
rect 2044 27474 2096 27480
rect 1952 26852 2004 26858
rect 1952 26794 2004 26800
rect 1964 26450 1992 26794
rect 2056 26586 2084 27474
rect 2044 26580 2096 26586
rect 2044 26522 2096 26528
rect 1952 26444 2004 26450
rect 1952 26386 2004 26392
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1964 25226 1992 26386
rect 1952 25220 2004 25226
rect 1952 25162 2004 25168
rect 1964 24750 1992 25162
rect 1952 24744 2004 24750
rect 1952 24686 2004 24692
rect 1860 24676 1912 24682
rect 1860 24618 1912 24624
rect 1872 23662 1900 24618
rect 1964 24410 1992 24686
rect 2056 24614 2084 26522
rect 2148 24682 2176 29566
rect 2516 29288 2544 30126
rect 2332 29260 2544 29288
rect 2332 28490 2360 29260
rect 2504 29164 2556 29170
rect 2504 29106 2556 29112
rect 2320 28484 2372 28490
rect 2320 28426 2372 28432
rect 2228 27532 2280 27538
rect 2332 27520 2360 28426
rect 2412 28416 2464 28422
rect 2412 28358 2464 28364
rect 2424 28218 2452 28358
rect 2412 28212 2464 28218
rect 2412 28154 2464 28160
rect 2280 27492 2360 27520
rect 2228 27474 2280 27480
rect 2136 24676 2188 24682
rect 2136 24618 2188 24624
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 2056 24410 2084 24550
rect 1952 24404 2004 24410
rect 1952 24346 2004 24352
rect 2044 24404 2096 24410
rect 2044 24346 2096 24352
rect 2240 24290 2268 27474
rect 2320 26240 2372 26246
rect 2320 26182 2372 26188
rect 2056 24274 2268 24290
rect 2044 24268 2268 24274
rect 2096 24262 2268 24268
rect 2044 24210 2096 24216
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2044 24132 2096 24138
rect 2044 24074 2096 24080
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1952 22772 2004 22778
rect 1952 22714 2004 22720
rect 1964 21554 1992 22714
rect 2056 22574 2084 24074
rect 2148 22636 2176 24142
rect 2240 23322 2268 24262
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 2148 22574 2179 22636
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 2139 22568 2191 22574
rect 2139 22510 2191 22516
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 1860 21072 1912 21078
rect 1860 21014 1912 21020
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1492 20052 1544 20058
rect 1492 19994 1544 20000
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1504 19446 1532 19858
rect 1492 19440 1544 19446
rect 1492 19382 1544 19388
rect 1412 18924 1532 18952
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17746 1440 18770
rect 1504 18630 1532 18924
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17746 1532 18022
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1492 17740 1544 17746
rect 1492 17682 1544 17688
rect 1412 16658 1440 17682
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1308 15904 1360 15910
rect 1308 15846 1360 15852
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1504 15366 1532 15506
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1400 13796 1452 13802
rect 1400 13738 1452 13744
rect 1412 13530 1440 13738
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12306 1440 13262
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7342 1440 8230
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1504 2106 1532 15302
rect 1596 12442 1624 20198
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1688 18834 1716 19858
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1780 19514 1808 19654
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 15162 1716 18566
rect 1780 17814 1808 18702
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1780 17338 1808 17750
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1780 14074 1808 14826
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1676 13456 1728 13462
rect 1676 13398 1728 13404
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1596 8480 1624 11154
rect 1688 9178 1716 13398
rect 1872 13274 1900 21014
rect 1964 18766 1992 21490
rect 2044 21480 2096 21486
rect 2148 21468 2176 22510
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2240 21486 2268 22374
rect 2332 22094 2360 26182
rect 2424 24614 2452 28154
rect 2516 27470 2544 29106
rect 2504 27464 2556 27470
rect 2504 27406 2556 27412
rect 2516 26926 2544 27406
rect 2504 26920 2556 26926
rect 2504 26862 2556 26868
rect 2608 26874 2636 31776
rect 2976 31754 3004 43046
rect 4172 42566 4200 43046
rect 3056 42560 3108 42566
rect 3056 42502 3108 42508
rect 4160 42560 4212 42566
rect 4160 42502 4212 42508
rect 4252 42560 4304 42566
rect 4252 42502 4304 42508
rect 3068 35766 3096 42502
rect 3700 41676 3752 41682
rect 3700 41618 3752 41624
rect 3240 41472 3292 41478
rect 3240 41414 3292 41420
rect 3252 41274 3280 41414
rect 3240 41268 3292 41274
rect 3240 41210 3292 41216
rect 3516 40996 3568 41002
rect 3516 40938 3568 40944
rect 3240 40588 3292 40594
rect 3240 40530 3292 40536
rect 3332 40588 3384 40594
rect 3332 40530 3384 40536
rect 3252 39642 3280 40530
rect 3240 39636 3292 39642
rect 3240 39578 3292 39584
rect 3344 39574 3372 40530
rect 3424 39976 3476 39982
rect 3424 39918 3476 39924
rect 3148 39568 3200 39574
rect 3148 39510 3200 39516
rect 3332 39568 3384 39574
rect 3332 39510 3384 39516
rect 3160 38418 3188 39510
rect 3436 39506 3464 39918
rect 3424 39500 3476 39506
rect 3424 39442 3476 39448
rect 3528 38826 3556 40938
rect 3608 40928 3660 40934
rect 3608 40870 3660 40876
rect 3620 39828 3648 40870
rect 3712 40662 3740 41618
rect 3976 41132 4028 41138
rect 3976 41074 4028 41080
rect 3792 40996 3844 41002
rect 3792 40938 3844 40944
rect 3700 40656 3752 40662
rect 3700 40598 3752 40604
rect 3804 40594 3832 40938
rect 3988 40730 4016 41074
rect 3976 40724 4028 40730
rect 3976 40666 4028 40672
rect 3792 40588 3844 40594
rect 3792 40530 3844 40536
rect 3988 40066 4016 40666
rect 4068 40520 4120 40526
rect 4068 40462 4120 40468
rect 4080 40186 4108 40462
rect 4068 40180 4120 40186
rect 4068 40122 4120 40128
rect 3712 40038 4016 40066
rect 3712 39982 3740 40038
rect 3988 39982 4016 40038
rect 4068 40044 4120 40050
rect 4068 39986 4120 39992
rect 3700 39976 3752 39982
rect 3700 39918 3752 39924
rect 3884 39976 3936 39982
rect 3884 39918 3936 39924
rect 3976 39976 4028 39982
rect 3976 39918 4028 39924
rect 3620 39800 3740 39828
rect 3516 38820 3568 38826
rect 3516 38762 3568 38768
rect 3148 38412 3200 38418
rect 3148 38354 3200 38360
rect 3160 37806 3188 38354
rect 3148 37800 3200 37806
rect 3148 37742 3200 37748
rect 3160 37466 3188 37742
rect 3516 37664 3568 37670
rect 3516 37606 3568 37612
rect 3148 37460 3200 37466
rect 3148 37402 3200 37408
rect 3240 36848 3292 36854
rect 3240 36790 3292 36796
rect 3148 36576 3200 36582
rect 3148 36518 3200 36524
rect 3056 35760 3108 35766
rect 3056 35702 3108 35708
rect 3068 35222 3096 35702
rect 3160 35630 3188 36518
rect 3148 35624 3200 35630
rect 3148 35566 3200 35572
rect 3056 35216 3108 35222
rect 3056 35158 3108 35164
rect 3252 34678 3280 36790
rect 3332 36304 3384 36310
rect 3332 36246 3384 36252
rect 3344 35154 3372 36246
rect 3424 36100 3476 36106
rect 3424 36042 3476 36048
rect 3332 35148 3384 35154
rect 3332 35090 3384 35096
rect 3240 34672 3292 34678
rect 3240 34614 3292 34620
rect 3332 34060 3384 34066
rect 3332 34002 3384 34008
rect 3056 33856 3108 33862
rect 3056 33798 3108 33804
rect 3068 33454 3096 33798
rect 3148 33516 3200 33522
rect 3148 33458 3200 33464
rect 3056 33448 3108 33454
rect 3056 33390 3108 33396
rect 3056 32768 3108 32774
rect 3056 32710 3108 32716
rect 2884 31726 3004 31754
rect 2780 31476 2832 31482
rect 2780 31418 2832 31424
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2700 29170 2728 30194
rect 2792 29782 2820 31418
rect 2780 29776 2832 29782
rect 2780 29718 2832 29724
rect 2688 29164 2740 29170
rect 2688 29106 2740 29112
rect 2688 28960 2740 28966
rect 2688 28902 2740 28908
rect 2700 28082 2728 28902
rect 2688 28076 2740 28082
rect 2688 28018 2740 28024
rect 2700 27674 2728 28018
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 2792 27878 2820 27950
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2688 27668 2740 27674
rect 2688 27610 2740 27616
rect 2792 27606 2820 27814
rect 2780 27600 2832 27606
rect 2780 27542 2832 27548
rect 2608 26846 2728 26874
rect 2596 26784 2648 26790
rect 2596 26726 2648 26732
rect 2608 26450 2636 26726
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 2504 26308 2556 26314
rect 2504 26250 2556 26256
rect 2516 25838 2544 26250
rect 2504 25832 2556 25838
rect 2504 25774 2556 25780
rect 2504 24676 2556 24682
rect 2504 24618 2556 24624
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2516 24410 2544 24618
rect 2504 24404 2556 24410
rect 2504 24346 2556 24352
rect 2608 24290 2636 26386
rect 2516 24262 2636 24290
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2424 22574 2452 23258
rect 2412 22568 2464 22574
rect 2412 22510 2464 22516
rect 2332 22066 2452 22094
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2332 21570 2360 21830
rect 2424 21690 2452 22066
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2332 21542 2452 21570
rect 2516 21554 2544 24262
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2608 22778 2636 23122
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2096 21440 2176 21468
rect 2044 21422 2096 21428
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2056 19310 2084 20334
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2056 18834 2084 19246
rect 2148 18902 2176 21440
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 2240 18970 2268 21422
rect 2424 21418 2452 21542
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2412 21412 2464 21418
rect 2412 21354 2464 21360
rect 2424 21010 2452 21354
rect 2700 21078 2728 26846
rect 2792 26790 2820 27542
rect 2780 26784 2832 26790
rect 2780 26726 2832 26732
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2792 24818 2820 25774
rect 2884 25362 2912 31726
rect 2964 31680 3016 31686
rect 2964 31622 3016 31628
rect 2976 31278 3004 31622
rect 3068 31278 3096 32710
rect 3160 32366 3188 33458
rect 3344 33386 3372 34002
rect 3436 33862 3464 36042
rect 3528 35034 3556 37606
rect 3608 35488 3660 35494
rect 3608 35430 3660 35436
rect 3620 35154 3648 35430
rect 3608 35148 3660 35154
rect 3608 35090 3660 35096
rect 3528 35006 3648 35034
rect 3516 34944 3568 34950
rect 3516 34886 3568 34892
rect 3424 33856 3476 33862
rect 3424 33798 3476 33804
rect 3528 33674 3556 34886
rect 3436 33646 3556 33674
rect 3332 33380 3384 33386
rect 3332 33322 3384 33328
rect 3240 33312 3292 33318
rect 3240 33254 3292 33260
rect 3252 32434 3280 33254
rect 3344 32570 3372 33322
rect 3332 32564 3384 32570
rect 3332 32506 3384 32512
rect 3240 32428 3292 32434
rect 3240 32370 3292 32376
rect 3332 32428 3384 32434
rect 3332 32370 3384 32376
rect 3148 32360 3200 32366
rect 3148 32302 3200 32308
rect 3160 31958 3188 32302
rect 3148 31952 3200 31958
rect 3148 31894 3200 31900
rect 3344 31822 3372 32370
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 3436 31498 3464 33646
rect 3516 32972 3568 32978
rect 3516 32914 3568 32920
rect 3528 32502 3556 32914
rect 3620 32842 3648 35006
rect 3712 34950 3740 39800
rect 3896 39506 3924 39918
rect 3884 39500 3936 39506
rect 3884 39442 3936 39448
rect 4080 39302 4108 39986
rect 3792 39296 3844 39302
rect 3792 39238 3844 39244
rect 4068 39296 4120 39302
rect 4068 39238 4120 39244
rect 3804 38894 3832 39238
rect 4172 38894 4200 42502
rect 4264 39642 4292 42502
rect 5000 42362 5028 45766
rect 5632 43444 5684 43450
rect 5632 43386 5684 43392
rect 5644 43110 5672 43386
rect 5632 43104 5684 43110
rect 5632 43046 5684 43052
rect 5172 42696 5224 42702
rect 5172 42638 5224 42644
rect 4988 42356 5040 42362
rect 4988 42298 5040 42304
rect 4804 42016 4856 42022
rect 4804 41958 4856 41964
rect 4528 41676 4580 41682
rect 4528 41618 4580 41624
rect 4344 41268 4396 41274
rect 4344 41210 4396 41216
rect 4436 41268 4488 41274
rect 4436 41210 4488 41216
rect 4356 40118 4384 41210
rect 4448 41070 4476 41210
rect 4436 41064 4488 41070
rect 4436 41006 4488 41012
rect 4344 40112 4396 40118
rect 4344 40054 4396 40060
rect 4344 39976 4396 39982
rect 4344 39918 4396 39924
rect 4252 39636 4304 39642
rect 4252 39578 4304 39584
rect 4356 39574 4384 39918
rect 4344 39568 4396 39574
rect 4344 39510 4396 39516
rect 4252 39432 4304 39438
rect 4252 39374 4304 39380
rect 3792 38888 3844 38894
rect 3792 38830 3844 38836
rect 4160 38888 4212 38894
rect 4160 38830 4212 38836
rect 4264 38486 4292 39374
rect 4356 38554 4384 39510
rect 4344 38548 4396 38554
rect 4344 38490 4396 38496
rect 4252 38480 4304 38486
rect 4252 38422 4304 38428
rect 3884 38412 3936 38418
rect 3884 38354 3936 38360
rect 3896 37942 3924 38354
rect 4160 38208 4212 38214
rect 4160 38150 4212 38156
rect 3884 37936 3936 37942
rect 3884 37878 3936 37884
rect 4172 37806 4200 38150
rect 4264 37874 4292 38422
rect 4448 38282 4476 41006
rect 4540 40050 4568 41618
rect 4816 40594 4844 41958
rect 5000 41414 5028 42298
rect 4908 41386 5028 41414
rect 4804 40588 4856 40594
rect 4804 40530 4856 40536
rect 4528 40044 4580 40050
rect 4528 39986 4580 39992
rect 4528 39636 4580 39642
rect 4528 39578 4580 39584
rect 4436 38276 4488 38282
rect 4436 38218 4488 38224
rect 4252 37868 4304 37874
rect 4252 37810 4304 37816
rect 4160 37800 4212 37806
rect 4160 37742 4212 37748
rect 3792 37664 3844 37670
rect 3792 37606 3844 37612
rect 3804 37398 3832 37606
rect 3792 37392 3844 37398
rect 3792 37334 3844 37340
rect 3884 37324 3936 37330
rect 3884 37266 3936 37272
rect 3896 36310 3924 37266
rect 3976 36712 4028 36718
rect 3976 36654 4028 36660
rect 3884 36304 3936 36310
rect 3884 36246 3936 36252
rect 3988 36242 4016 36654
rect 3976 36236 4028 36242
rect 3976 36178 4028 36184
rect 3792 36032 3844 36038
rect 3792 35974 3844 35980
rect 3700 34944 3752 34950
rect 3700 34886 3752 34892
rect 3608 32836 3660 32842
rect 3608 32778 3660 32784
rect 3516 32496 3568 32502
rect 3516 32438 3568 32444
rect 3608 32292 3660 32298
rect 3608 32234 3660 32240
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 3160 31470 3464 31498
rect 2964 31272 3016 31278
rect 2964 31214 3016 31220
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 2976 30598 3004 31214
rect 2964 30592 3016 30598
rect 2964 30534 3016 30540
rect 3160 29510 3188 31470
rect 3424 31408 3476 31414
rect 3424 31350 3476 31356
rect 3240 31340 3292 31346
rect 3240 31282 3292 31288
rect 3252 29850 3280 31282
rect 3332 30796 3384 30802
rect 3332 30738 3384 30744
rect 3344 30258 3372 30738
rect 3332 30252 3384 30258
rect 3332 30194 3384 30200
rect 3240 29844 3292 29850
rect 3240 29786 3292 29792
rect 3240 29708 3292 29714
rect 3240 29650 3292 29656
rect 3056 29504 3108 29510
rect 3056 29446 3108 29452
rect 3148 29504 3200 29510
rect 3148 29446 3200 29452
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 2976 28014 3004 29174
rect 3068 28626 3096 29446
rect 3056 28620 3108 28626
rect 3056 28562 3108 28568
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2792 23526 2820 24550
rect 3160 23798 3188 29446
rect 3252 27878 3280 29650
rect 3344 29102 3372 30194
rect 3332 29096 3384 29102
rect 3332 29038 3384 29044
rect 3332 28620 3384 28626
rect 3332 28562 3384 28568
rect 3344 28150 3372 28562
rect 3332 28144 3384 28150
rect 3332 28086 3384 28092
rect 3240 27872 3292 27878
rect 3240 27814 3292 27820
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 3252 26790 3280 27406
rect 3344 26926 3372 27474
rect 3332 26920 3384 26926
rect 3332 26862 3384 26868
rect 3240 26784 3292 26790
rect 3240 26726 3292 26732
rect 3252 26382 3280 26726
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3436 25498 3464 31350
rect 3528 30802 3556 31962
rect 3620 31482 3648 32234
rect 3804 31906 3832 35974
rect 3988 35766 4016 36178
rect 4172 36038 4200 37742
rect 4264 36174 4292 37810
rect 4344 37800 4396 37806
rect 4344 37742 4396 37748
rect 4436 37800 4488 37806
rect 4436 37742 4488 37748
rect 4356 36854 4384 37742
rect 4344 36848 4396 36854
rect 4344 36790 4396 36796
rect 4448 36242 4476 37742
rect 4436 36236 4488 36242
rect 4436 36178 4488 36184
rect 4252 36168 4304 36174
rect 4252 36110 4304 36116
rect 4160 36032 4212 36038
rect 4160 35974 4212 35980
rect 3976 35760 4028 35766
rect 3976 35702 4028 35708
rect 4172 35630 4200 35974
rect 4264 35698 4292 36110
rect 4252 35692 4304 35698
rect 4252 35634 4304 35640
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4068 33856 4120 33862
rect 4068 33798 4120 33804
rect 3884 33312 3936 33318
rect 3884 33254 3936 33260
rect 3896 32978 3924 33254
rect 3884 32972 3936 32978
rect 3884 32914 3936 32920
rect 3884 32836 3936 32842
rect 3884 32778 3936 32784
rect 3712 31878 3832 31906
rect 3608 31476 3660 31482
rect 3608 31418 3660 31424
rect 3608 31136 3660 31142
rect 3608 31078 3660 31084
rect 3516 30796 3568 30802
rect 3516 30738 3568 30744
rect 3516 30184 3568 30190
rect 3516 30126 3568 30132
rect 3528 29170 3556 30126
rect 3620 29510 3648 31078
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3516 29164 3568 29170
rect 3516 29106 3568 29112
rect 3528 27538 3556 29106
rect 3608 29096 3660 29102
rect 3608 29038 3660 29044
rect 3620 27606 3648 29038
rect 3608 27600 3660 27606
rect 3608 27542 3660 27548
rect 3516 27532 3568 27538
rect 3516 27474 3568 27480
rect 3424 25492 3476 25498
rect 3424 25434 3476 25440
rect 3332 25424 3384 25430
rect 3332 25366 3384 25372
rect 3148 23792 3200 23798
rect 3148 23734 3200 23740
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2964 23520 3016 23526
rect 2964 23462 3016 23468
rect 2688 21072 2740 21078
rect 2688 21014 2740 21020
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2332 19310 2360 20742
rect 2424 20398 2452 20946
rect 2792 20874 2820 23462
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2976 20806 3004 23462
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 3252 22098 3280 23054
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 3344 21350 3372 25366
rect 3436 25158 3464 25434
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3528 24614 3556 27474
rect 3712 26908 3740 31878
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3804 30938 3832 31758
rect 3792 30932 3844 30938
rect 3792 30874 3844 30880
rect 3792 30184 3844 30190
rect 3792 30126 3844 30132
rect 3804 29306 3832 30126
rect 3792 29300 3844 29306
rect 3792 29242 3844 29248
rect 3792 28960 3844 28966
rect 3792 28902 3844 28908
rect 3804 28014 3832 28902
rect 3896 28762 3924 32778
rect 3976 32768 4028 32774
rect 3976 32710 4028 32716
rect 3988 32366 4016 32710
rect 3976 32360 4028 32366
rect 3976 32302 4028 32308
rect 4080 32178 4108 33798
rect 3988 32150 4108 32178
rect 3884 28756 3936 28762
rect 3884 28698 3936 28704
rect 3884 28552 3936 28558
rect 3884 28494 3936 28500
rect 3896 28218 3924 28494
rect 3884 28212 3936 28218
rect 3884 28154 3936 28160
rect 3792 28008 3844 28014
rect 3792 27950 3844 27956
rect 3884 27532 3936 27538
rect 3884 27474 3936 27480
rect 3792 27328 3844 27334
rect 3792 27270 3844 27276
rect 3620 26880 3740 26908
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3528 23866 3556 24550
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3620 22098 3648 26880
rect 3700 26784 3752 26790
rect 3700 26726 3752 26732
rect 3712 25226 3740 26726
rect 3700 25220 3752 25226
rect 3700 25162 3752 25168
rect 3712 24682 3740 25162
rect 3700 24676 3752 24682
rect 3700 24618 3752 24624
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3608 22092 3660 22098
rect 3608 22034 3660 22040
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 2688 20528 2740 20534
rect 2688 20470 2740 20476
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2424 19990 2452 20334
rect 2412 19984 2464 19990
rect 2412 19926 2464 19932
rect 2504 19916 2556 19922
rect 2504 19858 2556 19864
rect 2412 19440 2464 19446
rect 2412 19382 2464 19388
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2332 18902 2360 19246
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 1952 18760 2004 18766
rect 1952 18702 2004 18708
rect 1964 17882 1992 18702
rect 2056 18086 2084 18770
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2240 18222 2268 18566
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1964 17048 1992 17818
rect 1964 17020 2084 17048
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 16114 1992 16594
rect 2056 16590 2084 17020
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 16250 2084 16526
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 2148 14550 2176 16594
rect 2240 14958 2268 16594
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1780 13246 1900 13274
rect 1780 12442 1808 13246
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1780 11218 1808 12378
rect 1872 11762 1900 13126
rect 1964 12714 1992 13670
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 2056 12434 2084 14010
rect 2148 14006 2176 14486
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2240 13870 2268 14894
rect 2228 13864 2280 13870
rect 2148 13824 2228 13852
rect 2148 13190 2176 13824
rect 2228 13806 2280 13812
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 1964 12406 2084 12434
rect 2332 12434 2360 18702
rect 2424 15450 2452 19382
rect 2516 19334 2544 19858
rect 2700 19514 2728 20470
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 2976 20058 3004 20402
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3068 19938 3096 21286
rect 3436 21146 3464 22034
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 2976 19910 3096 19938
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 2507 19306 2544 19334
rect 2507 19258 2535 19306
rect 2507 19230 2553 19258
rect 2525 19122 2553 19230
rect 2688 19168 2740 19174
rect 2525 19116 2688 19122
rect 2525 19110 2740 19116
rect 2525 19094 2728 19110
rect 2700 18834 2728 19094
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2792 18766 2820 19382
rect 2884 19310 2912 19722
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2700 17746 2728 18158
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2608 16522 2636 16730
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 15570 2544 16390
rect 2608 16114 2636 16458
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2424 15422 2544 15450
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2424 14414 2452 14758
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 14074 2452 14350
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2424 13462 2452 13670
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2516 12434 2544 15422
rect 2608 14822 2636 16050
rect 2700 15638 2728 17682
rect 2792 16998 2820 18022
rect 2884 17542 2912 19246
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 12714 2636 14554
rect 2700 13394 2728 15574
rect 2792 14618 2820 16934
rect 2976 15706 3004 19910
rect 3160 19242 3188 20878
rect 3252 20398 3280 21014
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3344 20806 3372 20878
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18970 3096 19110
rect 3252 18970 3280 20334
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3436 19922 3464 20198
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 13870 2820 14418
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2700 12782 2728 13330
rect 2792 12986 2820 13806
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2332 12406 2452 12434
rect 2516 12406 2636 12434
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1872 11150 1900 11698
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1768 11076 1820 11082
rect 1768 11018 1820 11024
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1596 8452 1716 8480
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 6866 1624 8298
rect 1688 8022 1716 8452
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7410 1716 7686
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 5778 1624 6802
rect 1688 6186 1716 7142
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1688 5658 1716 6122
rect 1596 5630 1716 5658
rect 1596 2650 1624 5630
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1688 4282 1716 5102
rect 1780 5098 1808 11018
rect 1964 10962 1992 12406
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 1872 10934 1992 10962
rect 1768 5092 1820 5098
rect 1768 5034 1820 5040
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1872 4146 1900 10934
rect 2056 10266 2084 11562
rect 2332 11218 2360 11630
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2332 10282 2360 11154
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2240 10254 2360 10282
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 7002 1992 7686
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1964 6390 1992 6802
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2056 2774 2084 8978
rect 2148 8566 2176 9862
rect 2240 9382 2268 10254
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9042 2268 9318
rect 2424 9178 2452 12406
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 9518 2544 11494
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2228 8832 2280 8838
rect 2280 8780 2360 8786
rect 2228 8774 2360 8780
rect 2240 8758 2360 8774
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 8294 2268 8366
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2228 7951 2280 7957
rect 2228 7893 2280 7899
rect 2240 5846 2268 7893
rect 2332 7410 2360 8758
rect 2424 8090 2452 9114
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2148 4826 2176 5578
rect 2332 5030 2360 7346
rect 2424 7342 2452 8026
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2424 5914 2452 6870
rect 2516 6798 2544 8434
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2516 5778 2544 6598
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2056 2746 2176 2774
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2148 2106 2176 2746
rect 1492 2100 1544 2106
rect 1492 2042 1544 2048
rect 2136 2100 2188 2106
rect 2136 2042 2188 2048
rect 2608 2038 2636 12406
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2700 10810 2728 12242
rect 2792 11830 2820 12922
rect 2884 12918 2912 14486
rect 2964 14000 3016 14006
rect 2964 13942 3016 13948
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2976 11898 3004 13942
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2792 11218 2820 11766
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2884 11286 2912 11698
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2976 11354 3004 11630
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2884 11150 2912 11222
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2884 10674 2912 11086
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2700 8498 2728 10202
rect 2976 10198 3004 10950
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 7954 2728 8434
rect 2792 8430 2820 8978
rect 2780 8424 2832 8430
rect 3068 8378 3096 17070
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3160 16658 3188 17002
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3160 10674 3188 15914
rect 3252 14890 3280 18770
rect 3344 18698 3372 19654
rect 3436 19446 3464 19858
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 3436 16998 3464 19246
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3252 11218 3280 14554
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3344 13326 3372 13874
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 11762 3372 13262
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10130 3188 10610
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3344 9722 3372 11290
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 2780 8366 2832 8372
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2700 7342 2728 7754
rect 2792 7750 2820 8366
rect 2884 8350 3096 8378
rect 3240 8356 3292 8362
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2700 6866 2728 7278
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6458 2728 6802
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2792 5914 2820 7210
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2884 5250 2912 8350
rect 3240 8298 3292 8304
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2976 6866 3004 7822
rect 3068 7410 3096 8230
rect 3252 7954 3280 8298
rect 3436 8072 3464 16730
rect 3344 8044 3464 8072
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7478 3188 7822
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3068 6798 3096 7346
rect 3344 7290 3372 8044
rect 3528 7970 3556 20946
rect 3620 19922 3648 21422
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3620 19514 3648 19858
rect 3608 19508 3660 19514
rect 3608 19450 3660 19456
rect 3620 18834 3648 19450
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3620 12442 3648 17138
rect 3712 16794 3740 24618
rect 3804 21486 3832 27270
rect 3896 26926 3924 27474
rect 3884 26920 3936 26926
rect 3884 26862 3936 26868
rect 3896 26586 3924 26862
rect 3884 26580 3936 26586
rect 3884 26522 3936 26528
rect 3792 21480 3844 21486
rect 3792 21422 3844 21428
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3792 21072 3844 21078
rect 3792 21014 3844 21020
rect 3804 19174 3832 21014
rect 3896 20942 3924 21286
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3896 20806 3924 20878
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 3896 18834 3924 19314
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3896 17882 3924 18770
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3884 17604 3936 17610
rect 3884 17546 3936 17552
rect 3896 17082 3924 17546
rect 3988 17202 4016 32150
rect 4172 32042 4200 35430
rect 4264 34542 4292 35634
rect 4448 35630 4476 36178
rect 4436 35624 4488 35630
rect 4436 35566 4488 35572
rect 4252 34536 4304 34542
rect 4252 34478 4304 34484
rect 4540 33658 4568 39578
rect 4620 38820 4672 38826
rect 4620 38762 4672 38768
rect 4528 33652 4580 33658
rect 4528 33594 4580 33600
rect 4252 33584 4304 33590
rect 4252 33526 4304 33532
rect 4080 32014 4200 32042
rect 4080 31414 4108 32014
rect 4264 31940 4292 33526
rect 4344 32768 4396 32774
rect 4344 32710 4396 32716
rect 4356 32230 4384 32710
rect 4528 32360 4580 32366
rect 4528 32302 4580 32308
rect 4344 32224 4396 32230
rect 4344 32166 4396 32172
rect 4172 31912 4292 31940
rect 4172 31686 4200 31912
rect 4252 31816 4304 31822
rect 4252 31758 4304 31764
rect 4160 31680 4212 31686
rect 4160 31622 4212 31628
rect 4172 31482 4200 31622
rect 4160 31476 4212 31482
rect 4160 31418 4212 31424
rect 4068 31408 4120 31414
rect 4068 31350 4120 31356
rect 4264 31210 4292 31758
rect 4252 31204 4304 31210
rect 4252 31146 4304 31152
rect 4356 30802 4384 32166
rect 4436 31952 4488 31958
rect 4436 31894 4488 31900
rect 4448 31346 4476 31894
rect 4436 31340 4488 31346
rect 4436 31282 4488 31288
rect 4436 30864 4488 30870
rect 4436 30806 4488 30812
rect 4068 30796 4120 30802
rect 4068 30738 4120 30744
rect 4160 30796 4212 30802
rect 4160 30738 4212 30744
rect 4344 30796 4396 30802
rect 4344 30738 4396 30744
rect 4080 29714 4108 30738
rect 4172 30054 4200 30738
rect 4252 30728 4304 30734
rect 4252 30670 4304 30676
rect 4264 30326 4292 30670
rect 4344 30388 4396 30394
rect 4344 30330 4396 30336
rect 4252 30320 4304 30326
rect 4252 30262 4304 30268
rect 4160 30048 4212 30054
rect 4160 29990 4212 29996
rect 4068 29708 4120 29714
rect 4068 29650 4120 29656
rect 4068 29572 4120 29578
rect 4068 29514 4120 29520
rect 4080 29102 4108 29514
rect 4172 29186 4200 29990
rect 4356 29850 4384 30330
rect 4344 29844 4396 29850
rect 4344 29786 4396 29792
rect 4252 29708 4304 29714
rect 4252 29650 4304 29656
rect 4264 29306 4292 29650
rect 4344 29640 4396 29646
rect 4344 29582 4396 29588
rect 4252 29300 4304 29306
rect 4252 29242 4304 29248
rect 4172 29158 4292 29186
rect 4356 29170 4384 29582
rect 4448 29306 4476 30806
rect 4540 30258 4568 32302
rect 4528 30252 4580 30258
rect 4528 30194 4580 30200
rect 4436 29300 4488 29306
rect 4436 29242 4488 29248
rect 4068 29096 4120 29102
rect 4068 29038 4120 29044
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 4080 27062 4108 28698
rect 4172 28694 4200 28902
rect 4160 28688 4212 28694
rect 4160 28630 4212 28636
rect 4264 28642 4292 29158
rect 4344 29164 4396 29170
rect 4344 29106 4396 29112
rect 4356 28762 4384 29106
rect 4344 28756 4396 28762
rect 4344 28698 4396 28704
rect 4264 28614 4384 28642
rect 4160 28416 4212 28422
rect 4160 28358 4212 28364
rect 4172 28150 4200 28358
rect 4160 28144 4212 28150
rect 4160 28086 4212 28092
rect 4252 27940 4304 27946
rect 4252 27882 4304 27888
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4172 26926 4200 27406
rect 4264 27130 4292 27882
rect 4356 27470 4384 28614
rect 4436 28076 4488 28082
rect 4436 28018 4488 28024
rect 4344 27464 4396 27470
rect 4344 27406 4396 27412
rect 4252 27124 4304 27130
rect 4252 27066 4304 27072
rect 4160 26920 4212 26926
rect 4344 26920 4396 26926
rect 4160 26862 4212 26868
rect 4264 26880 4344 26908
rect 4068 26784 4120 26790
rect 4068 26726 4120 26732
rect 4080 25770 4108 26726
rect 4172 26518 4200 26862
rect 4160 26512 4212 26518
rect 4160 26454 4212 26460
rect 4068 25764 4120 25770
rect 4068 25706 4120 25712
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4080 22098 4108 25434
rect 4172 24750 4200 26454
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4172 24342 4200 24686
rect 4160 24336 4212 24342
rect 4160 24278 4212 24284
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4172 22438 4200 24142
rect 4264 24138 4292 26880
rect 4344 26862 4396 26868
rect 4344 25152 4396 25158
rect 4344 25094 4396 25100
rect 4356 24886 4384 25094
rect 4344 24880 4396 24886
rect 4344 24822 4396 24828
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 4264 22574 4292 22918
rect 4252 22568 4304 22574
rect 4252 22510 4304 22516
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4080 18426 4108 20878
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4172 19922 4200 20742
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4264 20058 4292 20334
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4264 18834 4292 19314
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4080 18086 4108 18362
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4080 17270 4108 18022
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3896 17054 4016 17082
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3712 15638 3740 16390
rect 3700 15632 3752 15638
rect 3700 15574 3752 15580
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3620 11150 3648 12378
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3252 7262 3372 7290
rect 3436 7942 3556 7970
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6186 3004 6666
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2976 5778 3004 6122
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2976 5370 3004 5714
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2884 5222 3004 5250
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2700 4826 2728 4966
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2884 3738 2912 4218
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2884 3194 2912 3674
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2596 2032 2648 2038
rect 2596 1974 2648 1980
rect 1860 1420 1912 1426
rect 1860 1362 1912 1368
rect 1872 1018 1900 1362
rect 1860 1012 1912 1018
rect 1860 954 1912 960
rect 2792 800 2820 3062
rect 2976 1358 3004 5222
rect 3068 4826 3096 6394
rect 3160 5642 3188 6734
rect 3252 5914 3280 7262
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 2650 3188 4626
rect 3252 2650 3280 4694
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3344 2106 3372 6802
rect 3436 2106 3464 7942
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3528 7546 3556 7822
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3528 7002 3556 7278
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3620 6866 3648 10746
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3712 4826 3740 15574
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3804 14822 3832 15506
rect 3896 15434 3924 16934
rect 3884 15428 3936 15434
rect 3884 15370 3936 15376
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 12442 3832 14758
rect 3896 14414 3924 15370
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3896 14006 3924 14350
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3896 13734 3924 13806
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3884 13456 3936 13462
rect 3988 13444 4016 17054
rect 4080 16454 4108 17206
rect 4264 17116 4292 18022
rect 4356 17218 4384 24822
rect 4448 23322 4476 28018
rect 4540 27878 4568 30194
rect 4528 27872 4580 27878
rect 4528 27814 4580 27820
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4540 26518 4568 27270
rect 4528 26512 4580 26518
rect 4528 26454 4580 26460
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4540 23662 4568 24550
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4632 22574 4660 38762
rect 4712 38208 4764 38214
rect 4712 38150 4764 38156
rect 4724 37330 4752 38150
rect 4712 37324 4764 37330
rect 4712 37266 4764 37272
rect 4712 36304 4764 36310
rect 4712 36246 4764 36252
rect 4724 35562 4752 36246
rect 4712 35556 4764 35562
rect 4712 35498 4764 35504
rect 4724 35018 4752 35498
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4712 34536 4764 34542
rect 4712 34478 4764 34484
rect 4724 33862 4752 34478
rect 4712 33856 4764 33862
rect 4712 33798 4764 33804
rect 4724 31822 4752 33798
rect 4712 31816 4764 31822
rect 4712 31758 4764 31764
rect 4712 31680 4764 31686
rect 4712 31622 4764 31628
rect 4724 28558 4752 31622
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4724 27402 4752 28494
rect 4816 28422 4844 40530
rect 4908 38282 4936 41386
rect 5080 41064 5132 41070
rect 5080 41006 5132 41012
rect 5092 40594 5120 41006
rect 5080 40588 5132 40594
rect 5080 40530 5132 40536
rect 4988 40112 5040 40118
rect 4988 40054 5040 40060
rect 5000 39982 5028 40054
rect 4988 39976 5040 39982
rect 4988 39918 5040 39924
rect 5000 39506 5028 39918
rect 5092 39574 5120 40530
rect 5080 39568 5132 39574
rect 5080 39510 5132 39516
rect 4988 39500 5040 39506
rect 4988 39442 5040 39448
rect 4988 39364 5040 39370
rect 4988 39306 5040 39312
rect 4896 38276 4948 38282
rect 4896 38218 4948 38224
rect 5000 37670 5028 39306
rect 4988 37664 5040 37670
rect 4988 37606 5040 37612
rect 5184 37274 5212 42638
rect 5644 42226 5672 43046
rect 5736 42770 5764 47942
rect 6102 47900 6410 47920
rect 6102 47898 6108 47900
rect 6164 47898 6188 47900
rect 6244 47898 6268 47900
rect 6324 47898 6348 47900
rect 6404 47898 6410 47900
rect 6164 47846 6166 47898
rect 6346 47846 6348 47898
rect 6102 47844 6108 47846
rect 6164 47844 6188 47846
rect 6244 47844 6268 47846
rect 6324 47844 6348 47846
rect 6404 47844 6410 47846
rect 6102 47824 6410 47844
rect 8024 47524 8076 47530
rect 8024 47466 8076 47472
rect 6920 47456 6972 47462
rect 6920 47398 6972 47404
rect 6102 46812 6410 46832
rect 6102 46810 6108 46812
rect 6164 46810 6188 46812
rect 6244 46810 6268 46812
rect 6324 46810 6348 46812
rect 6404 46810 6410 46812
rect 6164 46758 6166 46810
rect 6346 46758 6348 46810
rect 6102 46756 6108 46758
rect 6164 46756 6188 46758
rect 6244 46756 6268 46758
rect 6324 46756 6348 46758
rect 6404 46756 6410 46758
rect 6102 46736 6410 46756
rect 6932 46578 6960 47398
rect 7748 47116 7800 47122
rect 7748 47058 7800 47064
rect 7840 47116 7892 47122
rect 7840 47058 7892 47064
rect 6920 46572 6972 46578
rect 6920 46514 6972 46520
rect 6102 45724 6410 45744
rect 6102 45722 6108 45724
rect 6164 45722 6188 45724
rect 6244 45722 6268 45724
rect 6324 45722 6348 45724
rect 6404 45722 6410 45724
rect 6164 45670 6166 45722
rect 6346 45670 6348 45722
rect 6102 45668 6108 45670
rect 6164 45668 6188 45670
rect 6244 45668 6268 45670
rect 6324 45668 6348 45670
rect 6404 45668 6410 45670
rect 6102 45648 6410 45668
rect 6932 45422 6960 46514
rect 7288 46504 7340 46510
rect 7288 46446 7340 46452
rect 7196 46028 7248 46034
rect 7196 45970 7248 45976
rect 6920 45416 6972 45422
rect 6920 45358 6972 45364
rect 7208 45082 7236 45970
rect 7300 45422 7328 46446
rect 7564 46436 7616 46442
rect 7564 46378 7616 46384
rect 7472 45892 7524 45898
rect 7472 45834 7524 45840
rect 7484 45422 7512 45834
rect 7576 45490 7604 46378
rect 7760 46102 7788 47058
rect 7852 46714 7880 47058
rect 7840 46708 7892 46714
rect 7840 46650 7892 46656
rect 7840 46504 7892 46510
rect 7840 46446 7892 46452
rect 7748 46096 7800 46102
rect 7748 46038 7800 46044
rect 7564 45484 7616 45490
rect 7564 45426 7616 45432
rect 7288 45416 7340 45422
rect 7288 45358 7340 45364
rect 7472 45416 7524 45422
rect 7472 45358 7524 45364
rect 7196 45076 7248 45082
rect 7196 45018 7248 45024
rect 7300 45014 7328 45358
rect 7380 45348 7432 45354
rect 7380 45290 7432 45296
rect 7288 45008 7340 45014
rect 7288 44950 7340 44956
rect 7196 44872 7248 44878
rect 7392 44860 7420 45290
rect 7484 44946 7512 45358
rect 7576 45098 7604 45426
rect 7852 45422 7880 46446
rect 8036 45558 8064 47466
rect 8392 45824 8444 45830
rect 8392 45766 8444 45772
rect 8024 45552 8076 45558
rect 8024 45494 8076 45500
rect 7840 45416 7892 45422
rect 7840 45358 7892 45364
rect 8024 45280 8076 45286
rect 8024 45222 8076 45228
rect 7576 45070 7696 45098
rect 7564 45008 7616 45014
rect 7564 44950 7616 44956
rect 7472 44940 7524 44946
rect 7472 44882 7524 44888
rect 7248 44832 7420 44860
rect 7196 44814 7248 44820
rect 6102 44636 6410 44656
rect 6102 44634 6108 44636
rect 6164 44634 6188 44636
rect 6244 44634 6268 44636
rect 6324 44634 6348 44636
rect 6404 44634 6410 44636
rect 6164 44582 6166 44634
rect 6346 44582 6348 44634
rect 6102 44580 6108 44582
rect 6164 44580 6188 44582
rect 6244 44580 6268 44582
rect 6324 44580 6348 44582
rect 6404 44580 6410 44582
rect 6102 44560 6410 44580
rect 7012 44464 7064 44470
rect 7012 44406 7064 44412
rect 5816 44328 5868 44334
rect 5816 44270 5868 44276
rect 5828 43314 5856 44270
rect 6828 44260 6880 44266
rect 6828 44202 6880 44208
rect 6840 43994 6868 44202
rect 6828 43988 6880 43994
rect 6828 43930 6880 43936
rect 7024 43858 7052 44406
rect 7012 43852 7064 43858
rect 7012 43794 7064 43800
rect 6736 43648 6788 43654
rect 6736 43590 6788 43596
rect 6102 43548 6410 43568
rect 6102 43546 6108 43548
rect 6164 43546 6188 43548
rect 6244 43546 6268 43548
rect 6324 43546 6348 43548
rect 6404 43546 6410 43548
rect 6164 43494 6166 43546
rect 6346 43494 6348 43546
rect 6102 43492 6108 43494
rect 6164 43492 6188 43494
rect 6244 43492 6268 43494
rect 6324 43492 6348 43494
rect 6404 43492 6410 43494
rect 6102 43472 6410 43492
rect 5816 43308 5868 43314
rect 5816 43250 5868 43256
rect 5724 42764 5776 42770
rect 5724 42706 5776 42712
rect 5632 42220 5684 42226
rect 5632 42162 5684 42168
rect 5540 42152 5592 42158
rect 5540 42094 5592 42100
rect 5356 41608 5408 41614
rect 5356 41550 5408 41556
rect 5264 40384 5316 40390
rect 5264 40326 5316 40332
rect 5276 38350 5304 40326
rect 5368 39030 5396 41550
rect 5448 41064 5500 41070
rect 5448 41006 5500 41012
rect 5460 40662 5488 41006
rect 5448 40656 5500 40662
rect 5448 40598 5500 40604
rect 5552 40474 5580 42094
rect 5828 41750 5856 43250
rect 6102 42460 6410 42480
rect 6102 42458 6108 42460
rect 6164 42458 6188 42460
rect 6244 42458 6268 42460
rect 6324 42458 6348 42460
rect 6404 42458 6410 42460
rect 6164 42406 6166 42458
rect 6346 42406 6348 42458
rect 6102 42404 6108 42406
rect 6164 42404 6188 42406
rect 6244 42404 6268 42406
rect 6324 42404 6348 42406
rect 6404 42404 6410 42406
rect 6102 42384 6410 42404
rect 6644 42152 6696 42158
rect 6644 42094 6696 42100
rect 6552 42084 6604 42090
rect 6552 42026 6604 42032
rect 6000 42016 6052 42022
rect 6000 41958 6052 41964
rect 5816 41744 5868 41750
rect 5816 41686 5868 41692
rect 5632 41472 5684 41478
rect 5632 41414 5684 41420
rect 5644 40594 5672 41414
rect 5724 40928 5776 40934
rect 5724 40870 5776 40876
rect 5632 40588 5684 40594
rect 5632 40530 5684 40536
rect 5460 40446 5580 40474
rect 5356 39024 5408 39030
rect 5356 38966 5408 38972
rect 5264 38344 5316 38350
rect 5264 38286 5316 38292
rect 5356 38276 5408 38282
rect 5356 38218 5408 38224
rect 5368 38010 5396 38218
rect 5356 38004 5408 38010
rect 5356 37946 5408 37952
rect 5000 37246 5212 37274
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 4908 32910 4936 33254
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 5000 32842 5028 37246
rect 5276 36786 5304 37266
rect 5264 36780 5316 36786
rect 5264 36722 5316 36728
rect 5080 36644 5132 36650
rect 5080 36586 5132 36592
rect 5092 36378 5120 36586
rect 5080 36372 5132 36378
rect 5080 36314 5132 36320
rect 5172 36032 5224 36038
rect 5172 35974 5224 35980
rect 5080 35624 5132 35630
rect 5080 35566 5132 35572
rect 5092 35494 5120 35566
rect 5184 35562 5212 35974
rect 5368 35850 5396 37946
rect 5460 37274 5488 40446
rect 5540 40384 5592 40390
rect 5540 40326 5592 40332
rect 5552 38418 5580 40326
rect 5644 40050 5672 40530
rect 5632 40044 5684 40050
rect 5632 39986 5684 39992
rect 5632 39840 5684 39846
rect 5736 39828 5764 40870
rect 5684 39800 5764 39828
rect 5632 39782 5684 39788
rect 5644 38826 5672 39782
rect 5828 39098 5856 41686
rect 5908 40996 5960 41002
rect 5908 40938 5960 40944
rect 5816 39092 5868 39098
rect 5816 39034 5868 39040
rect 5632 38820 5684 38826
rect 5632 38762 5684 38768
rect 5828 38418 5856 39034
rect 5540 38412 5592 38418
rect 5540 38354 5592 38360
rect 5816 38412 5868 38418
rect 5816 38354 5868 38360
rect 5724 38344 5776 38350
rect 5724 38286 5776 38292
rect 5736 37466 5764 38286
rect 5920 37874 5948 40938
rect 5908 37868 5960 37874
rect 5908 37810 5960 37816
rect 5816 37664 5868 37670
rect 5816 37606 5868 37612
rect 5724 37460 5776 37466
rect 5724 37402 5776 37408
rect 5460 37246 5672 37274
rect 5540 36168 5592 36174
rect 5540 36110 5592 36116
rect 5368 35834 5488 35850
rect 5368 35828 5500 35834
rect 5368 35822 5448 35828
rect 5448 35770 5500 35776
rect 5172 35556 5224 35562
rect 5172 35498 5224 35504
rect 5080 35488 5132 35494
rect 5080 35430 5132 35436
rect 4988 32836 5040 32842
rect 4988 32778 5040 32784
rect 4896 32564 4948 32570
rect 4896 32506 4948 32512
rect 4908 30682 4936 32506
rect 5092 31906 5120 35430
rect 5264 35148 5316 35154
rect 5264 35090 5316 35096
rect 5276 34542 5304 35090
rect 5356 34944 5408 34950
rect 5356 34886 5408 34892
rect 5264 34536 5316 34542
rect 5264 34478 5316 34484
rect 5172 34468 5224 34474
rect 5172 34410 5224 34416
rect 5184 34066 5212 34410
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 5276 33590 5304 34478
rect 5368 34202 5396 34886
rect 5356 34196 5408 34202
rect 5356 34138 5408 34144
rect 5368 34066 5396 34138
rect 5460 34066 5488 35770
rect 5356 34060 5408 34066
rect 5356 34002 5408 34008
rect 5448 34060 5500 34066
rect 5448 34002 5500 34008
rect 5460 33810 5488 34002
rect 5368 33782 5488 33810
rect 5264 33584 5316 33590
rect 5264 33526 5316 33532
rect 5368 33436 5396 33782
rect 5448 33652 5500 33658
rect 5448 33594 5500 33600
rect 5184 33408 5396 33436
rect 5184 32570 5212 33408
rect 5460 32910 5488 33594
rect 5552 32978 5580 36110
rect 5644 34388 5672 37246
rect 5736 35698 5764 37402
rect 5724 35692 5776 35698
rect 5724 35634 5776 35640
rect 5736 35154 5764 35634
rect 5828 35290 5856 37606
rect 5908 35692 5960 35698
rect 5908 35634 5960 35640
rect 5816 35284 5868 35290
rect 5816 35226 5868 35232
rect 5724 35148 5776 35154
rect 5724 35090 5776 35096
rect 5736 34542 5764 35090
rect 5816 34944 5868 34950
rect 5816 34886 5868 34892
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 5724 34400 5776 34406
rect 5644 34360 5724 34388
rect 5724 34342 5776 34348
rect 5632 33856 5684 33862
rect 5632 33798 5684 33804
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5448 32904 5500 32910
rect 5448 32846 5500 32852
rect 5356 32768 5408 32774
rect 5356 32710 5408 32716
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5264 32496 5316 32502
rect 5264 32438 5316 32444
rect 5172 32224 5224 32230
rect 5172 32166 5224 32172
rect 5184 32026 5212 32166
rect 5172 32020 5224 32026
rect 5172 31962 5224 31968
rect 5092 31878 5212 31906
rect 4988 31680 5040 31686
rect 4988 31622 5040 31628
rect 5000 30802 5028 31622
rect 5080 31272 5132 31278
rect 5080 31214 5132 31220
rect 5092 30938 5120 31214
rect 5080 30932 5132 30938
rect 5080 30874 5132 30880
rect 4988 30796 5040 30802
rect 4988 30738 5040 30744
rect 5080 30728 5132 30734
rect 4908 30654 5028 30682
rect 5080 30670 5132 30676
rect 4896 30116 4948 30122
rect 4896 30058 4948 30064
rect 4804 28416 4856 28422
rect 4804 28358 4856 28364
rect 4908 28218 4936 30058
rect 5000 29238 5028 30654
rect 5092 30598 5120 30670
rect 5080 30592 5132 30598
rect 5080 30534 5132 30540
rect 4988 29232 5040 29238
rect 4988 29174 5040 29180
rect 5000 28694 5028 29174
rect 4988 28688 5040 28694
rect 4988 28630 5040 28636
rect 4896 28212 4948 28218
rect 4896 28154 4948 28160
rect 4988 28212 5040 28218
rect 4988 28154 5040 28160
rect 5000 28098 5028 28154
rect 4816 28082 5028 28098
rect 4804 28076 5028 28082
rect 4856 28070 5028 28076
rect 4804 28018 4856 28024
rect 4896 28008 4948 28014
rect 4896 27950 4948 27956
rect 4804 27872 4856 27878
rect 4804 27814 4856 27820
rect 4712 27396 4764 27402
rect 4712 27338 4764 27344
rect 4712 27056 4764 27062
rect 4712 26998 4764 27004
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 4448 21894 4476 21966
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4448 21486 4476 21830
rect 4724 21690 4752 26998
rect 4816 26926 4844 27814
rect 4908 27538 4936 27950
rect 5092 27614 5120 30534
rect 5000 27586 5120 27614
rect 4896 27532 4948 27538
rect 4896 27474 4948 27480
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4816 25838 4844 26318
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4816 24818 4844 25774
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4816 24342 4844 24754
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4436 21480 4488 21486
rect 4436 21422 4488 21428
rect 4632 21350 4660 21626
rect 4620 21344 4672 21350
rect 4724 21332 4752 21626
rect 4816 21554 4844 22374
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4908 21418 4936 27270
rect 5000 26858 5028 27586
rect 5184 27010 5212 31878
rect 5276 30054 5304 32438
rect 5368 32366 5396 32710
rect 5356 32360 5408 32366
rect 5356 32302 5408 32308
rect 5356 31884 5408 31890
rect 5356 31826 5408 31832
rect 5368 30326 5396 31826
rect 5460 31822 5488 32846
rect 5552 32298 5580 32914
rect 5644 32910 5672 33798
rect 5736 33590 5764 34342
rect 5828 33998 5856 34886
rect 5816 33992 5868 33998
rect 5816 33934 5868 33940
rect 5724 33584 5776 33590
rect 5724 33526 5776 33532
rect 5828 33454 5856 33934
rect 5816 33448 5868 33454
rect 5816 33390 5868 33396
rect 5724 33380 5776 33386
rect 5724 33322 5776 33328
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5540 32292 5592 32298
rect 5540 32234 5592 32240
rect 5736 31958 5764 33322
rect 5920 33300 5948 35634
rect 6012 33658 6040 41958
rect 6102 41372 6410 41392
rect 6102 41370 6108 41372
rect 6164 41370 6188 41372
rect 6244 41370 6268 41372
rect 6324 41370 6348 41372
rect 6404 41370 6410 41372
rect 6164 41318 6166 41370
rect 6346 41318 6348 41370
rect 6102 41316 6108 41318
rect 6164 41316 6188 41318
rect 6244 41316 6268 41318
rect 6324 41316 6348 41318
rect 6404 41316 6410 41318
rect 6102 41296 6410 41316
rect 6102 40284 6410 40304
rect 6102 40282 6108 40284
rect 6164 40282 6188 40284
rect 6244 40282 6268 40284
rect 6324 40282 6348 40284
rect 6404 40282 6410 40284
rect 6164 40230 6166 40282
rect 6346 40230 6348 40282
rect 6102 40228 6108 40230
rect 6164 40228 6188 40230
rect 6244 40228 6268 40230
rect 6324 40228 6348 40230
rect 6404 40228 6410 40230
rect 6102 40208 6410 40228
rect 6368 39840 6420 39846
rect 6368 39782 6420 39788
rect 6380 39574 6408 39782
rect 6368 39568 6420 39574
rect 6368 39510 6420 39516
rect 6460 39432 6512 39438
rect 6460 39374 6512 39380
rect 6102 39196 6410 39216
rect 6102 39194 6108 39196
rect 6164 39194 6188 39196
rect 6244 39194 6268 39196
rect 6324 39194 6348 39196
rect 6404 39194 6410 39196
rect 6164 39142 6166 39194
rect 6346 39142 6348 39194
rect 6102 39140 6108 39142
rect 6164 39140 6188 39142
rect 6244 39140 6268 39142
rect 6324 39140 6348 39142
rect 6404 39140 6410 39142
rect 6102 39120 6410 39140
rect 6472 39098 6500 39374
rect 6460 39092 6512 39098
rect 6460 39034 6512 39040
rect 6276 39024 6328 39030
rect 6276 38966 6328 38972
rect 6288 38298 6316 38966
rect 6288 38270 6500 38298
rect 6102 38108 6410 38128
rect 6102 38106 6108 38108
rect 6164 38106 6188 38108
rect 6244 38106 6268 38108
rect 6324 38106 6348 38108
rect 6404 38106 6410 38108
rect 6164 38054 6166 38106
rect 6346 38054 6348 38106
rect 6102 38052 6108 38054
rect 6164 38052 6188 38054
rect 6244 38052 6268 38054
rect 6324 38052 6348 38054
rect 6404 38052 6410 38054
rect 6102 38032 6410 38052
rect 6472 37398 6500 38270
rect 6460 37392 6512 37398
rect 6460 37334 6512 37340
rect 6102 37020 6410 37040
rect 6102 37018 6108 37020
rect 6164 37018 6188 37020
rect 6244 37018 6268 37020
rect 6324 37018 6348 37020
rect 6404 37018 6410 37020
rect 6164 36966 6166 37018
rect 6346 36966 6348 37018
rect 6102 36964 6108 36966
rect 6164 36964 6188 36966
rect 6244 36964 6268 36966
rect 6324 36964 6348 36966
rect 6404 36964 6410 36966
rect 6102 36944 6410 36964
rect 6102 35932 6410 35952
rect 6102 35930 6108 35932
rect 6164 35930 6188 35932
rect 6244 35930 6268 35932
rect 6324 35930 6348 35932
rect 6404 35930 6410 35932
rect 6164 35878 6166 35930
rect 6346 35878 6348 35930
rect 6102 35876 6108 35878
rect 6164 35876 6188 35878
rect 6244 35876 6268 35878
rect 6324 35876 6348 35878
rect 6404 35876 6410 35878
rect 6102 35856 6410 35876
rect 6460 35624 6512 35630
rect 6460 35566 6512 35572
rect 6102 34844 6410 34864
rect 6102 34842 6108 34844
rect 6164 34842 6188 34844
rect 6244 34842 6268 34844
rect 6324 34842 6348 34844
rect 6404 34842 6410 34844
rect 6164 34790 6166 34842
rect 6346 34790 6348 34842
rect 6102 34788 6108 34790
rect 6164 34788 6188 34790
rect 6244 34788 6268 34790
rect 6324 34788 6348 34790
rect 6404 34788 6410 34790
rect 6102 34768 6410 34788
rect 6472 34728 6500 35566
rect 6196 34700 6500 34728
rect 6196 34202 6224 34700
rect 6368 34536 6420 34542
rect 6368 34478 6420 34484
rect 6564 34490 6592 42026
rect 6656 41682 6684 42094
rect 6644 41676 6696 41682
rect 6644 41618 6696 41624
rect 6656 41546 6684 41618
rect 6644 41540 6696 41546
rect 6644 41482 6696 41488
rect 6644 40044 6696 40050
rect 6644 39986 6696 39992
rect 6656 39914 6684 39986
rect 6644 39908 6696 39914
rect 6644 39850 6696 39856
rect 6644 38412 6696 38418
rect 6644 38354 6696 38360
rect 6656 37330 6684 38354
rect 6644 37324 6696 37330
rect 6644 37266 6696 37272
rect 6748 35766 6776 43590
rect 7024 42770 7052 43794
rect 7208 43790 7236 44814
rect 7380 44736 7432 44742
rect 7380 44678 7432 44684
rect 7196 43784 7248 43790
rect 7196 43726 7248 43732
rect 7288 43784 7340 43790
rect 7392 43772 7420 44678
rect 7576 43858 7604 44950
rect 7668 44878 7696 45070
rect 7748 44940 7800 44946
rect 7748 44882 7800 44888
rect 7656 44872 7708 44878
rect 7656 44814 7708 44820
rect 7760 44470 7788 44882
rect 7748 44464 7800 44470
rect 7748 44406 7800 44412
rect 8036 44334 8064 45222
rect 8404 44334 8432 45766
rect 8024 44328 8076 44334
rect 8024 44270 8076 44276
rect 8392 44328 8444 44334
rect 8392 44270 8444 44276
rect 7932 44260 7984 44266
rect 7932 44202 7984 44208
rect 7472 43852 7524 43858
rect 7472 43794 7524 43800
rect 7564 43852 7616 43858
rect 7564 43794 7616 43800
rect 7340 43744 7420 43772
rect 7288 43726 7340 43732
rect 7288 43172 7340 43178
rect 7288 43114 7340 43120
rect 7012 42764 7064 42770
rect 7012 42706 7064 42712
rect 7196 42628 7248 42634
rect 7196 42570 7248 42576
rect 7208 41414 7236 42570
rect 7300 42362 7328 43114
rect 7288 42356 7340 42362
rect 7288 42298 7340 42304
rect 7392 42226 7420 43744
rect 7484 43110 7512 43794
rect 7472 43104 7524 43110
rect 7472 43046 7524 43052
rect 7380 42220 7432 42226
rect 7380 42162 7432 42168
rect 7484 42158 7512 43046
rect 7576 42770 7604 43794
rect 7564 42764 7616 42770
rect 7564 42706 7616 42712
rect 7840 42696 7892 42702
rect 7840 42638 7892 42644
rect 7656 42288 7708 42294
rect 7656 42230 7708 42236
rect 7668 42158 7696 42230
rect 7472 42152 7524 42158
rect 7472 42094 7524 42100
rect 7656 42152 7708 42158
rect 7656 42094 7708 42100
rect 7208 41386 7328 41414
rect 6828 40928 6880 40934
rect 6828 40870 6880 40876
rect 7104 40928 7156 40934
rect 7104 40870 7156 40876
rect 6840 39098 6868 40870
rect 7012 39840 7064 39846
rect 7012 39782 7064 39788
rect 7024 39506 7052 39782
rect 7012 39500 7064 39506
rect 7012 39442 7064 39448
rect 6828 39092 6880 39098
rect 6828 39034 6880 39040
rect 7012 38820 7064 38826
rect 6932 38780 7012 38808
rect 6932 38486 6960 38780
rect 7012 38762 7064 38768
rect 6920 38480 6972 38486
rect 6920 38422 6972 38428
rect 6828 37800 6880 37806
rect 6932 37788 6960 38422
rect 6880 37760 6960 37788
rect 6828 37742 6880 37748
rect 6828 37664 6880 37670
rect 6828 37606 6880 37612
rect 6736 35760 6788 35766
rect 6736 35702 6788 35708
rect 6380 34218 6408 34478
rect 6564 34462 6684 34490
rect 6552 34400 6604 34406
rect 6552 34342 6604 34348
rect 6380 34202 6500 34218
rect 6184 34196 6236 34202
rect 6380 34196 6512 34202
rect 6380 34190 6460 34196
rect 6184 34138 6236 34144
rect 6460 34138 6512 34144
rect 6460 34060 6512 34066
rect 6460 34002 6512 34008
rect 6102 33756 6410 33776
rect 6102 33754 6108 33756
rect 6164 33754 6188 33756
rect 6244 33754 6268 33756
rect 6324 33754 6348 33756
rect 6404 33754 6410 33756
rect 6164 33702 6166 33754
rect 6346 33702 6348 33754
rect 6102 33700 6108 33702
rect 6164 33700 6188 33702
rect 6244 33700 6268 33702
rect 6324 33700 6348 33702
rect 6404 33700 6410 33702
rect 6102 33680 6410 33700
rect 6000 33652 6052 33658
rect 6000 33594 6052 33600
rect 5828 33272 5948 33300
rect 5828 32026 5856 33272
rect 6012 33130 6040 33594
rect 6472 33386 6500 34002
rect 6460 33380 6512 33386
rect 6460 33322 6512 33328
rect 5920 33102 6040 33130
rect 5816 32020 5868 32026
rect 5816 31962 5868 31968
rect 5540 31952 5592 31958
rect 5540 31894 5592 31900
rect 5724 31952 5776 31958
rect 5920 31906 5948 33102
rect 6000 32768 6052 32774
rect 6000 32710 6052 32716
rect 6012 32434 6040 32710
rect 6102 32668 6410 32688
rect 6102 32666 6108 32668
rect 6164 32666 6188 32668
rect 6244 32666 6268 32668
rect 6324 32666 6348 32668
rect 6404 32666 6410 32668
rect 6164 32614 6166 32666
rect 6346 32614 6348 32666
rect 6102 32612 6108 32614
rect 6164 32612 6188 32614
rect 6244 32612 6268 32614
rect 6324 32612 6348 32614
rect 6404 32612 6410 32614
rect 6102 32592 6410 32612
rect 6460 32496 6512 32502
rect 6460 32438 6512 32444
rect 6000 32428 6052 32434
rect 6000 32370 6052 32376
rect 6000 32292 6052 32298
rect 6000 32234 6052 32240
rect 5724 31894 5776 31900
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 5448 31680 5500 31686
rect 5448 31622 5500 31628
rect 5460 31346 5488 31622
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 5448 31204 5500 31210
rect 5448 31146 5500 31152
rect 5356 30320 5408 30326
rect 5356 30262 5408 30268
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 5356 30048 5408 30054
rect 5356 29990 5408 29996
rect 5276 29102 5304 29990
rect 5368 29782 5396 29990
rect 5356 29776 5408 29782
rect 5356 29718 5408 29724
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5264 29096 5316 29102
rect 5264 29038 5316 29044
rect 5368 28948 5396 29446
rect 5276 28920 5396 28948
rect 5276 27062 5304 28920
rect 5460 28064 5488 31146
rect 5552 30598 5580 31894
rect 5828 31878 5948 31906
rect 5724 30796 5776 30802
rect 5724 30738 5776 30744
rect 5540 30592 5592 30598
rect 5540 30534 5592 30540
rect 5552 30190 5580 30534
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 5736 30054 5764 30738
rect 5724 30048 5776 30054
rect 5724 29990 5776 29996
rect 5828 29764 5856 31878
rect 5908 31476 5960 31482
rect 5908 31418 5960 31424
rect 5920 30666 5948 31418
rect 5908 30660 5960 30666
rect 5908 30602 5960 30608
rect 5920 29782 5948 30602
rect 5552 29736 5856 29764
rect 5908 29776 5960 29782
rect 5552 28914 5580 29736
rect 5908 29718 5960 29724
rect 6012 29560 6040 32234
rect 6472 31754 6500 32438
rect 6460 31748 6512 31754
rect 6460 31690 6512 31696
rect 6102 31580 6410 31600
rect 6102 31578 6108 31580
rect 6164 31578 6188 31580
rect 6244 31578 6268 31580
rect 6324 31578 6348 31580
rect 6404 31578 6410 31580
rect 6164 31526 6166 31578
rect 6346 31526 6348 31578
rect 6102 31524 6108 31526
rect 6164 31524 6188 31526
rect 6244 31524 6268 31526
rect 6324 31524 6348 31526
rect 6404 31524 6410 31526
rect 6102 31504 6410 31524
rect 6564 31482 6592 34342
rect 6656 32910 6684 34462
rect 6840 34406 6868 37606
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 6932 36378 6960 37266
rect 7012 36576 7064 36582
rect 7012 36518 7064 36524
rect 6920 36372 6972 36378
rect 6920 36314 6972 36320
rect 7024 36258 7052 36518
rect 6932 36242 7052 36258
rect 6920 36236 7052 36242
rect 6972 36230 7052 36236
rect 6920 36178 6972 36184
rect 6932 35562 6960 36178
rect 6920 35556 6972 35562
rect 6920 35498 6972 35504
rect 6736 34400 6788 34406
rect 6736 34342 6788 34348
rect 6828 34400 6880 34406
rect 6828 34342 6880 34348
rect 6748 33046 6776 34342
rect 6828 34196 6880 34202
rect 6828 34138 6880 34144
rect 6736 33040 6788 33046
rect 6736 32982 6788 32988
rect 6840 32978 6868 34138
rect 6932 33998 6960 35498
rect 7012 35148 7064 35154
rect 7012 35090 7064 35096
rect 7024 34542 7052 35090
rect 7012 34536 7064 34542
rect 7012 34478 7064 34484
rect 6920 33992 6972 33998
rect 6920 33934 6972 33940
rect 7024 33504 7052 34478
rect 6932 33476 7052 33504
rect 6828 32972 6880 32978
rect 6932 32960 6960 33476
rect 7116 33402 7144 40870
rect 7196 39432 7248 39438
rect 7196 39374 7248 39380
rect 7208 38554 7236 39374
rect 7196 38548 7248 38554
rect 7196 38490 7248 38496
rect 7300 37806 7328 41386
rect 7852 41002 7880 42638
rect 7944 41414 7972 44202
rect 8024 42764 8076 42770
rect 8024 42706 8076 42712
rect 8036 42158 8064 42706
rect 8024 42152 8076 42158
rect 8024 42094 8076 42100
rect 8116 42084 8168 42090
rect 8116 42026 8168 42032
rect 8128 41682 8156 42026
rect 8116 41676 8168 41682
rect 8116 41618 8168 41624
rect 8300 41608 8352 41614
rect 8300 41550 8352 41556
rect 7944 41386 8064 41414
rect 7840 40996 7892 41002
rect 7840 40938 7892 40944
rect 7840 39976 7892 39982
rect 7840 39918 7892 39924
rect 7472 39500 7524 39506
rect 7472 39442 7524 39448
rect 7380 39092 7432 39098
rect 7380 39034 7432 39040
rect 7288 37800 7340 37806
rect 7288 37742 7340 37748
rect 7392 37738 7420 39034
rect 7484 38010 7512 39442
rect 7852 38894 7880 39918
rect 7840 38888 7892 38894
rect 7840 38830 7892 38836
rect 7852 38554 7880 38830
rect 7840 38548 7892 38554
rect 7840 38490 7892 38496
rect 7656 38208 7708 38214
rect 7656 38150 7708 38156
rect 7472 38004 7524 38010
rect 7472 37946 7524 37952
rect 7564 37800 7616 37806
rect 7564 37742 7616 37748
rect 7380 37732 7432 37738
rect 7380 37674 7432 37680
rect 7196 37664 7248 37670
rect 7196 37606 7248 37612
rect 7208 36922 7236 37606
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 7196 36916 7248 36922
rect 7196 36858 7248 36864
rect 7300 36242 7328 37402
rect 7472 36304 7524 36310
rect 7472 36246 7524 36252
rect 7288 36236 7340 36242
rect 7288 36178 7340 36184
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 7288 36100 7340 36106
rect 7288 36042 7340 36048
rect 7300 35578 7328 36042
rect 7392 35698 7420 36110
rect 7380 35692 7432 35698
rect 7380 35634 7432 35640
rect 7300 35550 7420 35578
rect 7196 35488 7248 35494
rect 7196 35430 7248 35436
rect 7288 35488 7340 35494
rect 7288 35430 7340 35436
rect 6828 32914 6880 32920
rect 6923 32932 6960 32960
rect 7024 33374 7144 33402
rect 6644 32904 6696 32910
rect 6696 32864 6776 32892
rect 6644 32846 6696 32852
rect 6644 32768 6696 32774
rect 6644 32710 6696 32716
rect 6656 31890 6684 32710
rect 6748 32570 6776 32864
rect 6923 32858 6951 32932
rect 7024 32892 7052 33374
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 7116 33046 7144 33254
rect 7104 33040 7156 33046
rect 7104 32982 7156 32988
rect 7024 32864 7144 32892
rect 6828 32836 6880 32842
rect 6923 32830 6960 32858
rect 6828 32778 6880 32784
rect 6736 32564 6788 32570
rect 6736 32506 6788 32512
rect 6840 32366 6868 32778
rect 6828 32360 6880 32366
rect 6828 32302 6880 32308
rect 6932 32298 6960 32830
rect 7116 32484 7144 32864
rect 7024 32456 7144 32484
rect 6920 32292 6972 32298
rect 6920 32234 6972 32240
rect 6920 32020 6972 32026
rect 6920 31962 6972 31968
rect 6736 31952 6788 31958
rect 6736 31894 6788 31900
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6644 31680 6696 31686
rect 6644 31622 6696 31628
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6552 31272 6604 31278
rect 6552 31214 6604 31220
rect 6460 31136 6512 31142
rect 6460 31078 6512 31084
rect 6102 30492 6410 30512
rect 6102 30490 6108 30492
rect 6164 30490 6188 30492
rect 6244 30490 6268 30492
rect 6324 30490 6348 30492
rect 6404 30490 6410 30492
rect 6164 30438 6166 30490
rect 6346 30438 6348 30490
rect 6102 30436 6108 30438
rect 6164 30436 6188 30438
rect 6244 30436 6268 30438
rect 6324 30436 6348 30438
rect 6404 30436 6410 30438
rect 6102 30416 6410 30436
rect 6184 30320 6236 30326
rect 6184 30262 6236 30268
rect 6092 30048 6144 30054
rect 6092 29990 6144 29996
rect 6104 29714 6132 29990
rect 6092 29708 6144 29714
rect 6092 29650 6144 29656
rect 6196 29646 6224 30262
rect 6472 30122 6500 31078
rect 6564 30802 6592 31214
rect 6552 30796 6604 30802
rect 6552 30738 6604 30744
rect 6276 30116 6328 30122
rect 6276 30058 6328 30064
rect 6460 30116 6512 30122
rect 6460 30058 6512 30064
rect 6288 29850 6316 30058
rect 6276 29844 6328 29850
rect 6276 29786 6328 29792
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 5828 29532 6040 29560
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5736 29238 5764 29446
rect 5828 29238 5856 29532
rect 6102 29404 6410 29424
rect 6102 29402 6108 29404
rect 6164 29402 6188 29404
rect 6244 29402 6268 29404
rect 6324 29402 6348 29404
rect 6404 29402 6410 29404
rect 6164 29350 6166 29402
rect 6346 29350 6348 29402
rect 6102 29348 6108 29350
rect 6164 29348 6188 29350
rect 6244 29348 6268 29350
rect 6324 29348 6348 29350
rect 6404 29348 6410 29350
rect 6102 29328 6410 29348
rect 5724 29232 5776 29238
rect 5724 29174 5776 29180
rect 5816 29232 5868 29238
rect 5816 29174 5868 29180
rect 6092 29232 6144 29238
rect 6092 29174 6144 29180
rect 5908 29096 5960 29102
rect 5908 29038 5960 29044
rect 5816 29028 5868 29034
rect 5816 28970 5868 28976
rect 5521 28886 5580 28914
rect 5521 28608 5549 28886
rect 5521 28580 5580 28608
rect 5552 28506 5580 28580
rect 5552 28478 5764 28506
rect 5632 28416 5684 28422
rect 5632 28358 5684 28364
rect 5368 28036 5488 28064
rect 5092 26982 5212 27010
rect 5264 27056 5316 27062
rect 5264 26998 5316 27004
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 5092 25498 5120 26982
rect 5172 26920 5224 26926
rect 5172 26862 5224 26868
rect 5184 26042 5212 26862
rect 5172 26036 5224 26042
rect 5172 25978 5224 25984
rect 5080 25492 5132 25498
rect 5080 25434 5132 25440
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5080 24676 5132 24682
rect 5080 24618 5132 24624
rect 5092 24410 5120 24618
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 5172 23656 5224 23662
rect 5172 23598 5224 23604
rect 5184 23254 5212 23598
rect 5172 23248 5224 23254
rect 5172 23190 5224 23196
rect 5184 22778 5212 23190
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5276 22658 5304 25094
rect 5368 24954 5396 28036
rect 5428 27940 5480 27946
rect 5480 27900 5589 27928
rect 5428 27882 5480 27888
rect 5561 27690 5589 27900
rect 5552 27662 5589 27690
rect 5552 26586 5580 27662
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5540 25696 5592 25702
rect 5540 25638 5592 25644
rect 5356 24948 5408 24954
rect 5356 24890 5408 24896
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 5460 23746 5488 24210
rect 5552 23866 5580 25638
rect 5644 24274 5672 28358
rect 5736 25430 5764 28478
rect 5724 25424 5776 25430
rect 5724 25366 5776 25372
rect 5828 24290 5856 28970
rect 5920 28762 5948 29038
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 5908 28756 5960 28762
rect 5908 28698 5960 28704
rect 6012 27606 6040 28970
rect 6104 28490 6132 29174
rect 6472 28626 6500 30058
rect 6564 29714 6592 30738
rect 6656 30394 6684 31622
rect 6748 31142 6776 31894
rect 6736 31136 6788 31142
rect 6736 31078 6788 31084
rect 6644 30388 6696 30394
rect 6644 30330 6696 30336
rect 6552 29708 6604 29714
rect 6604 29668 6684 29696
rect 6552 29650 6604 29656
rect 6656 29306 6684 29668
rect 6736 29572 6788 29578
rect 6736 29514 6788 29520
rect 6644 29300 6696 29306
rect 6644 29242 6696 29248
rect 6748 29050 6776 29514
rect 6552 29028 6604 29034
rect 6552 28970 6604 28976
rect 6656 29022 6776 29050
rect 6932 29034 6960 31962
rect 7024 31482 7052 32456
rect 7208 32366 7236 35430
rect 7300 33930 7328 35430
rect 7392 34678 7420 35550
rect 7484 35154 7512 36246
rect 7472 35148 7524 35154
rect 7472 35090 7524 35096
rect 7380 34672 7432 34678
rect 7432 34632 7512 34660
rect 7380 34614 7432 34620
rect 7380 34536 7432 34542
rect 7380 34478 7432 34484
rect 7288 33924 7340 33930
rect 7288 33866 7340 33872
rect 7300 33454 7328 33866
rect 7288 33448 7340 33454
rect 7288 33390 7340 33396
rect 7288 33312 7340 33318
rect 7288 33254 7340 33260
rect 7196 32360 7248 32366
rect 7196 32302 7248 32308
rect 7196 32224 7248 32230
rect 7116 32184 7196 32212
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 7024 31210 7052 31418
rect 7012 31204 7064 31210
rect 7012 31146 7064 31152
rect 7116 30190 7144 32184
rect 7196 32166 7248 32172
rect 7300 32042 7328 33254
rect 7392 32502 7420 34478
rect 7380 32496 7432 32502
rect 7380 32438 7432 32444
rect 7380 32292 7432 32298
rect 7380 32234 7432 32240
rect 7208 32014 7328 32042
rect 7012 30184 7064 30190
rect 7012 30126 7064 30132
rect 7104 30184 7156 30190
rect 7104 30126 7156 30132
rect 7024 29510 7052 30126
rect 7012 29504 7064 29510
rect 7012 29446 7064 29452
rect 6920 29028 6972 29034
rect 6460 28620 6512 28626
rect 6460 28562 6512 28568
rect 6092 28484 6144 28490
rect 6092 28426 6144 28432
rect 6102 28316 6410 28336
rect 6102 28314 6108 28316
rect 6164 28314 6188 28316
rect 6244 28314 6268 28316
rect 6324 28314 6348 28316
rect 6404 28314 6410 28316
rect 6164 28262 6166 28314
rect 6346 28262 6348 28314
rect 6102 28260 6108 28262
rect 6164 28260 6188 28262
rect 6244 28260 6268 28262
rect 6324 28260 6348 28262
rect 6404 28260 6410 28262
rect 6102 28240 6410 28260
rect 6184 28144 6236 28150
rect 6184 28086 6236 28092
rect 6196 27614 6224 28086
rect 6472 28082 6500 28562
rect 6460 28076 6512 28082
rect 6460 28018 6512 28024
rect 6460 27940 6512 27946
rect 6460 27882 6512 27888
rect 6000 27600 6052 27606
rect 6196 27586 6316 27614
rect 6000 27542 6052 27548
rect 6288 27470 6316 27586
rect 6472 27470 6500 27882
rect 6276 27464 6328 27470
rect 6276 27406 6328 27412
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6102 27228 6410 27248
rect 6102 27226 6108 27228
rect 6164 27226 6188 27228
rect 6244 27226 6268 27228
rect 6324 27226 6348 27228
rect 6404 27226 6410 27228
rect 6164 27174 6166 27226
rect 6346 27174 6348 27226
rect 6102 27172 6108 27174
rect 6164 27172 6188 27174
rect 6244 27172 6268 27174
rect 6324 27172 6348 27174
rect 6404 27172 6410 27174
rect 6102 27152 6410 27172
rect 5908 26444 5960 26450
rect 5908 26386 5960 26392
rect 5920 26246 5948 26386
rect 6472 26246 6500 27406
rect 5908 26240 5960 26246
rect 5908 26182 5960 26188
rect 6460 26240 6512 26246
rect 6460 26182 6512 26188
rect 6102 26140 6410 26160
rect 6102 26138 6108 26140
rect 6164 26138 6188 26140
rect 6244 26138 6268 26140
rect 6324 26138 6348 26140
rect 6404 26138 6410 26140
rect 6164 26086 6166 26138
rect 6346 26086 6348 26138
rect 6102 26084 6108 26086
rect 6164 26084 6188 26086
rect 6244 26084 6268 26086
rect 6324 26084 6348 26086
rect 6404 26084 6410 26086
rect 6102 26064 6410 26084
rect 6564 25498 6592 28970
rect 6656 27606 6684 29022
rect 6920 28970 6972 28976
rect 6828 28620 6880 28626
rect 6828 28562 6880 28568
rect 6644 27600 6696 27606
rect 6644 27542 6696 27548
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6748 26450 6776 27066
rect 6840 26586 6868 28562
rect 6920 28552 6972 28558
rect 6920 28494 6972 28500
rect 6932 27538 6960 28494
rect 6920 27532 6972 27538
rect 6920 27474 6972 27480
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6828 26444 6880 26450
rect 6828 26386 6880 26392
rect 6840 26042 6868 26386
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 5908 25492 5960 25498
rect 5908 25434 5960 25440
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 5736 24262 5856 24290
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5460 23718 5580 23746
rect 5552 23594 5580 23718
rect 5540 23588 5592 23594
rect 5540 23530 5592 23536
rect 5736 23066 5764 24262
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 5552 23038 5764 23066
rect 5552 22658 5580 23038
rect 5724 22976 5776 22982
rect 5724 22918 5776 22924
rect 5184 22630 5304 22658
rect 5368 22630 5580 22658
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 4896 21412 4948 21418
rect 4896 21354 4948 21360
rect 4724 21304 4844 21332
rect 4620 21286 4672 21292
rect 4528 21004 4580 21010
rect 4528 20946 4580 20952
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 4448 20466 4476 20742
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 4448 18970 4476 19246
rect 4540 19174 4568 20946
rect 4632 19990 4660 21286
rect 4712 20936 4764 20942
rect 4712 20878 4764 20884
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4436 18964 4488 18970
rect 4436 18906 4488 18912
rect 4632 18834 4660 19382
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4356 17190 4476 17218
rect 4264 17088 4384 17116
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16794 4200 16934
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4264 16250 4292 16526
rect 4252 16244 4304 16250
rect 4172 16204 4252 16232
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 14414 4108 15846
rect 4172 14550 4200 16204
rect 4252 16186 4304 16192
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4264 15502 4292 15982
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4356 15366 4384 17088
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4172 13734 4200 14486
rect 4264 14482 4292 14758
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4080 13530 4108 13670
rect 4264 13530 4292 14214
rect 4068 13524 4120 13530
rect 4252 13524 4304 13530
rect 4068 13466 4120 13472
rect 4172 13484 4252 13512
rect 3936 13416 4016 13444
rect 3884 13398 3936 13404
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3896 12986 3924 13262
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 4080 12782 4108 13194
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3896 12322 3924 12650
rect 4172 12374 4200 13484
rect 4252 13466 4304 13472
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4264 12918 4292 13330
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 3804 12294 3924 12322
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 3804 10180 3832 12294
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3896 11286 3924 11562
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3896 10690 3924 10950
rect 3988 10810 4016 12174
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3896 10674 4016 10690
rect 3896 10668 4028 10674
rect 3896 10662 3976 10668
rect 3976 10610 4028 10616
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3896 10248 3924 10542
rect 4080 10248 4108 11290
rect 3896 10220 4108 10248
rect 3804 10152 4016 10180
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9518 3832 9998
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3804 8430 3832 9454
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3804 5166 3832 8366
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3896 4690 3924 9658
rect 3988 7750 4016 10152
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7546 4016 7686
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3988 6934 4016 7210
rect 4080 6934 4108 10220
rect 4172 7256 4200 12038
rect 4264 9518 4292 12718
rect 4356 11286 4384 14350
rect 4448 12102 4476 17190
rect 4540 15314 4568 18158
rect 4724 18086 4752 20878
rect 4816 18766 4844 21304
rect 4896 20868 4948 20874
rect 4896 20810 4948 20816
rect 4908 20398 4936 20810
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4816 17134 4844 18702
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4632 16046 4660 17070
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4724 15706 4752 16594
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4712 15360 4764 15366
rect 4540 15286 4660 15314
rect 4712 15302 4764 15308
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4540 14278 4568 15098
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4540 13190 4568 13942
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4540 12306 4568 13126
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4264 8430 4292 8774
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4252 7268 4304 7274
rect 4172 7228 4252 7256
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4080 6390 4108 6870
rect 4172 6866 4200 7228
rect 4252 7210 4304 7216
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5166 4108 5510
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4172 5098 4200 6802
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 4172 3738 4200 5034
rect 4356 4214 4384 11018
rect 4448 10538 4476 11630
rect 4632 11354 4660 15286
rect 4724 15162 4752 15302
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4724 13954 4752 15098
rect 4816 14958 4844 16594
rect 4908 16250 4936 19926
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 5000 18290 5028 19654
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 5092 16726 5120 21490
rect 5184 20942 5212 22630
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5276 21690 5304 22034
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 5172 20528 5224 20534
rect 5224 20488 5304 20516
rect 5172 20470 5224 20476
rect 5276 20482 5304 20488
rect 5368 20482 5396 22630
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5460 22094 5488 22510
rect 5460 22066 5580 22094
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5276 20454 5396 20482
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5184 19854 5212 20266
rect 5276 19938 5304 20454
rect 5460 20398 5488 21422
rect 5448 20392 5500 20398
rect 5368 20352 5448 20380
rect 5368 20058 5396 20352
rect 5448 20334 5500 20340
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5276 19910 5396 19938
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5184 19446 5212 19790
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5172 19440 5224 19446
rect 5172 19382 5224 19388
rect 5276 18834 5304 19722
rect 5368 19334 5396 19910
rect 5460 19446 5488 20198
rect 5448 19440 5500 19446
rect 5448 19382 5500 19388
rect 5368 19306 5488 19334
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5184 17678 5212 18566
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 17270 5304 17478
rect 5264 17264 5316 17270
rect 5264 17206 5316 17212
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4908 14074 4936 16050
rect 4988 15972 5040 15978
rect 5092 15960 5120 16662
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5040 15932 5120 15960
rect 4988 15914 5040 15920
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5000 14482 5028 15438
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5092 14550 5120 14894
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4724 13926 4936 13954
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 11354 4752 13262
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4816 11234 4844 13738
rect 4540 11206 4844 11234
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4448 9518 4476 10474
rect 4540 9654 4568 11206
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4632 9722 4660 10542
rect 4724 10130 4752 11086
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4540 8906 4568 9590
rect 4632 9518 4660 9658
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4620 9036 4672 9042
rect 4724 9024 4752 9862
rect 4816 9178 4844 11086
rect 4908 11082 4936 13926
rect 5000 12986 5028 14418
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 5092 13802 5120 14350
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 5000 10724 5028 12786
rect 5092 12782 5120 13330
rect 5184 13326 5212 16186
rect 5276 16046 5304 16934
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5276 15570 5304 15982
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5276 14890 5304 15506
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 13802 5304 14418
rect 5368 14414 5396 17070
rect 5460 16114 5488 19306
rect 5552 18358 5580 22066
rect 5644 21554 5672 22646
rect 5736 22098 5764 22918
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5828 21978 5856 24074
rect 5920 23662 5948 25434
rect 6102 25052 6410 25072
rect 6102 25050 6108 25052
rect 6164 25050 6188 25052
rect 6244 25050 6268 25052
rect 6324 25050 6348 25052
rect 6404 25050 6410 25052
rect 6164 24998 6166 25050
rect 6346 24998 6348 25050
rect 6102 24996 6108 24998
rect 6164 24996 6188 24998
rect 6244 24996 6268 24998
rect 6324 24996 6348 24998
rect 6404 24996 6410 24998
rect 6102 24976 6410 24996
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 6012 23730 6040 24210
rect 6380 24138 6408 24550
rect 6564 24206 6592 24754
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6368 24132 6420 24138
rect 6368 24074 6420 24080
rect 6102 23964 6410 23984
rect 6102 23962 6108 23964
rect 6164 23962 6188 23964
rect 6244 23962 6268 23964
rect 6324 23962 6348 23964
rect 6404 23962 6410 23964
rect 6164 23910 6166 23962
rect 6346 23910 6348 23962
rect 6102 23908 6108 23910
rect 6164 23908 6188 23910
rect 6244 23908 6268 23910
rect 6324 23908 6348 23910
rect 6404 23908 6410 23910
rect 6102 23888 6410 23908
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 5908 23656 5960 23662
rect 5908 23598 5960 23604
rect 5920 23050 5948 23598
rect 6012 23186 6040 23666
rect 6000 23180 6052 23186
rect 6000 23122 6052 23128
rect 5908 23044 5960 23050
rect 5908 22986 5960 22992
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 5920 22166 5948 22714
rect 6012 22574 6040 23122
rect 6564 23050 6592 24142
rect 6552 23044 6604 23050
rect 6552 22986 6604 22992
rect 6102 22876 6410 22896
rect 6102 22874 6108 22876
rect 6164 22874 6188 22876
rect 6244 22874 6268 22876
rect 6324 22874 6348 22876
rect 6404 22874 6410 22876
rect 6164 22822 6166 22874
rect 6346 22822 6348 22874
rect 6102 22820 6108 22822
rect 6164 22820 6188 22822
rect 6244 22820 6268 22822
rect 6324 22820 6348 22822
rect 6404 22820 6410 22822
rect 6102 22800 6410 22820
rect 6564 22642 6592 22986
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6552 22636 6604 22642
rect 6552 22578 6604 22584
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 5908 22160 5960 22166
rect 5908 22102 5960 22108
rect 5736 21950 5856 21978
rect 6288 21962 6316 22578
rect 6460 22568 6512 22574
rect 6460 22510 6512 22516
rect 5908 21956 5960 21962
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5736 21434 5764 21950
rect 5908 21898 5960 21904
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5828 21622 5856 21830
rect 5816 21616 5868 21622
rect 5816 21558 5868 21564
rect 5816 21480 5868 21486
rect 5736 21428 5816 21434
rect 5736 21422 5868 21428
rect 5736 21406 5856 21422
rect 5828 20466 5856 21406
rect 5920 21078 5948 21898
rect 6102 21788 6410 21808
rect 6102 21786 6108 21788
rect 6164 21786 6188 21788
rect 6244 21786 6268 21788
rect 6324 21786 6348 21788
rect 6404 21786 6410 21788
rect 6164 21734 6166 21786
rect 6346 21734 6348 21786
rect 6102 21732 6108 21734
rect 6164 21732 6188 21734
rect 6244 21732 6268 21734
rect 6324 21732 6348 21734
rect 6404 21732 6410 21734
rect 6102 21712 6410 21732
rect 6472 21486 6500 22510
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 21554 6592 21966
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 6012 21010 6040 21422
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5644 18426 5672 19246
rect 5828 18834 5856 20402
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 17746 5672 18226
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5552 17202 5580 17614
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5736 17134 5764 18022
rect 5920 17626 5948 20878
rect 6102 20700 6410 20720
rect 6102 20698 6108 20700
rect 6164 20698 6188 20700
rect 6244 20698 6268 20700
rect 6324 20698 6348 20700
rect 6404 20698 6410 20700
rect 6164 20646 6166 20698
rect 6346 20646 6348 20698
rect 6102 20644 6108 20646
rect 6164 20644 6188 20646
rect 6244 20644 6268 20646
rect 6324 20644 6348 20646
rect 6404 20644 6410 20646
rect 6102 20624 6410 20644
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6012 19786 6040 20198
rect 6564 19922 6592 20334
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6012 19310 6040 19722
rect 6102 19612 6410 19632
rect 6102 19610 6108 19612
rect 6164 19610 6188 19612
rect 6244 19610 6268 19612
rect 6324 19610 6348 19612
rect 6404 19610 6410 19612
rect 6164 19558 6166 19610
rect 6346 19558 6348 19610
rect 6102 19556 6108 19558
rect 6164 19556 6188 19558
rect 6244 19556 6268 19558
rect 6324 19556 6348 19558
rect 6404 19556 6410 19558
rect 6102 19536 6410 19556
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6102 18524 6410 18544
rect 6102 18522 6108 18524
rect 6164 18522 6188 18524
rect 6244 18522 6268 18524
rect 6324 18522 6348 18524
rect 6404 18522 6410 18524
rect 6164 18470 6166 18522
rect 6346 18470 6348 18522
rect 6102 18468 6108 18470
rect 6164 18468 6188 18470
rect 6244 18468 6268 18470
rect 6324 18468 6348 18470
rect 6404 18468 6410 18470
rect 6102 18448 6410 18468
rect 6472 18222 6500 18566
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5828 17598 5948 17626
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5460 14260 5488 16050
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15026 5580 15846
rect 5632 15496 5684 15502
rect 5828 15450 5856 17598
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5632 15438 5684 15444
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5644 14618 5672 15438
rect 5736 15422 5856 15450
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5368 14232 5488 14260
rect 5540 14272 5592 14278
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 12306 5120 12582
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4908 10696 5028 10724
rect 4908 9674 4936 10696
rect 5092 10470 5120 11290
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4908 9654 5028 9674
rect 4908 9648 5040 9654
rect 4908 9646 4988 9648
rect 4988 9590 5040 9596
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4908 9042 4936 9386
rect 4672 8996 4752 9024
rect 4620 8978 4672 8984
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4448 6254 4476 6666
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4448 4690 4476 6190
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5778 4568 6054
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4632 5710 4660 8978
rect 4724 8838 4752 8996
rect 4896 9036 4948 9042
rect 5080 9036 5132 9042
rect 4948 8996 5080 9024
rect 4896 8978 4948 8984
rect 5080 8978 5132 8984
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 5092 8566 5120 8978
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 7546 4752 7822
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4816 6458 4844 7890
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4816 5846 4844 6394
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 4826 4660 5646
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4436 4684 4488 4690
rect 4632 4672 4660 4762
rect 4712 4684 4764 4690
rect 4632 4644 4712 4672
rect 4436 4626 4488 4632
rect 4712 4626 4764 4632
rect 4448 4282 4476 4626
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4908 4010 4936 7142
rect 5000 5778 5028 7822
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5092 6458 5120 7278
rect 5184 7206 5212 13126
rect 5276 12374 5304 13466
rect 5368 13190 5396 14232
rect 5540 14214 5592 14220
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13258 5488 13806
rect 5552 13410 5580 14214
rect 5644 13938 5672 14214
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5736 13530 5764 15422
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5828 14958 5856 15302
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5828 13530 5856 14282
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5552 13382 5856 13410
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5276 6866 5304 12174
rect 5368 11354 5396 12242
rect 5460 11830 5488 13194
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12986 5764 13126
rect 5828 13002 5856 13382
rect 5920 13190 5948 17478
rect 6012 17270 6040 18022
rect 6460 17604 6512 17610
rect 6460 17546 6512 17552
rect 6102 17436 6410 17456
rect 6102 17434 6108 17436
rect 6164 17434 6188 17436
rect 6244 17434 6268 17436
rect 6324 17434 6348 17436
rect 6404 17434 6410 17436
rect 6164 17382 6166 17434
rect 6346 17382 6348 17434
rect 6102 17380 6108 17382
rect 6164 17380 6188 17382
rect 6244 17380 6268 17382
rect 6324 17380 6348 17382
rect 6404 17380 6410 17382
rect 6102 17360 6410 17380
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 6472 17066 6500 17546
rect 6564 17134 6592 19110
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6012 15094 6040 17002
rect 6656 16640 6684 25842
rect 6932 25770 6960 27474
rect 7024 26994 7052 29446
rect 7208 29238 7236 32014
rect 7288 30932 7340 30938
rect 7288 30874 7340 30880
rect 7300 30326 7328 30874
rect 7392 30870 7420 32234
rect 7380 30864 7432 30870
rect 7380 30806 7432 30812
rect 7288 30320 7340 30326
rect 7288 30262 7340 30268
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7196 29028 7248 29034
rect 7116 28976 7196 28994
rect 7116 28970 7248 28976
rect 7116 28966 7236 28970
rect 7116 28218 7144 28966
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7104 28212 7156 28218
rect 7104 28154 7156 28160
rect 7208 28082 7236 28494
rect 7300 28490 7328 30262
rect 7288 28484 7340 28490
rect 7288 28426 7340 28432
rect 7196 28076 7248 28082
rect 7196 28018 7248 28024
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 7116 27674 7144 27950
rect 7104 27668 7156 27674
rect 7104 27610 7156 27616
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 7012 26240 7064 26246
rect 7012 26182 7064 26188
rect 7024 25838 7052 26182
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 6920 25764 6972 25770
rect 6920 25706 6972 25712
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6840 25362 6868 25638
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 6736 23792 6788 23798
rect 6736 23734 6788 23740
rect 6748 23662 6776 23734
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 6748 23186 6776 23598
rect 6840 23322 6868 25298
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 7024 23254 7052 24006
rect 7012 23248 7064 23254
rect 7012 23190 7064 23196
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 6748 22710 6776 23122
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6736 22704 6788 22710
rect 6736 22646 6788 22652
rect 6840 22098 6868 22918
rect 6932 22574 6960 23122
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 7116 22438 7144 27610
rect 7208 27402 7236 28018
rect 7300 28014 7328 28426
rect 7288 28008 7340 28014
rect 7288 27950 7340 27956
rect 7196 27396 7248 27402
rect 7196 27338 7248 27344
rect 7208 26518 7236 27338
rect 7196 26512 7248 26518
rect 7196 26454 7248 26460
rect 7208 25838 7236 26454
rect 7196 25832 7248 25838
rect 7196 25774 7248 25780
rect 7288 25764 7340 25770
rect 7288 25706 7340 25712
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6748 19310 6776 21082
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 7024 20398 7052 21014
rect 7012 20392 7064 20398
rect 6932 20352 7012 20380
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6748 18290 6776 19246
rect 6840 19242 6868 19654
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6840 18970 6868 19178
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6932 18766 6960 20352
rect 7012 20334 7064 20340
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 7024 19514 7052 19654
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 7024 18222 7052 18770
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6932 17610 6960 17682
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6472 16612 6684 16640
rect 6102 16348 6410 16368
rect 6102 16346 6108 16348
rect 6164 16346 6188 16348
rect 6244 16346 6268 16348
rect 6324 16346 6348 16348
rect 6404 16346 6410 16348
rect 6164 16294 6166 16346
rect 6346 16294 6348 16346
rect 6102 16292 6108 16294
rect 6164 16292 6188 16294
rect 6244 16292 6268 16294
rect 6324 16292 6348 16294
rect 6404 16292 6410 16294
rect 6102 16272 6410 16292
rect 6472 16046 6500 16612
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 16114 6592 16458
rect 6552 16108 6604 16114
rect 6604 16068 6684 16096
rect 6552 16050 6604 16056
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6102 15260 6410 15280
rect 6102 15258 6108 15260
rect 6164 15258 6188 15260
rect 6244 15258 6268 15260
rect 6324 15258 6348 15260
rect 6404 15258 6410 15260
rect 6164 15206 6166 15258
rect 6346 15206 6348 15258
rect 6102 15204 6108 15206
rect 6164 15204 6188 15206
rect 6244 15204 6268 15206
rect 6324 15204 6348 15206
rect 6404 15204 6410 15206
rect 6102 15184 6410 15204
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 6012 14550 6040 15030
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6472 14414 6500 15982
rect 6656 14482 6684 16068
rect 6748 16046 6776 16730
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7024 16250 7052 16594
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6460 14408 6512 14414
rect 6512 14368 6592 14396
rect 6460 14350 6512 14356
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6102 14172 6410 14192
rect 6102 14170 6108 14172
rect 6164 14170 6188 14172
rect 6244 14170 6268 14172
rect 6324 14170 6348 14172
rect 6404 14170 6410 14172
rect 6164 14118 6166 14170
rect 6346 14118 6348 14170
rect 6102 14116 6108 14118
rect 6164 14116 6188 14118
rect 6244 14116 6268 14118
rect 6324 14116 6348 14118
rect 6404 14116 6410 14118
rect 6102 14096 6410 14116
rect 6472 13870 6500 14214
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5724 12980 5776 12986
rect 5828 12974 5948 13002
rect 5724 12922 5776 12928
rect 5736 12832 5764 12922
rect 5736 12804 5856 12832
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5552 11830 5580 12650
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5460 11626 5488 11766
rect 5644 11676 5672 12242
rect 5552 11648 5672 11676
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5368 10266 5396 11154
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5460 10130 5488 11562
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5368 9178 5396 10066
rect 5552 9874 5580 11648
rect 5736 10606 5764 12650
rect 5828 12238 5856 12804
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 10810 5856 11290
rect 5920 11098 5948 12974
rect 6012 11354 6040 13670
rect 6564 13258 6592 14368
rect 6656 13870 6684 14418
rect 6748 14346 6776 15030
rect 6840 14498 6868 15914
rect 6840 14482 7052 14498
rect 6840 14476 7064 14482
rect 6840 14470 7012 14476
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6102 13084 6410 13104
rect 6102 13082 6108 13084
rect 6164 13082 6188 13084
rect 6244 13082 6268 13084
rect 6324 13082 6348 13084
rect 6404 13082 6410 13084
rect 6164 13030 6166 13082
rect 6346 13030 6348 13082
rect 6102 13028 6108 13030
rect 6164 13028 6188 13030
rect 6244 13028 6268 13030
rect 6324 13028 6348 13030
rect 6404 13028 6410 13030
rect 6102 13008 6410 13028
rect 6564 12850 6592 13194
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6656 12782 6684 13398
rect 6748 13394 6776 14010
rect 6840 13462 6868 14470
rect 7012 14418 7064 14424
rect 7116 14346 7144 22374
rect 7208 21434 7236 23530
rect 7300 23338 7328 25706
rect 7392 23526 7420 30806
rect 7484 30326 7512 34632
rect 7576 33522 7604 37742
rect 7668 36922 7696 38150
rect 8036 37274 8064 41386
rect 8312 41138 8340 41550
rect 8496 41414 8524 48146
rect 14924 48068 14976 48074
rect 14924 48010 14976 48016
rect 11612 48000 11664 48006
rect 11612 47942 11664 47948
rect 11624 47734 11652 47942
rect 14936 47734 14964 48010
rect 11612 47728 11664 47734
rect 11612 47670 11664 47676
rect 14924 47728 14976 47734
rect 14924 47670 14976 47676
rect 10416 47592 10468 47598
rect 10416 47534 10468 47540
rect 10428 47190 10456 47534
rect 10968 47524 11020 47530
rect 10968 47466 11020 47472
rect 10876 47456 10928 47462
rect 10796 47416 10876 47444
rect 10416 47184 10468 47190
rect 10416 47126 10468 47132
rect 9864 47116 9916 47122
rect 9864 47058 9916 47064
rect 9220 46912 9272 46918
rect 9220 46854 9272 46860
rect 9232 46578 9260 46854
rect 9220 46572 9272 46578
rect 9220 46514 9272 46520
rect 9496 46572 9548 46578
rect 9496 46514 9548 46520
rect 9036 46504 9088 46510
rect 9036 46446 9088 46452
rect 9048 46034 9076 46446
rect 9232 46034 9260 46514
rect 9404 46504 9456 46510
rect 9404 46446 9456 46452
rect 9416 46170 9444 46446
rect 9404 46164 9456 46170
rect 9404 46106 9456 46112
rect 9508 46034 9536 46514
rect 9680 46504 9732 46510
rect 9680 46446 9732 46452
rect 9692 46102 9720 46446
rect 9772 46436 9824 46442
rect 9772 46378 9824 46384
rect 9680 46096 9732 46102
rect 9680 46038 9732 46044
rect 9784 46034 9812 46378
rect 9876 46170 9904 47058
rect 10428 46510 10456 47126
rect 10416 46504 10468 46510
rect 10416 46446 10468 46452
rect 9864 46164 9916 46170
rect 9864 46106 9916 46112
rect 10796 46034 10824 47416
rect 10876 47398 10928 47404
rect 10876 46912 10928 46918
rect 10876 46854 10928 46860
rect 9036 46028 9088 46034
rect 9036 45970 9088 45976
rect 9220 46028 9272 46034
rect 9220 45970 9272 45976
rect 9496 46028 9548 46034
rect 9496 45970 9548 45976
rect 9772 46028 9824 46034
rect 9772 45970 9824 45976
rect 10232 46028 10284 46034
rect 10784 46028 10836 46034
rect 10232 45970 10284 45976
rect 10704 45988 10784 46016
rect 9232 45422 9260 45970
rect 9508 45626 9536 45970
rect 9784 45898 9812 45970
rect 9772 45892 9824 45898
rect 9772 45834 9824 45840
rect 10244 45830 10272 45970
rect 10508 45960 10560 45966
rect 10508 45902 10560 45908
rect 10600 45960 10652 45966
rect 10600 45902 10652 45908
rect 10232 45824 10284 45830
rect 10232 45766 10284 45772
rect 9496 45620 9548 45626
rect 9496 45562 9548 45568
rect 9864 45552 9916 45558
rect 9864 45494 9916 45500
rect 9220 45416 9272 45422
rect 9220 45358 9272 45364
rect 9496 45348 9548 45354
rect 9496 45290 9548 45296
rect 9312 44872 9364 44878
rect 9312 44814 9364 44820
rect 9128 44192 9180 44198
rect 9128 44134 9180 44140
rect 9220 44192 9272 44198
rect 9220 44134 9272 44140
rect 8576 43784 8628 43790
rect 8576 43726 8628 43732
rect 8588 42294 8616 43726
rect 9140 42770 9168 44134
rect 9232 43246 9260 44134
rect 9324 43790 9352 44814
rect 9508 44470 9536 45290
rect 9772 45280 9824 45286
rect 9772 45222 9824 45228
rect 9496 44464 9548 44470
rect 9496 44406 9548 44412
rect 9508 43858 9536 44406
rect 9496 43852 9548 43858
rect 9496 43794 9548 43800
rect 9312 43784 9364 43790
rect 9312 43726 9364 43732
rect 9324 43450 9352 43726
rect 9312 43444 9364 43450
rect 9312 43386 9364 43392
rect 9220 43240 9272 43246
rect 9220 43182 9272 43188
rect 9232 42906 9260 43182
rect 9496 43104 9548 43110
rect 9496 43046 9548 43052
rect 9220 42900 9272 42906
rect 9220 42842 9272 42848
rect 9404 42900 9456 42906
rect 9404 42842 9456 42848
rect 9128 42764 9180 42770
rect 9128 42706 9180 42712
rect 9128 42560 9180 42566
rect 9128 42502 9180 42508
rect 8576 42288 8628 42294
rect 8576 42230 8628 42236
rect 8588 41682 8616 42230
rect 9140 42158 9168 42502
rect 9416 42294 9444 42842
rect 9404 42288 9456 42294
rect 9404 42230 9456 42236
rect 8944 42152 8996 42158
rect 8944 42094 8996 42100
rect 9128 42152 9180 42158
rect 9128 42094 9180 42100
rect 8956 41818 8984 42094
rect 9416 42090 9444 42230
rect 9508 42158 9536 43046
rect 9784 42770 9812 45222
rect 9876 44266 9904 45494
rect 10244 44946 10272 45766
rect 10232 44940 10284 44946
rect 10232 44882 10284 44888
rect 9956 44872 10008 44878
rect 9956 44814 10008 44820
rect 9864 44260 9916 44266
rect 9864 44202 9916 44208
rect 9876 43314 9904 44202
rect 9968 43790 9996 44814
rect 10140 44736 10192 44742
rect 10140 44678 10192 44684
rect 9956 43784 10008 43790
rect 9956 43726 10008 43732
rect 9968 43314 9996 43726
rect 9864 43308 9916 43314
rect 9864 43250 9916 43256
rect 9956 43308 10008 43314
rect 9956 43250 10008 43256
rect 9956 42900 10008 42906
rect 9956 42842 10008 42848
rect 9772 42764 9824 42770
rect 9772 42706 9824 42712
rect 9588 42696 9640 42702
rect 9588 42638 9640 42644
rect 9496 42152 9548 42158
rect 9496 42094 9548 42100
rect 9600 42090 9628 42638
rect 9968 42362 9996 42842
rect 10152 42650 10180 44678
rect 10244 43246 10272 44882
rect 10520 44878 10548 45902
rect 10612 45626 10640 45902
rect 10600 45620 10652 45626
rect 10600 45562 10652 45568
rect 10612 44878 10640 45562
rect 10704 45082 10732 45988
rect 10784 45970 10836 45976
rect 10888 45898 10916 46854
rect 10980 46170 11008 47466
rect 11253 47356 11561 47376
rect 11253 47354 11259 47356
rect 11315 47354 11339 47356
rect 11395 47354 11419 47356
rect 11475 47354 11499 47356
rect 11555 47354 11561 47356
rect 11315 47302 11317 47354
rect 11497 47302 11499 47354
rect 11253 47300 11259 47302
rect 11315 47300 11339 47302
rect 11395 47300 11419 47302
rect 11475 47300 11499 47302
rect 11555 47300 11561 47302
rect 11253 47280 11561 47300
rect 11624 46986 11652 47670
rect 12900 47660 12952 47666
rect 12900 47602 12952 47608
rect 12808 47456 12860 47462
rect 12808 47398 12860 47404
rect 12820 47190 12848 47398
rect 12808 47184 12860 47190
rect 12808 47126 12860 47132
rect 12164 47048 12216 47054
rect 12164 46990 12216 46996
rect 11612 46980 11664 46986
rect 11612 46922 11664 46928
rect 11253 46268 11561 46288
rect 11253 46266 11259 46268
rect 11315 46266 11339 46268
rect 11395 46266 11419 46268
rect 11475 46266 11499 46268
rect 11555 46266 11561 46268
rect 11315 46214 11317 46266
rect 11497 46214 11499 46266
rect 11253 46212 11259 46214
rect 11315 46212 11339 46214
rect 11395 46212 11419 46214
rect 11475 46212 11499 46214
rect 11555 46212 11561 46214
rect 11253 46192 11561 46212
rect 10968 46164 11020 46170
rect 10968 46106 11020 46112
rect 10876 45892 10928 45898
rect 10876 45834 10928 45840
rect 10888 45422 10916 45834
rect 10968 45824 11020 45830
rect 10968 45766 11020 45772
rect 10876 45416 10928 45422
rect 10876 45358 10928 45364
rect 10784 45280 10836 45286
rect 10784 45222 10836 45228
rect 10692 45076 10744 45082
rect 10692 45018 10744 45024
rect 10704 44946 10732 45018
rect 10692 44940 10744 44946
rect 10692 44882 10744 44888
rect 10508 44872 10560 44878
rect 10508 44814 10560 44820
rect 10600 44872 10652 44878
rect 10600 44814 10652 44820
rect 10600 44396 10652 44402
rect 10600 44338 10652 44344
rect 10508 44328 10560 44334
rect 10508 44270 10560 44276
rect 10324 43376 10376 43382
rect 10324 43318 10376 43324
rect 10232 43240 10284 43246
rect 10232 43182 10284 43188
rect 10152 42622 10272 42650
rect 10048 42560 10100 42566
rect 10048 42502 10100 42508
rect 10140 42560 10192 42566
rect 10140 42502 10192 42508
rect 9956 42356 10008 42362
rect 9956 42298 10008 42304
rect 9404 42084 9456 42090
rect 9404 42026 9456 42032
rect 9588 42084 9640 42090
rect 9588 42026 9640 42032
rect 8760 41812 8812 41818
rect 8760 41754 8812 41760
rect 8944 41812 8996 41818
rect 8944 41754 8996 41760
rect 8576 41676 8628 41682
rect 8576 41618 8628 41624
rect 8668 41608 8720 41614
rect 8668 41550 8720 41556
rect 8404 41386 8524 41414
rect 8300 41132 8352 41138
rect 8300 41074 8352 41080
rect 8312 40662 8340 41074
rect 8300 40656 8352 40662
rect 8300 40598 8352 40604
rect 8312 39506 8340 40598
rect 8404 39658 8432 41386
rect 8484 41064 8536 41070
rect 8484 41006 8536 41012
rect 8496 40730 8524 41006
rect 8576 40996 8628 41002
rect 8576 40938 8628 40944
rect 8484 40724 8536 40730
rect 8484 40666 8536 40672
rect 8496 40594 8524 40666
rect 8484 40588 8536 40594
rect 8484 40530 8536 40536
rect 8404 39630 8524 39658
rect 8300 39500 8352 39506
rect 8300 39442 8352 39448
rect 8392 39500 8444 39506
rect 8392 39442 8444 39448
rect 8208 39364 8260 39370
rect 8208 39306 8260 39312
rect 8116 38888 8168 38894
rect 8116 38830 8168 38836
rect 8128 38350 8156 38830
rect 8116 38344 8168 38350
rect 8116 38286 8168 38292
rect 8036 37246 8156 37274
rect 7656 36916 7708 36922
rect 7656 36858 7708 36864
rect 7748 36848 7800 36854
rect 7748 36790 7800 36796
rect 7656 36236 7708 36242
rect 7656 36178 7708 36184
rect 7668 34678 7696 36178
rect 7656 34672 7708 34678
rect 7656 34614 7708 34620
rect 7656 34468 7708 34474
rect 7656 34410 7708 34416
rect 7564 33516 7616 33522
rect 7564 33458 7616 33464
rect 7564 33312 7616 33318
rect 7564 33254 7616 33260
rect 7576 31822 7604 33254
rect 7668 32570 7696 34410
rect 7656 32564 7708 32570
rect 7656 32506 7708 32512
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7656 31816 7708 31822
rect 7656 31758 7708 31764
rect 7668 31482 7696 31758
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7760 30938 7788 36790
rect 8128 35894 8156 37246
rect 8220 36650 8248 39306
rect 8404 39098 8432 39442
rect 8392 39092 8444 39098
rect 8392 39034 8444 39040
rect 8496 37482 8524 39630
rect 8404 37466 8524 37482
rect 8392 37460 8524 37466
rect 8444 37454 8524 37460
rect 8392 37402 8444 37408
rect 8208 36644 8260 36650
rect 8208 36586 8260 36592
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 8404 36378 8432 36518
rect 8392 36372 8444 36378
rect 8392 36314 8444 36320
rect 8128 35866 8248 35894
rect 7932 35624 7984 35630
rect 7932 35566 7984 35572
rect 7840 35148 7892 35154
rect 7840 35090 7892 35096
rect 7852 34746 7880 35090
rect 7840 34740 7892 34746
rect 7840 34682 7892 34688
rect 7944 34610 7972 35566
rect 7932 34604 7984 34610
rect 7932 34546 7984 34552
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 7852 31958 7880 33390
rect 7840 31952 7892 31958
rect 7840 31894 7892 31900
rect 7840 31340 7892 31346
rect 7840 31282 7892 31288
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7852 30394 7880 31282
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 7472 30320 7524 30326
rect 7472 30262 7524 30268
rect 7484 29646 7512 30262
rect 7944 30258 7972 34546
rect 8116 34536 8168 34542
rect 8116 34478 8168 34484
rect 8024 33312 8076 33318
rect 8024 33254 8076 33260
rect 8036 32366 8064 33254
rect 8128 32774 8156 34478
rect 8116 32768 8168 32774
rect 8116 32710 8168 32716
rect 8116 32496 8168 32502
rect 8116 32438 8168 32444
rect 8024 32360 8076 32366
rect 8024 32302 8076 32308
rect 8024 32224 8076 32230
rect 8024 32166 8076 32172
rect 8036 31482 8064 32166
rect 8128 31872 8156 32438
rect 8220 32230 8248 35866
rect 8484 35216 8536 35222
rect 8484 35158 8536 35164
rect 8300 34060 8352 34066
rect 8300 34002 8352 34008
rect 8312 33046 8340 34002
rect 8300 33040 8352 33046
rect 8300 32982 8352 32988
rect 8312 32774 8340 32982
rect 8300 32768 8352 32774
rect 8300 32710 8352 32716
rect 8208 32224 8260 32230
rect 8208 32166 8260 32172
rect 8300 32224 8352 32230
rect 8300 32166 8352 32172
rect 8208 31884 8260 31890
rect 8128 31844 8208 31872
rect 8208 31826 8260 31832
rect 8116 31680 8168 31686
rect 8116 31622 8168 31628
rect 8024 31476 8076 31482
rect 8024 31418 8076 31424
rect 8024 30796 8076 30802
rect 8024 30738 8076 30744
rect 8036 30394 8064 30738
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 8128 30274 8156 31622
rect 8220 30938 8248 31826
rect 8312 31822 8340 32166
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 8496 31686 8524 35158
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8484 31204 8536 31210
rect 8484 31146 8536 31152
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 8036 30246 8156 30274
rect 7564 30048 7616 30054
rect 7564 29990 7616 29996
rect 7576 29714 7604 29990
rect 7840 29776 7892 29782
rect 7840 29718 7892 29724
rect 7564 29708 7616 29714
rect 7564 29650 7616 29656
rect 7656 29708 7708 29714
rect 7656 29650 7708 29656
rect 7472 29640 7524 29646
rect 7472 29582 7524 29588
rect 7484 24818 7512 29582
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7576 27470 7604 28018
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7564 27056 7616 27062
rect 7564 26998 7616 27004
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7484 23730 7512 24754
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7380 23520 7432 23526
rect 7380 23462 7432 23468
rect 7300 23310 7420 23338
rect 7208 21406 7328 21434
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7208 17610 7236 21286
rect 7300 21146 7328 21406
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7208 14890 7236 16050
rect 7300 15978 7328 19450
rect 7392 19334 7420 23310
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7484 23186 7512 23258
rect 7472 23180 7524 23186
rect 7472 23122 7524 23128
rect 7484 22234 7512 23122
rect 7576 22642 7604 26998
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7668 22574 7696 29650
rect 7852 28966 7880 29718
rect 7944 29646 7972 30194
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7944 28626 7972 29582
rect 8036 29510 8064 30246
rect 8220 30190 8248 30874
rect 8208 30184 8260 30190
rect 8208 30126 8260 30132
rect 8312 30054 8340 31078
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8116 30048 8168 30054
rect 8116 29990 8168 29996
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8024 29504 8076 29510
rect 8024 29446 8076 29452
rect 7932 28620 7984 28626
rect 7932 28562 7984 28568
rect 7840 28484 7892 28490
rect 7840 28426 7892 28432
rect 7852 28014 7880 28426
rect 7840 28008 7892 28014
rect 7760 27968 7840 27996
rect 7760 27606 7788 27968
rect 7840 27950 7892 27956
rect 7748 27600 7800 27606
rect 7748 27542 7800 27548
rect 7760 26450 7788 27542
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 7852 26586 7880 27474
rect 8036 26602 8064 29446
rect 7840 26580 7892 26586
rect 7840 26522 7892 26528
rect 7944 26574 8064 26602
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 7760 25922 7788 26386
rect 7760 25906 7880 25922
rect 7748 25900 7880 25906
rect 7800 25894 7880 25900
rect 7748 25842 7800 25848
rect 7748 25764 7800 25770
rect 7748 25706 7800 25712
rect 7760 25158 7788 25706
rect 7852 25362 7880 25894
rect 7840 25356 7892 25362
rect 7840 25298 7892 25304
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 7944 24410 7972 26574
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 8036 24750 8064 25774
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 7852 23866 7880 24210
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7852 23254 7880 23598
rect 8036 23322 8064 24686
rect 8128 24410 8156 29990
rect 8312 28150 8340 29990
rect 8404 29170 8432 30534
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 8300 28144 8352 28150
rect 8300 28086 8352 28092
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8220 27878 8248 28018
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 8220 26926 8248 27814
rect 8404 27538 8432 29106
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8404 27130 8432 27474
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 8220 26382 8248 26862
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8220 26042 8248 26318
rect 8300 26308 8352 26314
rect 8300 26250 8352 26256
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8208 25696 8260 25702
rect 8208 25638 8260 25644
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 8220 23882 8248 25638
rect 8312 25362 8340 26250
rect 8496 25702 8524 31146
rect 8588 28994 8616 40938
rect 8680 40662 8708 41550
rect 8668 40656 8720 40662
rect 8668 40598 8720 40604
rect 8680 38962 8708 40598
rect 8668 38956 8720 38962
rect 8668 38898 8720 38904
rect 8680 38554 8708 38898
rect 8668 38548 8720 38554
rect 8668 38490 8720 38496
rect 8772 36632 8800 41754
rect 8852 41676 8904 41682
rect 8852 41618 8904 41624
rect 9312 41676 9364 41682
rect 9312 41618 9364 41624
rect 8864 41070 8892 41618
rect 9220 41608 9272 41614
rect 9220 41550 9272 41556
rect 9232 41274 9260 41550
rect 9220 41268 9272 41274
rect 9220 41210 9272 41216
rect 9324 41070 9352 41618
rect 9416 41562 9444 42026
rect 9496 42016 9548 42022
rect 9496 41958 9548 41964
rect 9508 41682 9536 41958
rect 9496 41676 9548 41682
rect 9496 41618 9548 41624
rect 9416 41534 9536 41562
rect 8852 41064 8904 41070
rect 8852 41006 8904 41012
rect 9312 41064 9364 41070
rect 9312 41006 9364 41012
rect 9324 40594 9352 41006
rect 8944 40588 8996 40594
rect 8944 40530 8996 40536
rect 9312 40588 9364 40594
rect 9312 40530 9364 40536
rect 8852 40452 8904 40458
rect 8852 40394 8904 40400
rect 8864 38350 8892 40394
rect 8956 39302 8984 40530
rect 8944 39296 8996 39302
rect 8944 39238 8996 39244
rect 8956 38894 8984 39238
rect 8944 38888 8996 38894
rect 8944 38830 8996 38836
rect 8852 38344 8904 38350
rect 8852 38286 8904 38292
rect 8956 37806 8984 38830
rect 9324 38826 9352 40530
rect 9404 40112 9456 40118
rect 9404 40054 9456 40060
rect 9312 38820 9364 38826
rect 9312 38762 9364 38768
rect 9220 38480 9272 38486
rect 9220 38422 9272 38428
rect 9128 38412 9180 38418
rect 9128 38354 9180 38360
rect 8944 37800 8996 37806
rect 8944 37742 8996 37748
rect 9140 37466 9168 38354
rect 9128 37460 9180 37466
rect 9128 37402 9180 37408
rect 9232 36854 9260 38422
rect 9324 38418 9352 38762
rect 9312 38412 9364 38418
rect 9312 38354 9364 38360
rect 9324 36922 9352 38354
rect 9416 38010 9444 40054
rect 9508 39960 9536 41534
rect 9600 39960 9628 42026
rect 9680 42016 9732 42022
rect 9680 41958 9732 41964
rect 9692 41206 9720 41958
rect 9772 41744 9824 41750
rect 9772 41686 9824 41692
rect 9680 41200 9732 41206
rect 9680 41142 9732 41148
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 9496 39954 9548 39960
rect 9496 39896 9548 39902
rect 9588 39954 9640 39960
rect 9588 39896 9640 39902
rect 9508 38010 9536 39896
rect 9600 39642 9628 39896
rect 9588 39636 9640 39642
rect 9588 39578 9640 39584
rect 9692 38554 9720 39986
rect 9784 39098 9812 41686
rect 10060 41682 10088 42502
rect 10152 42158 10180 42502
rect 10244 42158 10272 42622
rect 10140 42152 10192 42158
rect 10140 42094 10192 42100
rect 10232 42152 10284 42158
rect 10232 42094 10284 42100
rect 10048 41676 10100 41682
rect 10048 41618 10100 41624
rect 10336 41614 10364 43318
rect 10520 42770 10548 44270
rect 10508 42764 10560 42770
rect 10508 42706 10560 42712
rect 10520 42106 10548 42706
rect 10612 42566 10640 44338
rect 10692 43648 10744 43654
rect 10692 43590 10744 43596
rect 10600 42560 10652 42566
rect 10600 42502 10652 42508
rect 10428 42078 10548 42106
rect 10428 41750 10456 42078
rect 10416 41744 10468 41750
rect 10416 41686 10468 41692
rect 10324 41608 10376 41614
rect 10324 41550 10376 41556
rect 10140 41540 10192 41546
rect 10140 41482 10192 41488
rect 9864 41472 9916 41478
rect 9864 41414 9916 41420
rect 9876 40526 9904 41414
rect 10152 41002 10180 41482
rect 10232 41064 10284 41070
rect 10232 41006 10284 41012
rect 10140 40996 10192 41002
rect 10140 40938 10192 40944
rect 10244 40730 10272 41006
rect 10232 40724 10284 40730
rect 10232 40666 10284 40672
rect 10336 40662 10364 41550
rect 10612 41546 10640 42502
rect 10704 42140 10732 43590
rect 10796 42634 10824 45222
rect 10876 44940 10928 44946
rect 10876 44882 10928 44888
rect 10888 43858 10916 44882
rect 10876 43852 10928 43858
rect 10876 43794 10928 43800
rect 10888 43246 10916 43794
rect 10876 43240 10928 43246
rect 10876 43182 10928 43188
rect 10980 42770 11008 45766
rect 11624 45558 11652 46922
rect 12176 46510 12204 46990
rect 12164 46504 12216 46510
rect 12164 46446 12216 46452
rect 12808 46504 12860 46510
rect 12808 46446 12860 46452
rect 11704 46368 11756 46374
rect 11704 46310 11756 46316
rect 11716 46034 11744 46310
rect 11704 46028 11756 46034
rect 11704 45970 11756 45976
rect 11612 45552 11664 45558
rect 11612 45494 11664 45500
rect 11980 45416 12032 45422
rect 11980 45358 12032 45364
rect 11253 45180 11561 45200
rect 11253 45178 11259 45180
rect 11315 45178 11339 45180
rect 11395 45178 11419 45180
rect 11475 45178 11499 45180
rect 11555 45178 11561 45180
rect 11315 45126 11317 45178
rect 11497 45126 11499 45178
rect 11253 45124 11259 45126
rect 11315 45124 11339 45126
rect 11395 45124 11419 45126
rect 11475 45124 11499 45126
rect 11555 45124 11561 45126
rect 11253 45104 11561 45124
rect 11152 45008 11204 45014
rect 11152 44950 11204 44956
rect 11060 43240 11112 43246
rect 11060 43182 11112 43188
rect 10968 42764 11020 42770
rect 10968 42706 11020 42712
rect 10784 42628 10836 42634
rect 10784 42570 10836 42576
rect 11072 42362 11100 43182
rect 11164 42702 11192 44950
rect 11612 44260 11664 44266
rect 11612 44202 11664 44208
rect 11253 44092 11561 44112
rect 11253 44090 11259 44092
rect 11315 44090 11339 44092
rect 11395 44090 11419 44092
rect 11475 44090 11499 44092
rect 11555 44090 11561 44092
rect 11315 44038 11317 44090
rect 11497 44038 11499 44090
rect 11253 44036 11259 44038
rect 11315 44036 11339 44038
rect 11395 44036 11419 44038
rect 11475 44036 11499 44038
rect 11555 44036 11561 44038
rect 11253 44016 11561 44036
rect 11624 43790 11652 44202
rect 11612 43784 11664 43790
rect 11612 43726 11664 43732
rect 11253 43004 11561 43024
rect 11253 43002 11259 43004
rect 11315 43002 11339 43004
rect 11395 43002 11419 43004
rect 11475 43002 11499 43004
rect 11555 43002 11561 43004
rect 11315 42950 11317 43002
rect 11497 42950 11499 43002
rect 11253 42948 11259 42950
rect 11315 42948 11339 42950
rect 11395 42948 11419 42950
rect 11475 42948 11499 42950
rect 11555 42948 11561 42950
rect 11253 42928 11561 42948
rect 11624 42770 11652 43726
rect 11704 43172 11756 43178
rect 11704 43114 11756 43120
rect 11612 42764 11664 42770
rect 11612 42706 11664 42712
rect 11152 42696 11204 42702
rect 11152 42638 11204 42644
rect 11060 42356 11112 42362
rect 11060 42298 11112 42304
rect 10784 42152 10836 42158
rect 10704 42112 10784 42140
rect 10784 42094 10836 42100
rect 10968 42016 11020 42022
rect 10968 41958 11020 41964
rect 10600 41540 10652 41546
rect 10600 41482 10652 41488
rect 10416 41472 10468 41478
rect 10416 41414 10468 41420
rect 10784 41472 10836 41478
rect 10784 41414 10836 41420
rect 10428 41070 10456 41414
rect 10416 41064 10468 41070
rect 10416 41006 10468 41012
rect 10600 41064 10652 41070
rect 10600 41006 10652 41012
rect 10692 41064 10744 41070
rect 10692 41006 10744 41012
rect 10324 40656 10376 40662
rect 10324 40598 10376 40604
rect 10140 40588 10192 40594
rect 10140 40530 10192 40536
rect 9864 40520 9916 40526
rect 9864 40462 9916 40468
rect 9772 39092 9824 39098
rect 9772 39034 9824 39040
rect 9876 39030 9904 40462
rect 10152 40118 10180 40530
rect 10324 40520 10376 40526
rect 10324 40462 10376 40468
rect 10232 40384 10284 40390
rect 10232 40326 10284 40332
rect 10140 40112 10192 40118
rect 10140 40054 10192 40060
rect 9864 39024 9916 39030
rect 9864 38966 9916 38972
rect 10048 38888 10100 38894
rect 10048 38830 10100 38836
rect 9956 38820 10008 38826
rect 9956 38762 10008 38768
rect 9680 38548 9732 38554
rect 9680 38490 9732 38496
rect 9968 38298 9996 38762
rect 10060 38418 10088 38830
rect 10048 38412 10100 38418
rect 10048 38354 10100 38360
rect 9588 38276 9640 38282
rect 9968 38270 10088 38298
rect 9588 38218 9640 38224
rect 9404 38004 9456 38010
rect 9404 37946 9456 37952
rect 9496 38004 9548 38010
rect 9496 37946 9548 37952
rect 9404 37460 9456 37466
rect 9404 37402 9456 37408
rect 9312 36916 9364 36922
rect 9312 36858 9364 36864
rect 9416 36854 9444 37402
rect 9220 36848 9272 36854
rect 9220 36790 9272 36796
rect 9404 36848 9456 36854
rect 9404 36790 9456 36796
rect 8772 36604 9076 36632
rect 8944 34944 8996 34950
rect 8944 34886 8996 34892
rect 8956 34610 8984 34886
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 8956 34490 8984 34546
rect 8864 34462 8984 34490
rect 8864 33998 8892 34462
rect 8944 34128 8996 34134
rect 8944 34070 8996 34076
rect 8852 33992 8904 33998
rect 8852 33934 8904 33940
rect 8956 33454 8984 34070
rect 8668 33448 8720 33454
rect 8668 33390 8720 33396
rect 8944 33448 8996 33454
rect 8944 33390 8996 33396
rect 8680 32502 8708 33390
rect 8760 32904 8812 32910
rect 8760 32846 8812 32852
rect 8668 32496 8720 32502
rect 8668 32438 8720 32444
rect 8680 31278 8708 32438
rect 8772 32026 8800 32846
rect 8760 32020 8812 32026
rect 8760 31962 8812 31968
rect 8956 31958 8984 33390
rect 8944 31952 8996 31958
rect 8944 31894 8996 31900
rect 8944 31476 8996 31482
rect 8944 31418 8996 31424
rect 8668 31272 8720 31278
rect 8668 31214 8720 31220
rect 8680 30394 8708 31214
rect 8956 30938 8984 31418
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 8668 30388 8720 30394
rect 8668 30330 8720 30336
rect 8680 30122 8708 30330
rect 8668 30116 8720 30122
rect 8668 30058 8720 30064
rect 8680 29714 8708 30058
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 8852 29504 8904 29510
rect 8852 29446 8904 29452
rect 8864 29102 8892 29446
rect 8852 29096 8904 29102
rect 8852 29038 8904 29044
rect 8588 28966 8708 28994
rect 8576 28620 8628 28626
rect 8576 28562 8628 28568
rect 8588 27538 8616 28562
rect 8576 27532 8628 27538
rect 8576 27474 8628 27480
rect 8484 25696 8536 25702
rect 8484 25638 8536 25644
rect 8484 25424 8536 25430
rect 8484 25366 8536 25372
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 8128 23854 8248 23882
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7668 22438 7696 22510
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7656 22432 7708 22438
rect 7656 22374 7708 22380
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7576 21486 7604 22374
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7668 21350 7696 22170
rect 7760 21894 7788 22442
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7392 19306 7512 19334
rect 7484 18850 7512 19306
rect 7392 18822 7512 18850
rect 7392 16794 7420 18822
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7484 18222 7512 18702
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7484 17134 7512 18158
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7576 16946 7604 20402
rect 7668 19990 7696 20538
rect 7656 19984 7708 19990
rect 7656 19926 7708 19932
rect 7760 19922 7788 21830
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 18970 7696 19246
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7656 18828 7708 18834
rect 7760 18816 7788 19858
rect 7852 18834 7880 23190
rect 8128 23118 8156 23854
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8036 21010 8064 22374
rect 8024 21004 8076 21010
rect 8024 20946 8076 20952
rect 7932 20392 7984 20398
rect 8036 20380 8064 20946
rect 8220 20584 8248 23734
rect 8312 22438 8340 25298
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8404 22642 8432 23462
rect 8496 23186 8524 25366
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 8496 22710 8524 23122
rect 8588 23118 8616 24142
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8312 21146 8340 22374
rect 8588 21842 8616 22918
rect 8496 21814 8616 21842
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8404 21010 8432 21286
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 8220 20556 8340 20584
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 7984 20352 8064 20380
rect 7932 20334 7984 20340
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 19922 7972 20198
rect 8036 19990 8064 20352
rect 8220 20058 8248 20402
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8024 19984 8076 19990
rect 8312 19938 8340 20556
rect 8496 20398 8524 21814
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8588 20244 8616 21626
rect 8024 19926 8076 19932
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 7708 18788 7788 18816
rect 7840 18828 7892 18834
rect 7656 18770 7708 18776
rect 7840 18770 7892 18776
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7852 17542 7880 18634
rect 7944 18222 7972 19858
rect 8036 19378 8064 19926
rect 8220 19910 8340 19938
rect 8404 20216 8616 20244
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8128 19174 8156 19790
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8220 18986 8248 19910
rect 8404 19802 8432 20216
rect 8128 18958 8248 18986
rect 8312 19774 8432 19802
rect 8484 19780 8536 19786
rect 8128 18902 8156 18958
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7944 17814 7972 18158
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7484 16918 7604 16946
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15026 7328 15302
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7116 14006 7144 14282
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6932 13326 6960 13806
rect 7116 13394 7144 13806
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6932 12918 6960 13262
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6102 11996 6410 12016
rect 6102 11994 6108 11996
rect 6164 11994 6188 11996
rect 6244 11994 6268 11996
rect 6324 11994 6348 11996
rect 6404 11994 6410 11996
rect 6164 11942 6166 11994
rect 6346 11942 6348 11994
rect 6102 11940 6108 11942
rect 6164 11940 6188 11942
rect 6244 11940 6268 11942
rect 6324 11940 6348 11942
rect 6404 11940 6410 11942
rect 6102 11920 6410 11940
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5920 11070 6040 11098
rect 6104 11082 6132 11698
rect 6472 11642 6500 12718
rect 6656 12306 6684 12718
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6380 11614 6500 11642
rect 6380 11098 6408 11614
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 11286 6500 11494
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6460 11144 6512 11150
rect 6380 11092 6460 11098
rect 6380 11086 6512 11092
rect 6012 11014 6040 11070
rect 6092 11076 6144 11082
rect 6380 11070 6500 11086
rect 6092 11018 6144 11024
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5920 10742 5948 10950
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5460 9846 5580 9874
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5460 8616 5488 9846
rect 5644 9518 5672 9862
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5368 8588 5488 8616
rect 5368 8362 5396 8588
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 7818 5396 8298
rect 5552 7886 5580 8910
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5368 7002 5396 7346
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5460 6866 5488 7482
rect 5264 6860 5316 6866
rect 5448 6860 5500 6866
rect 5264 6802 5316 6808
rect 5368 6820 5448 6848
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5000 4672 5028 5714
rect 5092 5556 5120 6190
rect 5184 5914 5212 6734
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5368 5778 5396 6820
rect 5448 6802 5500 6808
rect 5552 6254 5580 7686
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5644 6186 5672 9318
rect 5828 9042 5856 10610
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5828 8634 5856 8978
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5920 8430 5948 10406
rect 6012 9654 6040 10950
rect 6102 10908 6410 10928
rect 6102 10906 6108 10908
rect 6164 10906 6188 10908
rect 6244 10906 6268 10908
rect 6324 10906 6348 10908
rect 6404 10906 6410 10908
rect 6164 10854 6166 10906
rect 6346 10854 6348 10906
rect 6102 10852 6108 10854
rect 6164 10852 6188 10854
rect 6244 10852 6268 10854
rect 6324 10852 6348 10854
rect 6404 10852 6410 10854
rect 6102 10832 6410 10852
rect 6184 10600 6236 10606
rect 6472 10588 6500 11070
rect 6552 10600 6604 10606
rect 6472 10560 6552 10588
rect 6184 10542 6236 10548
rect 6552 10542 6604 10548
rect 6196 9908 6224 10542
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6472 10198 6500 10406
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6196 9880 6500 9908
rect 6102 9820 6410 9840
rect 6102 9818 6108 9820
rect 6164 9818 6188 9820
rect 6244 9818 6268 9820
rect 6324 9818 6348 9820
rect 6404 9818 6410 9820
rect 6164 9766 6166 9818
rect 6346 9766 6348 9818
rect 6102 9764 6108 9766
rect 6164 9764 6188 9766
rect 6244 9764 6268 9766
rect 6324 9764 6348 9766
rect 6404 9764 6410 9766
rect 6102 9744 6410 9764
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 9042 6408 9318
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6472 8974 6500 9880
rect 6564 9450 6592 10542
rect 6748 10470 6776 11222
rect 6932 10674 6960 12854
rect 7116 12714 7144 13330
rect 7208 12782 7236 14826
rect 7392 14414 7420 15506
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7484 13716 7512 16918
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7576 15502 7604 15846
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7576 14482 7604 14826
rect 7668 14618 7696 15982
rect 7852 15162 7880 17478
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7760 14498 7788 14894
rect 7840 14544 7892 14550
rect 7760 14492 7840 14498
rect 7760 14486 7892 14492
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7760 14470 7880 14486
rect 7576 13870 7604 14418
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7484 13688 7604 13716
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7208 12306 7236 12718
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11218 7052 11698
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6840 10266 6868 10542
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6840 9586 6868 10202
rect 7024 9722 7052 10406
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 7208 9110 7236 12242
rect 7300 11694 7328 13126
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7392 9654 7420 12174
rect 7484 11286 7512 12582
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7392 9450 7420 9590
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6102 8732 6410 8752
rect 6102 8730 6108 8732
rect 6164 8730 6188 8732
rect 6244 8730 6268 8732
rect 6324 8730 6348 8732
rect 6404 8730 6410 8732
rect 6164 8678 6166 8730
rect 6346 8678 6348 8730
rect 6102 8676 6108 8678
rect 6164 8676 6188 8678
rect 6244 8676 6268 8678
rect 6324 8676 6348 8678
rect 6404 8676 6410 8678
rect 6102 8656 6410 8676
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5920 8072 5948 8366
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5736 8044 5948 8072
rect 5736 7342 5764 8044
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 7002 5764 7142
rect 5828 7002 5856 7890
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5724 6860 5776 6866
rect 5776 6820 5856 6848
rect 5724 6802 5776 6808
rect 5828 6730 5856 6820
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5460 5914 5488 6054
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5172 5568 5224 5574
rect 5092 5528 5172 5556
rect 5172 5510 5224 5516
rect 5184 5370 5212 5510
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 4684 5132 4690
rect 5000 4644 5080 4672
rect 5080 4626 5132 4632
rect 5184 4604 5212 5306
rect 5368 5030 5396 5578
rect 5736 5166 5764 6258
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5264 4616 5316 4622
rect 5184 4576 5264 4604
rect 5264 4558 5316 4564
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4172 2650 4200 3130
rect 5368 3058 5396 4966
rect 5644 4622 5672 5034
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4078 5580 4422
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5828 3670 5856 6666
rect 5920 6390 5948 7822
rect 6012 7478 6040 8230
rect 6102 7644 6410 7664
rect 6102 7642 6108 7644
rect 6164 7642 6188 7644
rect 6244 7642 6268 7644
rect 6324 7642 6348 7644
rect 6404 7642 6410 7644
rect 6164 7590 6166 7642
rect 6346 7590 6348 7642
rect 6102 7588 6108 7590
rect 6164 7588 6188 7590
rect 6244 7588 6268 7590
rect 6324 7588 6348 7590
rect 6404 7588 6410 7590
rect 6102 7568 6410 7588
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 6730 6132 7278
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 6012 6254 6040 6598
rect 6102 6556 6410 6576
rect 6102 6554 6108 6556
rect 6164 6554 6188 6556
rect 6244 6554 6268 6556
rect 6324 6554 6348 6556
rect 6404 6554 6410 6556
rect 6164 6502 6166 6554
rect 6346 6502 6348 6554
rect 6102 6500 6108 6502
rect 6164 6500 6188 6502
rect 6244 6500 6268 6502
rect 6324 6500 6348 6502
rect 6404 6500 6410 6502
rect 6102 6480 6410 6500
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5098 6040 5646
rect 6102 5468 6410 5488
rect 6102 5466 6108 5468
rect 6164 5466 6188 5468
rect 6244 5466 6268 5468
rect 6324 5466 6348 5468
rect 6404 5466 6410 5468
rect 6164 5414 6166 5466
rect 6346 5414 6348 5466
rect 6102 5412 6108 5414
rect 6164 5412 6188 5414
rect 6244 5412 6268 5414
rect 6324 5412 6348 5414
rect 6404 5412 6410 5414
rect 6102 5392 6410 5412
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6472 4554 6500 8910
rect 6840 8566 6868 8978
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 7116 8430 7144 8774
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6564 7546 6592 7754
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6656 7478 6684 7754
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6656 7274 6684 7414
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6748 5846 6776 7958
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6102 4380 6410 4400
rect 6102 4378 6108 4380
rect 6164 4378 6188 4380
rect 6244 4378 6268 4380
rect 6324 4378 6348 4380
rect 6404 4378 6410 4380
rect 6164 4326 6166 4378
rect 6346 4326 6348 4378
rect 6102 4324 6108 4326
rect 6164 4324 6188 4326
rect 6244 4324 6268 4326
rect 6324 4324 6348 4326
rect 6404 4324 6410 4326
rect 6102 4304 6410 4324
rect 6748 3738 6776 5782
rect 6840 5166 6868 7890
rect 7576 7834 7604 13688
rect 7760 13530 7788 14470
rect 7944 14278 7972 15506
rect 8036 14822 8064 18770
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8128 18426 8156 18566
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8220 18086 8248 18770
rect 8312 18154 8340 19774
rect 8484 19722 8536 19728
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8220 17882 8248 18022
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8312 16250 8340 18090
rect 8404 17882 8432 19314
rect 8496 18222 8524 19722
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8496 17338 8524 18158
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8208 16108 8260 16114
rect 8260 16068 8340 16096
rect 8208 16050 8260 16056
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 14006 7972 14214
rect 8036 14006 8064 14758
rect 8128 14482 8156 15506
rect 8312 15502 8340 16068
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8404 15706 8432 15982
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8128 14074 8156 14418
rect 8220 14414 8248 14894
rect 8496 14482 8524 15574
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 14074 8248 14350
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 8128 13394 8156 14010
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7668 11558 7696 12650
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10198 7696 10406
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7668 9042 7696 9998
rect 7852 9926 7880 12718
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 12374 7972 12582
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 10266 8524 11494
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7668 8412 7696 8978
rect 8404 8634 8432 9522
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 7748 8424 7800 8430
rect 7668 8384 7748 8412
rect 7748 8366 7800 8372
rect 7484 7806 7604 7834
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7342 6960 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6932 5030 6960 5646
rect 7024 5642 7052 7278
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7116 5778 7144 7142
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4690 6960 4966
rect 7116 4826 7144 5034
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4282 6960 4626
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 7300 3942 7328 7482
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 6102 3292 6410 3312
rect 6102 3290 6108 3292
rect 6164 3290 6188 3292
rect 6244 3290 6268 3292
rect 6324 3290 6348 3292
rect 6404 3290 6410 3292
rect 6164 3238 6166 3290
rect 6346 3238 6348 3290
rect 6102 3236 6108 3238
rect 6164 3236 6188 3238
rect 6244 3236 6268 3238
rect 6324 3236 6348 3238
rect 6404 3236 6410 3238
rect 6102 3216 6410 3236
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5460 2650 5488 3130
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 5460 2038 5488 2586
rect 6012 2106 6040 2858
rect 7116 2650 7144 3674
rect 7300 3194 7328 3878
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6102 2204 6410 2224
rect 6102 2202 6108 2204
rect 6164 2202 6188 2204
rect 6244 2202 6268 2204
rect 6324 2202 6348 2204
rect 6404 2202 6410 2204
rect 6164 2150 6166 2202
rect 6346 2150 6348 2202
rect 6102 2148 6108 2150
rect 6164 2148 6188 2150
rect 6244 2148 6268 2150
rect 6324 2148 6348 2150
rect 6404 2148 6410 2150
rect 6102 2128 6410 2148
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 2964 1352 3016 1358
rect 2964 1294 3016 1300
rect 7392 1290 7420 3606
rect 7484 3534 7512 7806
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 6322 7604 7686
rect 7760 6730 7788 8366
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8036 7002 8064 7142
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7760 5778 7788 6666
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 5846 8064 6054
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7760 5234 7788 5714
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7760 4690 7788 5170
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7760 4214 7788 4626
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 8312 4146 8340 7754
rect 8404 7410 8432 7890
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7944 3738 7972 4014
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3058 7512 3470
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 8404 2038 8432 6802
rect 8588 4468 8616 19654
rect 8680 17814 8708 28966
rect 8852 28756 8904 28762
rect 8852 28698 8904 28704
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8772 26586 8800 27270
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8772 26450 8800 26522
rect 8760 26444 8812 26450
rect 8760 26386 8812 26392
rect 8772 24750 8800 26386
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8760 22568 8812 22574
rect 8760 22510 8812 22516
rect 8772 19718 8800 22510
rect 8864 21894 8892 28698
rect 9048 28098 9076 36604
rect 9232 36242 9260 36790
rect 9404 36712 9456 36718
rect 9600 36700 9628 38218
rect 10060 38214 10088 38270
rect 10048 38208 10100 38214
rect 10048 38150 10100 38156
rect 10060 37738 10088 38150
rect 10048 37732 10100 37738
rect 10048 37674 10100 37680
rect 9956 37460 10008 37466
rect 9956 37402 10008 37408
rect 9772 37324 9824 37330
rect 9772 37266 9824 37272
rect 9784 36922 9812 37266
rect 9772 36916 9824 36922
rect 9772 36858 9824 36864
rect 9456 36672 9628 36700
rect 9404 36654 9456 36660
rect 9220 36236 9272 36242
rect 9220 36178 9272 36184
rect 9220 36100 9272 36106
rect 9220 36042 9272 36048
rect 9232 35494 9260 36042
rect 9416 35494 9444 36654
rect 9496 35760 9548 35766
rect 9496 35702 9548 35708
rect 9220 35488 9272 35494
rect 9220 35430 9272 35436
rect 9404 35488 9456 35494
rect 9404 35430 9456 35436
rect 9232 34950 9260 35430
rect 9404 35216 9456 35222
rect 9404 35158 9456 35164
rect 9220 34944 9272 34950
rect 9220 34886 9272 34892
rect 9232 34490 9260 34886
rect 9140 34462 9260 34490
rect 9312 34536 9364 34542
rect 9312 34478 9364 34484
rect 9140 34134 9168 34462
rect 9220 34400 9272 34406
rect 9220 34342 9272 34348
rect 9128 34128 9180 34134
rect 9128 34070 9180 34076
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9140 32570 9168 33934
rect 9232 33454 9260 34342
rect 9324 34202 9352 34478
rect 9312 34196 9364 34202
rect 9312 34138 9364 34144
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 9128 32564 9180 32570
rect 9128 32506 9180 32512
rect 9232 32450 9260 33390
rect 9312 33380 9364 33386
rect 9312 33322 9364 33328
rect 9324 32978 9352 33322
rect 9312 32972 9364 32978
rect 9312 32914 9364 32920
rect 9416 32858 9444 35158
rect 9140 32422 9260 32450
rect 9324 32830 9444 32858
rect 9140 31346 9168 32422
rect 9220 32360 9272 32366
rect 9220 32302 9272 32308
rect 9232 31754 9260 32302
rect 9220 31748 9272 31754
rect 9220 31690 9272 31696
rect 9324 31498 9352 32830
rect 9404 32768 9456 32774
rect 9404 32710 9456 32716
rect 9232 31470 9352 31498
rect 9128 31340 9180 31346
rect 9128 31282 9180 31288
rect 8956 28070 9076 28098
rect 8956 23254 8984 28070
rect 9036 28008 9088 28014
rect 9036 27950 9088 27956
rect 9048 26926 9076 27950
rect 9036 26920 9088 26926
rect 9036 26862 9088 26868
rect 9048 25906 9076 26862
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 9048 24614 9076 25230
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9048 23730 9076 24550
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9140 23594 9168 31282
rect 9232 28762 9260 31470
rect 9416 31362 9444 32710
rect 9508 31906 9536 35702
rect 9680 34672 9732 34678
rect 9680 34614 9732 34620
rect 9588 33856 9640 33862
rect 9588 33798 9640 33804
rect 9600 32366 9628 33798
rect 9692 33454 9720 34614
rect 9772 33856 9824 33862
rect 9772 33798 9824 33804
rect 9784 33522 9812 33798
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9680 33448 9732 33454
rect 9680 33390 9732 33396
rect 9968 33046 9996 37402
rect 10060 33590 10088 37674
rect 10244 36174 10272 40326
rect 10336 40186 10364 40462
rect 10612 40390 10640 41006
rect 10704 40458 10732 41006
rect 10692 40452 10744 40458
rect 10692 40394 10744 40400
rect 10600 40384 10652 40390
rect 10600 40326 10652 40332
rect 10324 40180 10376 40186
rect 10324 40122 10376 40128
rect 10704 39914 10732 40394
rect 10796 39982 10824 41414
rect 10876 40928 10928 40934
rect 10876 40870 10928 40876
rect 10784 39976 10836 39982
rect 10784 39918 10836 39924
rect 10692 39908 10744 39914
rect 10692 39850 10744 39856
rect 10416 39500 10468 39506
rect 10416 39442 10468 39448
rect 10428 38418 10456 39442
rect 10416 38412 10468 38418
rect 10416 38354 10468 38360
rect 10428 37806 10456 38354
rect 10416 37800 10468 37806
rect 10416 37742 10468 37748
rect 10784 37664 10836 37670
rect 10784 37606 10836 37612
rect 10600 37120 10652 37126
rect 10600 37062 10652 37068
rect 10416 36644 10468 36650
rect 10416 36586 10468 36592
rect 10324 36372 10376 36378
rect 10324 36314 10376 36320
rect 10232 36168 10284 36174
rect 10232 36110 10284 36116
rect 10336 35698 10364 36314
rect 10428 36310 10456 36586
rect 10612 36378 10640 37062
rect 10796 36650 10824 37606
rect 10888 37330 10916 40870
rect 10980 40526 11008 41958
rect 11253 41916 11561 41936
rect 11253 41914 11259 41916
rect 11315 41914 11339 41916
rect 11395 41914 11419 41916
rect 11475 41914 11499 41916
rect 11555 41914 11561 41916
rect 11315 41862 11317 41914
rect 11497 41862 11499 41914
rect 11253 41860 11259 41862
rect 11315 41860 11339 41862
rect 11395 41860 11419 41862
rect 11475 41860 11499 41862
rect 11555 41860 11561 41862
rect 11253 41840 11561 41860
rect 11624 41138 11652 42706
rect 11060 41132 11112 41138
rect 11060 41074 11112 41080
rect 11612 41132 11664 41138
rect 11612 41074 11664 41080
rect 10968 40520 11020 40526
rect 10968 40462 11020 40468
rect 10968 38412 11020 38418
rect 10968 38354 11020 38360
rect 10980 37670 11008 38354
rect 10968 37664 11020 37670
rect 10968 37606 11020 37612
rect 11072 37398 11100 41074
rect 11253 40828 11561 40848
rect 11253 40826 11259 40828
rect 11315 40826 11339 40828
rect 11395 40826 11419 40828
rect 11475 40826 11499 40828
rect 11555 40826 11561 40828
rect 11315 40774 11317 40826
rect 11497 40774 11499 40826
rect 11253 40772 11259 40774
rect 11315 40772 11339 40774
rect 11395 40772 11419 40774
rect 11475 40772 11499 40774
rect 11555 40772 11561 40774
rect 11253 40752 11561 40772
rect 11428 40384 11480 40390
rect 11428 40326 11480 40332
rect 11440 39982 11468 40326
rect 11428 39976 11480 39982
rect 11428 39918 11480 39924
rect 11253 39740 11561 39760
rect 11253 39738 11259 39740
rect 11315 39738 11339 39740
rect 11395 39738 11419 39740
rect 11475 39738 11499 39740
rect 11555 39738 11561 39740
rect 11315 39686 11317 39738
rect 11497 39686 11499 39738
rect 11253 39684 11259 39686
rect 11315 39684 11339 39686
rect 11395 39684 11419 39686
rect 11475 39684 11499 39686
rect 11555 39684 11561 39686
rect 11253 39664 11561 39684
rect 11152 39500 11204 39506
rect 11152 39442 11204 39448
rect 11164 38826 11192 39442
rect 11152 38820 11204 38826
rect 11152 38762 11204 38768
rect 11164 38554 11192 38762
rect 11253 38652 11561 38672
rect 11716 38654 11744 43114
rect 11796 43104 11848 43110
rect 11796 43046 11848 43052
rect 11808 42838 11836 43046
rect 11796 42832 11848 42838
rect 11796 42774 11848 42780
rect 11888 42356 11940 42362
rect 11888 42298 11940 42304
rect 11796 38752 11848 38758
rect 11796 38694 11848 38700
rect 11253 38650 11259 38652
rect 11315 38650 11339 38652
rect 11395 38650 11419 38652
rect 11475 38650 11499 38652
rect 11555 38650 11561 38652
rect 11315 38598 11317 38650
rect 11497 38598 11499 38650
rect 11253 38596 11259 38598
rect 11315 38596 11339 38598
rect 11395 38596 11419 38598
rect 11475 38596 11499 38598
rect 11555 38596 11561 38598
rect 11253 38576 11561 38596
rect 11624 38626 11744 38654
rect 11152 38548 11204 38554
rect 11152 38490 11204 38496
rect 11152 37936 11204 37942
rect 11152 37878 11204 37884
rect 11164 37806 11192 37878
rect 11152 37800 11204 37806
rect 11152 37742 11204 37748
rect 11253 37564 11561 37584
rect 11253 37562 11259 37564
rect 11315 37562 11339 37564
rect 11395 37562 11419 37564
rect 11475 37562 11499 37564
rect 11555 37562 11561 37564
rect 11315 37510 11317 37562
rect 11497 37510 11499 37562
rect 11253 37508 11259 37510
rect 11315 37508 11339 37510
rect 11395 37508 11419 37510
rect 11475 37508 11499 37510
rect 11555 37508 11561 37510
rect 11253 37488 11561 37508
rect 11060 37392 11112 37398
rect 11060 37334 11112 37340
rect 10876 37324 10928 37330
rect 10876 37266 10928 37272
rect 11152 37324 11204 37330
rect 11152 37266 11204 37272
rect 11060 36712 11112 36718
rect 11060 36654 11112 36660
rect 10784 36644 10836 36650
rect 10784 36586 10836 36592
rect 10600 36372 10652 36378
rect 10600 36314 10652 36320
rect 10416 36304 10468 36310
rect 10416 36246 10468 36252
rect 10324 35692 10376 35698
rect 10324 35634 10376 35640
rect 10140 35624 10192 35630
rect 10140 35566 10192 35572
rect 10232 35624 10284 35630
rect 10232 35566 10284 35572
rect 10152 35494 10180 35566
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 10152 34746 10180 35430
rect 10244 35290 10272 35566
rect 10232 35284 10284 35290
rect 10232 35226 10284 35232
rect 10232 35148 10284 35154
rect 10232 35090 10284 35096
rect 10140 34740 10192 34746
rect 10140 34682 10192 34688
rect 10244 33998 10272 35090
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 10336 33930 10364 35634
rect 10428 35630 10456 36246
rect 10416 35624 10468 35630
rect 10416 35566 10468 35572
rect 10600 35556 10652 35562
rect 10600 35498 10652 35504
rect 10416 35488 10468 35494
rect 10416 35430 10468 35436
rect 10428 35222 10456 35430
rect 10416 35216 10468 35222
rect 10416 35158 10468 35164
rect 10324 33924 10376 33930
rect 10324 33866 10376 33872
rect 10048 33584 10100 33590
rect 10048 33526 10100 33532
rect 9864 33040 9916 33046
rect 9864 32982 9916 32988
rect 9956 33040 10008 33046
rect 9956 32982 10008 32988
rect 9680 32904 9732 32910
rect 9680 32846 9732 32852
rect 9692 32570 9720 32846
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9588 32360 9640 32366
rect 9588 32302 9640 32308
rect 9876 32298 9904 32982
rect 9864 32292 9916 32298
rect 9864 32234 9916 32240
rect 9508 31878 9628 31906
rect 9496 31816 9548 31822
rect 9496 31758 9548 31764
rect 9324 31334 9444 31362
rect 9220 28756 9272 28762
rect 9220 28698 9272 28704
rect 9220 28416 9272 28422
rect 9220 28358 9272 28364
rect 9232 26858 9260 28358
rect 9324 27826 9352 31334
rect 9404 31272 9456 31278
rect 9508 31260 9536 31758
rect 9456 31232 9536 31260
rect 9404 31214 9456 31220
rect 9416 30122 9444 31214
rect 9404 30116 9456 30122
rect 9404 30058 9456 30064
rect 9496 30116 9548 30122
rect 9496 30058 9548 30064
rect 9416 29646 9444 30058
rect 9508 29850 9536 30058
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 9600 29782 9628 31878
rect 9588 29776 9640 29782
rect 9588 29718 9640 29724
rect 9404 29640 9456 29646
rect 9404 29582 9456 29588
rect 9416 28014 9444 29582
rect 9680 29028 9732 29034
rect 9680 28970 9732 28976
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9508 28558 9536 28902
rect 9692 28626 9720 28970
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 9508 27878 9536 28494
rect 9496 27872 9548 27878
rect 9324 27798 9444 27826
rect 9496 27814 9548 27820
rect 9220 26852 9272 26858
rect 9220 26794 9272 26800
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9324 25838 9352 26182
rect 9312 25832 9364 25838
rect 9312 25774 9364 25780
rect 9220 24064 9272 24070
rect 9220 24006 9272 24012
rect 9232 23662 9260 24006
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9128 23588 9180 23594
rect 9128 23530 9180 23536
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 8956 22094 8984 23190
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 8956 22066 9076 22094
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8864 20602 8892 21830
rect 8956 21622 8984 21966
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8956 20398 8984 20946
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8864 19310 8892 20198
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8772 18630 8800 19110
rect 8956 18766 8984 20334
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 8668 17808 8720 17814
rect 8668 17750 8720 17756
rect 8680 15026 8708 17750
rect 8864 16590 8892 18362
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8772 14890 8800 16186
rect 8864 16046 8892 16390
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8864 15162 8892 15438
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8956 14618 8984 16594
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8772 13870 8800 14282
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8680 6322 8708 13738
rect 8772 12306 8800 13806
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8772 11354 8800 12242
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 7954 8892 10542
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7478 8892 7890
rect 8956 7546 8984 8978
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8680 5846 8708 6258
rect 8864 6254 8892 7414
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 5914 8800 6122
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8496 4440 8616 4468
rect 8496 3670 8524 4440
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8496 3194 8524 3606
rect 8588 3398 8616 4014
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8588 2650 8616 3334
rect 9048 3126 9076 22066
rect 9140 21962 9168 22646
rect 9128 21956 9180 21962
rect 9128 21898 9180 21904
rect 9140 21554 9168 21898
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9128 21412 9180 21418
rect 9232 21400 9260 23598
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9324 22778 9352 23122
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9416 22094 9444 27798
rect 9508 27402 9536 27814
rect 9692 27674 9720 28562
rect 9876 28490 9904 32234
rect 10336 31890 10364 33866
rect 10416 32972 10468 32978
rect 10416 32914 10468 32920
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10336 29306 10364 29786
rect 10324 29300 10376 29306
rect 10324 29242 10376 29248
rect 9864 28484 9916 28490
rect 9864 28426 9916 28432
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10244 28014 10272 28358
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 9496 27396 9548 27402
rect 9496 27338 9548 27344
rect 10244 27130 10272 27474
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 9496 26444 9548 26450
rect 9496 26386 9548 26392
rect 9508 25430 9536 26386
rect 9496 25424 9548 25430
rect 9496 25366 9548 25372
rect 9680 25424 9732 25430
rect 9680 25366 9732 25372
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9600 24818 9628 25298
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 9508 24342 9536 24686
rect 9496 24336 9548 24342
rect 9496 24278 9548 24284
rect 9600 24274 9628 24754
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9508 22234 9536 23122
rect 9692 22710 9720 25366
rect 9772 25220 9824 25226
rect 9772 25162 9824 25168
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9416 22066 9536 22094
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9180 21372 9260 21400
rect 9128 21354 9180 21360
rect 9140 21146 9168 21354
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9140 18970 9168 19858
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 9140 9518 9168 18294
rect 9232 16794 9260 20878
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9232 15502 9260 16526
rect 9324 16182 9352 21490
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9416 19378 9444 19654
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9416 18426 9444 18702
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9508 18358 9536 22066
rect 9600 21554 9628 22374
rect 9692 22094 9720 22646
rect 9784 22574 9812 25162
rect 10244 24750 10272 27066
rect 10428 25786 10456 32914
rect 10508 32496 10560 32502
rect 10508 32438 10560 32444
rect 10520 30122 10548 32438
rect 10612 32314 10640 35498
rect 10876 35488 10928 35494
rect 10876 35430 10928 35436
rect 10692 34944 10744 34950
rect 10692 34886 10744 34892
rect 10704 34746 10732 34886
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 10888 34474 10916 35430
rect 11072 35154 11100 36654
rect 11164 35562 11192 37266
rect 11253 36476 11561 36496
rect 11253 36474 11259 36476
rect 11315 36474 11339 36476
rect 11395 36474 11419 36476
rect 11475 36474 11499 36476
rect 11555 36474 11561 36476
rect 11315 36422 11317 36474
rect 11497 36422 11499 36474
rect 11253 36420 11259 36422
rect 11315 36420 11339 36422
rect 11395 36420 11419 36422
rect 11475 36420 11499 36422
rect 11555 36420 11561 36422
rect 11253 36400 11561 36420
rect 11152 35556 11204 35562
rect 11152 35498 11204 35504
rect 11253 35388 11561 35408
rect 11253 35386 11259 35388
rect 11315 35386 11339 35388
rect 11395 35386 11419 35388
rect 11475 35386 11499 35388
rect 11555 35386 11561 35388
rect 11315 35334 11317 35386
rect 11497 35334 11499 35386
rect 11253 35332 11259 35334
rect 11315 35332 11339 35334
rect 11395 35332 11419 35334
rect 11475 35332 11499 35334
rect 11555 35332 11561 35334
rect 11253 35312 11561 35332
rect 11624 35306 11652 38626
rect 11704 38412 11756 38418
rect 11704 38354 11756 38360
rect 11716 37806 11744 38354
rect 11808 37942 11836 38694
rect 11900 37942 11928 42298
rect 11992 39982 12020 45358
rect 12072 44464 12124 44470
rect 12072 44406 12124 44412
rect 12084 42158 12112 44406
rect 12176 44334 12204 46446
rect 12624 46368 12676 46374
rect 12624 46310 12676 46316
rect 12636 46034 12664 46310
rect 12820 46034 12848 46446
rect 12624 46028 12676 46034
rect 12624 45970 12676 45976
rect 12808 46028 12860 46034
rect 12808 45970 12860 45976
rect 12912 45966 12940 47602
rect 13084 47592 13136 47598
rect 13084 47534 13136 47540
rect 13728 47592 13780 47598
rect 13728 47534 13780 47540
rect 14372 47592 14424 47598
rect 14372 47534 14424 47540
rect 13096 46050 13124 47534
rect 13544 47456 13596 47462
rect 13544 47398 13596 47404
rect 13360 47116 13412 47122
rect 13360 47058 13412 47064
rect 13372 46170 13400 47058
rect 13556 46918 13584 47398
rect 13544 46912 13596 46918
rect 13544 46854 13596 46860
rect 13556 46578 13584 46854
rect 13544 46572 13596 46578
rect 13544 46514 13596 46520
rect 13740 46374 13768 47534
rect 13820 47524 13872 47530
rect 13820 47466 13872 47472
rect 13832 46714 13860 47466
rect 14384 46918 14412 47534
rect 15752 47524 15804 47530
rect 15752 47466 15804 47472
rect 15384 47252 15436 47258
rect 15384 47194 15436 47200
rect 14372 46912 14424 46918
rect 14372 46854 14424 46860
rect 13820 46708 13872 46714
rect 13820 46650 13872 46656
rect 13728 46368 13780 46374
rect 13728 46310 13780 46316
rect 13360 46164 13412 46170
rect 13360 46106 13412 46112
rect 13004 46022 13124 46050
rect 13740 46034 13768 46310
rect 13728 46028 13780 46034
rect 13004 45966 13032 46022
rect 13648 45988 13728 46016
rect 12900 45960 12952 45966
rect 12900 45902 12952 45908
rect 12992 45960 13044 45966
rect 12992 45902 13044 45908
rect 12912 45778 12940 45902
rect 13084 45892 13136 45898
rect 13084 45834 13136 45840
rect 13096 45778 13124 45834
rect 12912 45750 13124 45778
rect 12912 45490 12940 45750
rect 12900 45484 12952 45490
rect 12900 45426 12952 45432
rect 12532 45416 12584 45422
rect 12532 45358 12584 45364
rect 12348 44804 12400 44810
rect 12348 44746 12400 44752
rect 12360 44334 12388 44746
rect 12164 44328 12216 44334
rect 12164 44270 12216 44276
rect 12348 44328 12400 44334
rect 12348 44270 12400 44276
rect 12256 44192 12308 44198
rect 12256 44134 12308 44140
rect 12268 43926 12296 44134
rect 12256 43920 12308 43926
rect 12256 43862 12308 43868
rect 12544 43314 12572 45358
rect 13648 45082 13676 45988
rect 13728 45970 13780 45976
rect 13728 45892 13780 45898
rect 13728 45834 13780 45840
rect 13740 45626 13768 45834
rect 13728 45620 13780 45626
rect 13728 45562 13780 45568
rect 13832 45422 13860 46650
rect 14384 46510 14412 46854
rect 14372 46504 14424 46510
rect 14372 46446 14424 46452
rect 14096 46436 14148 46442
rect 14096 46378 14148 46384
rect 13912 45892 13964 45898
rect 13912 45834 13964 45840
rect 13820 45416 13872 45422
rect 13820 45358 13872 45364
rect 13924 45354 13952 45834
rect 14108 45490 14136 46378
rect 14188 45960 14240 45966
rect 14188 45902 14240 45908
rect 14200 45830 14228 45902
rect 14188 45824 14240 45830
rect 14188 45766 14240 45772
rect 14200 45642 14228 45766
rect 14200 45614 14320 45642
rect 14292 45558 14320 45614
rect 14188 45552 14240 45558
rect 14188 45494 14240 45500
rect 14280 45552 14332 45558
rect 14280 45494 14332 45500
rect 14096 45484 14148 45490
rect 14096 45426 14148 45432
rect 13912 45348 13964 45354
rect 13912 45290 13964 45296
rect 13636 45076 13688 45082
rect 13636 45018 13688 45024
rect 13648 44946 13676 45018
rect 13636 44940 13688 44946
rect 13636 44882 13688 44888
rect 12624 44872 12676 44878
rect 12624 44814 12676 44820
rect 13452 44872 13504 44878
rect 13452 44814 13504 44820
rect 12532 43308 12584 43314
rect 12532 43250 12584 43256
rect 12544 43194 12572 43250
rect 12452 43166 12572 43194
rect 12636 43178 12664 44814
rect 12624 43172 12676 43178
rect 12072 42152 12124 42158
rect 12072 42094 12124 42100
rect 12256 40996 12308 41002
rect 12256 40938 12308 40944
rect 12268 40730 12296 40938
rect 12256 40724 12308 40730
rect 12256 40666 12308 40672
rect 12072 40452 12124 40458
rect 12072 40394 12124 40400
rect 11980 39976 12032 39982
rect 11980 39918 12032 39924
rect 11796 37936 11848 37942
rect 11796 37878 11848 37884
rect 11888 37936 11940 37942
rect 11888 37878 11940 37884
rect 11704 37800 11756 37806
rect 11704 37742 11756 37748
rect 11704 37664 11756 37670
rect 11704 37606 11756 37612
rect 11716 35578 11744 37606
rect 11808 36310 11836 37878
rect 11888 37800 11940 37806
rect 11888 37742 11940 37748
rect 11900 36922 11928 37742
rect 11992 37652 12020 39918
rect 12084 39828 12112 40394
rect 12452 40050 12480 43166
rect 12624 43114 12676 43120
rect 13268 43172 13320 43178
rect 13268 43114 13320 43120
rect 12992 42764 13044 42770
rect 12992 42706 13044 42712
rect 13004 42090 13032 42706
rect 13280 42566 13308 43114
rect 13464 42702 13492 44814
rect 13912 44260 13964 44266
rect 13912 44202 13964 44208
rect 13452 42696 13504 42702
rect 13452 42638 13504 42644
rect 13268 42560 13320 42566
rect 13268 42502 13320 42508
rect 13084 42220 13136 42226
rect 13084 42162 13136 42168
rect 12992 42084 13044 42090
rect 12992 42026 13044 42032
rect 12532 41812 12584 41818
rect 12532 41754 12584 41760
rect 12544 40458 12572 41754
rect 12808 41676 12860 41682
rect 12808 41618 12860 41624
rect 12624 41608 12676 41614
rect 12624 41550 12676 41556
rect 12636 40526 12664 41550
rect 12820 41206 12848 41618
rect 12808 41200 12860 41206
rect 12808 41142 12860 41148
rect 12820 40594 12848 41142
rect 13004 40594 13032 42026
rect 13096 41682 13124 42162
rect 13084 41676 13136 41682
rect 13084 41618 13136 41624
rect 13280 41414 13308 42502
rect 13360 42152 13412 42158
rect 13360 42094 13412 42100
rect 13372 41682 13400 42094
rect 13360 41676 13412 41682
rect 13360 41618 13412 41624
rect 13280 41386 13400 41414
rect 13084 41064 13136 41070
rect 13084 41006 13136 41012
rect 12808 40588 12860 40594
rect 12808 40530 12860 40536
rect 12992 40588 13044 40594
rect 12992 40530 13044 40536
rect 13096 40526 13124 41006
rect 12624 40520 12676 40526
rect 12624 40462 12676 40468
rect 13084 40520 13136 40526
rect 13084 40462 13136 40468
rect 12532 40452 12584 40458
rect 12532 40394 12584 40400
rect 12636 40050 12664 40462
rect 12440 40044 12492 40050
rect 12440 39986 12492 39992
rect 12624 40044 12676 40050
rect 12624 39986 12676 39992
rect 12084 39800 12204 39828
rect 12072 37936 12124 37942
rect 12072 37878 12124 37884
rect 12084 37806 12112 37878
rect 12072 37800 12124 37806
rect 12072 37742 12124 37748
rect 11992 37624 12112 37652
rect 11888 36916 11940 36922
rect 11888 36858 11940 36864
rect 11796 36304 11848 36310
rect 11796 36246 11848 36252
rect 11900 35698 11928 36858
rect 11980 36032 12032 36038
rect 11980 35974 12032 35980
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11992 35630 12020 35974
rect 11980 35624 12032 35630
rect 11716 35550 11928 35578
rect 11980 35566 12032 35572
rect 11624 35278 11836 35306
rect 11704 35216 11756 35222
rect 11704 35158 11756 35164
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 10876 34468 10928 34474
rect 10876 34410 10928 34416
rect 10692 33448 10744 33454
rect 10692 33390 10744 33396
rect 10704 33114 10732 33390
rect 10692 33108 10744 33114
rect 10692 33050 10744 33056
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 10796 32366 10824 32710
rect 11072 32502 11100 35090
rect 11253 34300 11561 34320
rect 11253 34298 11259 34300
rect 11315 34298 11339 34300
rect 11395 34298 11419 34300
rect 11475 34298 11499 34300
rect 11555 34298 11561 34300
rect 11315 34246 11317 34298
rect 11497 34246 11499 34298
rect 11253 34244 11259 34246
rect 11315 34244 11339 34246
rect 11395 34244 11419 34246
rect 11475 34244 11499 34246
rect 11555 34244 11561 34246
rect 11253 34224 11561 34244
rect 11520 33856 11572 33862
rect 11520 33798 11572 33804
rect 11152 33516 11204 33522
rect 11152 33458 11204 33464
rect 11164 32774 11192 33458
rect 11532 33402 11560 33798
rect 11532 33374 11652 33402
rect 11253 33212 11561 33232
rect 11253 33210 11259 33212
rect 11315 33210 11339 33212
rect 11395 33210 11419 33212
rect 11475 33210 11499 33212
rect 11555 33210 11561 33212
rect 11315 33158 11317 33210
rect 11497 33158 11499 33210
rect 11253 33156 11259 33158
rect 11315 33156 11339 33158
rect 11395 33156 11419 33158
rect 11475 33156 11499 33158
rect 11555 33156 11561 33158
rect 11253 33136 11561 33156
rect 11624 33114 11652 33374
rect 11716 33114 11744 35158
rect 11808 33658 11836 35278
rect 11796 33652 11848 33658
rect 11796 33594 11848 33600
rect 11808 33454 11836 33594
rect 11796 33448 11848 33454
rect 11796 33390 11848 33396
rect 11900 33130 11928 35550
rect 12084 35222 12112 37624
rect 12176 37074 12204 39800
rect 12452 39574 12480 39986
rect 12440 39568 12492 39574
rect 12440 39510 12492 39516
rect 12440 39432 12492 39438
rect 12440 39374 12492 39380
rect 12452 38962 12480 39374
rect 12440 38956 12492 38962
rect 12440 38898 12492 38904
rect 12452 38350 12480 38898
rect 12532 38548 12584 38554
rect 12532 38490 12584 38496
rect 12440 38344 12492 38350
rect 12440 38286 12492 38292
rect 12452 37874 12480 38286
rect 12440 37868 12492 37874
rect 12440 37810 12492 37816
rect 12348 37664 12400 37670
rect 12348 37606 12400 37612
rect 12360 37330 12388 37606
rect 12348 37324 12400 37330
rect 12348 37266 12400 37272
rect 12176 37046 12296 37074
rect 12268 35894 12296 37046
rect 12544 36786 12572 38490
rect 12636 38418 12664 39986
rect 12992 39976 13044 39982
rect 12992 39918 13044 39924
rect 12624 38412 12676 38418
rect 12624 38354 12676 38360
rect 12808 37936 12860 37942
rect 12808 37878 12860 37884
rect 12716 37868 12768 37874
rect 12716 37810 12768 37816
rect 12624 37800 12676 37806
rect 12624 37742 12676 37748
rect 12636 37466 12664 37742
rect 12624 37460 12676 37466
rect 12624 37402 12676 37408
rect 12532 36780 12584 36786
rect 12532 36722 12584 36728
rect 12636 36718 12664 37402
rect 12728 36718 12756 37810
rect 12820 36786 12848 37878
rect 13004 37806 13032 39918
rect 13096 39030 13124 40462
rect 13084 39024 13136 39030
rect 13084 38966 13136 38972
rect 13096 38350 13124 38966
rect 13372 38894 13400 41386
rect 13464 39846 13492 42638
rect 13728 42016 13780 42022
rect 13728 41958 13780 41964
rect 13740 40662 13768 41958
rect 13820 41268 13872 41274
rect 13820 41210 13872 41216
rect 13832 40730 13860 41210
rect 13820 40724 13872 40730
rect 13820 40666 13872 40672
rect 13728 40656 13780 40662
rect 13728 40598 13780 40604
rect 13544 40588 13596 40594
rect 13544 40530 13596 40536
rect 13556 39914 13584 40530
rect 13544 39908 13596 39914
rect 13544 39850 13596 39856
rect 13452 39840 13504 39846
rect 13452 39782 13504 39788
rect 13728 39840 13780 39846
rect 13728 39782 13780 39788
rect 13740 39438 13768 39782
rect 13832 39506 13860 40666
rect 13820 39500 13872 39506
rect 13820 39442 13872 39448
rect 13452 39432 13504 39438
rect 13452 39374 13504 39380
rect 13728 39432 13780 39438
rect 13728 39374 13780 39380
rect 13176 38888 13228 38894
rect 13176 38830 13228 38836
rect 13360 38888 13412 38894
rect 13360 38830 13412 38836
rect 13084 38344 13136 38350
rect 13084 38286 13136 38292
rect 12992 37800 13044 37806
rect 12992 37742 13044 37748
rect 12992 37664 13044 37670
rect 12992 37606 13044 37612
rect 12900 36848 12952 36854
rect 12900 36790 12952 36796
rect 12808 36780 12860 36786
rect 12808 36722 12860 36728
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12716 36712 12768 36718
rect 12716 36654 12768 36660
rect 12268 35866 12388 35894
rect 12164 35488 12216 35494
rect 12164 35430 12216 35436
rect 12072 35216 12124 35222
rect 12072 35158 12124 35164
rect 12176 35154 12204 35430
rect 12164 35148 12216 35154
rect 12164 35090 12216 35096
rect 12164 34604 12216 34610
rect 12164 34546 12216 34552
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 11992 33522 12020 33934
rect 12084 33862 12112 34342
rect 12072 33856 12124 33862
rect 12072 33798 12124 33804
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 12084 33402 12112 33798
rect 11612 33108 11664 33114
rect 11612 33050 11664 33056
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 11808 33102 11928 33130
rect 11992 33374 12112 33402
rect 11612 32972 11664 32978
rect 11612 32914 11664 32920
rect 11152 32768 11204 32774
rect 11152 32710 11204 32716
rect 11060 32496 11112 32502
rect 11060 32438 11112 32444
rect 10968 32428 11020 32434
rect 10968 32370 11020 32376
rect 10784 32360 10836 32366
rect 10612 32286 10732 32314
rect 10784 32302 10836 32308
rect 10876 32360 10928 32366
rect 10876 32302 10928 32308
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10612 31958 10640 32166
rect 10600 31952 10652 31958
rect 10600 31894 10652 31900
rect 10704 31906 10732 32286
rect 10796 32026 10824 32302
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10704 31878 10824 31906
rect 10692 31816 10744 31822
rect 10692 31758 10744 31764
rect 10508 30116 10560 30122
rect 10508 30058 10560 30064
rect 10600 29844 10652 29850
rect 10600 29786 10652 29792
rect 10612 29714 10640 29786
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10600 29708 10652 29714
rect 10600 29650 10652 29656
rect 10520 29306 10548 29650
rect 10600 29572 10652 29578
rect 10600 29514 10652 29520
rect 10508 29300 10560 29306
rect 10508 29242 10560 29248
rect 10612 29170 10640 29514
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10612 28694 10640 29106
rect 10600 28688 10652 28694
rect 10600 28630 10652 28636
rect 10612 27062 10640 28630
rect 10600 27056 10652 27062
rect 10600 26998 10652 27004
rect 10612 26382 10640 26998
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10428 25758 10548 25786
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 10428 25430 10456 25638
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 10416 24948 10468 24954
rect 10416 24890 10468 24896
rect 10324 24880 10376 24886
rect 10324 24822 10376 24828
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 9968 24274 9996 24686
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 9968 24154 9996 24210
rect 9876 24126 9996 24154
rect 9876 23662 9904 24126
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9968 22642 9996 24006
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10060 22778 10088 23122
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9772 22568 9824 22574
rect 9824 22528 9904 22556
rect 9772 22510 9824 22516
rect 9692 22066 9812 22094
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9784 21010 9812 22066
rect 9876 21418 9904 22528
rect 9968 22098 9996 22578
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10244 22098 10272 22510
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 9864 21412 9916 21418
rect 9864 21354 9916 21360
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9968 20534 9996 20810
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9784 19378 9812 19654
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9416 17338 9444 17614
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9416 16658 9444 17274
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9416 12102 9444 16594
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9232 11218 9260 12038
rect 9508 11898 9536 18090
rect 9876 17814 9904 18226
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9600 15638 9628 17478
rect 9968 17338 9996 17682
rect 10060 17678 10088 18022
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9876 16794 9904 17138
rect 9968 17134 9996 17274
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9968 16522 9996 17070
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9692 15706 9720 15982
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9600 13870 9628 15302
rect 10060 15094 10088 15982
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9600 12782 9628 13806
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9600 11898 9628 12582
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9692 10606 9720 14894
rect 9784 14890 9812 14962
rect 10152 14958 10180 21490
rect 10244 21486 10272 22034
rect 10232 21480 10284 21486
rect 10232 21422 10284 21428
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10244 16726 10272 18294
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10244 16114 10272 16662
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 10152 14618 10180 14894
rect 10140 14612 10192 14618
rect 10060 14572 10140 14600
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9876 13530 9904 13738
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9968 13394 9996 13670
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 11694 9812 12582
rect 10060 12442 10088 14572
rect 10140 14554 10192 14560
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9968 10742 9996 11630
rect 10060 11354 10088 12378
rect 10244 11830 10272 16050
rect 10336 15162 10364 24822
rect 10428 23526 10456 24890
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10428 22098 10456 23462
rect 10520 23050 10548 25758
rect 10612 25430 10640 26318
rect 10600 25424 10652 25430
rect 10600 25366 10652 25372
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10612 24070 10640 24754
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10508 23044 10560 23050
rect 10508 22986 10560 22992
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10428 19922 10456 20198
rect 10520 20058 10548 22986
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10612 21554 10640 21966
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10520 18630 10548 19246
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10428 17746 10456 18158
rect 10520 17814 10548 18566
rect 10612 17882 10640 18906
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10416 17604 10468 17610
rect 10416 17546 10468 17552
rect 10428 16590 10456 17546
rect 10520 17112 10548 17750
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10508 17106 10560 17112
rect 10508 17048 10560 17054
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10520 16454 10548 17048
rect 10612 16794 10640 17478
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10704 16640 10732 31758
rect 10796 24886 10824 31878
rect 10888 29578 10916 32302
rect 10980 31822 11008 32370
rect 11152 32360 11204 32366
rect 11152 32302 11204 32308
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10968 31408 11020 31414
rect 10968 31350 11020 31356
rect 10876 29572 10928 29578
rect 10876 29514 10928 29520
rect 10876 29096 10928 29102
rect 10980 29084 11008 31350
rect 11072 31278 11100 31962
rect 11164 31890 11192 32302
rect 11253 32124 11561 32144
rect 11253 32122 11259 32124
rect 11315 32122 11339 32124
rect 11395 32122 11419 32124
rect 11475 32122 11499 32124
rect 11555 32122 11561 32124
rect 11315 32070 11317 32122
rect 11497 32070 11499 32122
rect 11253 32068 11259 32070
rect 11315 32068 11339 32070
rect 11395 32068 11419 32070
rect 11475 32068 11499 32070
rect 11555 32068 11561 32070
rect 11253 32048 11561 32068
rect 11152 31884 11204 31890
rect 11152 31826 11204 31832
rect 11624 31414 11652 32914
rect 11704 31816 11756 31822
rect 11704 31758 11756 31764
rect 11612 31408 11664 31414
rect 11612 31350 11664 31356
rect 11716 31278 11744 31758
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 11704 31272 11756 31278
rect 11704 31214 11756 31220
rect 11612 31136 11664 31142
rect 11612 31078 11664 31084
rect 11253 31036 11561 31056
rect 11253 31034 11259 31036
rect 11315 31034 11339 31036
rect 11395 31034 11419 31036
rect 11475 31034 11499 31036
rect 11555 31034 11561 31036
rect 11315 30982 11317 31034
rect 11497 30982 11499 31034
rect 11253 30980 11259 30982
rect 11315 30980 11339 30982
rect 11395 30980 11419 30982
rect 11475 30980 11499 30982
rect 11555 30980 11561 30982
rect 11253 30960 11561 30980
rect 11152 30184 11204 30190
rect 11152 30126 11204 30132
rect 11164 29850 11192 30126
rect 11253 29948 11561 29968
rect 11253 29946 11259 29948
rect 11315 29946 11339 29948
rect 11395 29946 11419 29948
rect 11475 29946 11499 29948
rect 11555 29946 11561 29948
rect 11315 29894 11317 29946
rect 11497 29894 11499 29946
rect 11253 29892 11259 29894
rect 11315 29892 11339 29894
rect 11395 29892 11419 29894
rect 11475 29892 11499 29894
rect 11555 29892 11561 29894
rect 11253 29872 11561 29892
rect 11152 29844 11204 29850
rect 11152 29786 11204 29792
rect 11060 29096 11112 29102
rect 10980 29056 11060 29084
rect 10876 29038 10928 29044
rect 11060 29038 11112 29044
rect 10888 28490 10916 29038
rect 11164 29034 11192 29786
rect 11624 29730 11652 31078
rect 11716 30802 11744 31214
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 11808 29782 11836 33102
rect 11888 32292 11940 32298
rect 11888 32234 11940 32240
rect 11900 32026 11928 32234
rect 11888 32020 11940 32026
rect 11888 31962 11940 31968
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11336 29708 11388 29714
rect 11336 29650 11388 29656
rect 11532 29702 11652 29730
rect 11796 29776 11848 29782
rect 11796 29718 11848 29724
rect 11704 29708 11756 29714
rect 11348 29102 11376 29650
rect 11428 29572 11480 29578
rect 11428 29514 11480 29520
rect 11440 29306 11468 29514
rect 11428 29300 11480 29306
rect 11428 29242 11480 29248
rect 11336 29096 11388 29102
rect 11336 29038 11388 29044
rect 11152 29028 11204 29034
rect 11152 28970 11204 28976
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 10980 28626 11008 28902
rect 11072 28762 11100 28902
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 10968 28620 11020 28626
rect 10968 28562 11020 28568
rect 10876 28484 10928 28490
rect 10876 28426 10928 28432
rect 10980 27606 11008 28562
rect 11072 28218 11100 28698
rect 11164 28694 11192 28970
rect 11532 28948 11560 29702
rect 11704 29650 11756 29656
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11624 29016 11652 29582
rect 11716 29306 11744 29650
rect 11704 29300 11756 29306
rect 11704 29242 11756 29248
rect 11900 29238 11928 29990
rect 11888 29232 11940 29238
rect 11888 29174 11940 29180
rect 11624 28988 11928 29016
rect 11532 28920 11744 28948
rect 11253 28860 11561 28880
rect 11253 28858 11259 28860
rect 11315 28858 11339 28860
rect 11395 28858 11419 28860
rect 11475 28858 11499 28860
rect 11555 28858 11561 28860
rect 11315 28806 11317 28858
rect 11497 28806 11499 28858
rect 11253 28804 11259 28806
rect 11315 28804 11339 28806
rect 11395 28804 11419 28806
rect 11475 28804 11499 28806
rect 11555 28804 11561 28806
rect 11253 28784 11561 28804
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 11072 26994 11100 28154
rect 11152 27940 11204 27946
rect 11152 27882 11204 27888
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 11164 26926 11192 27882
rect 11253 27772 11561 27792
rect 11253 27770 11259 27772
rect 11315 27770 11339 27772
rect 11395 27770 11419 27772
rect 11475 27770 11499 27772
rect 11555 27770 11561 27772
rect 11315 27718 11317 27770
rect 11497 27718 11499 27770
rect 11253 27716 11259 27718
rect 11315 27716 11339 27718
rect 11395 27716 11419 27718
rect 11475 27716 11499 27718
rect 11555 27716 11561 27718
rect 11253 27696 11561 27716
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 11256 26926 11284 27542
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11060 26852 11112 26858
rect 11060 26794 11112 26800
rect 11072 26330 11100 26794
rect 11256 26772 11284 26862
rect 11164 26744 11284 26772
rect 11164 26450 11192 26744
rect 11253 26684 11561 26704
rect 11253 26682 11259 26684
rect 11315 26682 11339 26684
rect 11395 26682 11419 26684
rect 11475 26682 11499 26684
rect 11555 26682 11561 26684
rect 11315 26630 11317 26682
rect 11497 26630 11499 26682
rect 11253 26628 11259 26630
rect 11315 26628 11339 26630
rect 11395 26628 11419 26630
rect 11475 26628 11499 26630
rect 11555 26628 11561 26630
rect 11253 26608 11561 26628
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 11520 26444 11572 26450
rect 11520 26386 11572 26392
rect 11072 26302 11192 26330
rect 10876 25968 10928 25974
rect 10876 25910 10928 25916
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10796 24274 10824 24550
rect 10784 24268 10836 24274
rect 10784 24210 10836 24216
rect 10796 21978 10824 24210
rect 10888 22778 10916 25910
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11072 25362 11100 25638
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 10968 24744 11020 24750
rect 10968 24686 11020 24692
rect 10980 24342 11008 24686
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 11072 24274 11100 25298
rect 11164 24750 11192 26302
rect 11532 26246 11560 26386
rect 11520 26240 11572 26246
rect 11716 26234 11744 28920
rect 11900 28762 11928 28988
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11808 28422 11836 28494
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11888 28416 11940 28422
rect 11992 28404 12020 33374
rect 12072 33108 12124 33114
rect 12072 33050 12124 33056
rect 12084 29510 12112 33050
rect 12176 31754 12204 34546
rect 12256 33448 12308 33454
rect 12256 33390 12308 33396
rect 12268 32978 12296 33390
rect 12256 32972 12308 32978
rect 12256 32914 12308 32920
rect 12176 31726 12296 31754
rect 12164 31680 12216 31686
rect 12164 31622 12216 31628
rect 12176 31346 12204 31622
rect 12164 31340 12216 31346
rect 12164 31282 12216 31288
rect 12176 30598 12204 31282
rect 12164 30592 12216 30598
rect 12164 30534 12216 30540
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 12072 29504 12124 29510
rect 12072 29446 12124 29452
rect 12072 29232 12124 29238
rect 12072 29174 12124 29180
rect 12084 28626 12112 29174
rect 12072 28620 12124 28626
rect 12072 28562 12124 28568
rect 12176 28558 12204 30194
rect 12268 29050 12296 31726
rect 12360 31142 12388 35866
rect 12636 35562 12664 36654
rect 12912 36106 12940 36790
rect 12900 36100 12952 36106
rect 12900 36042 12952 36048
rect 12624 35556 12676 35562
rect 12624 35498 12676 35504
rect 12636 34678 12664 35498
rect 13004 35290 13032 37606
rect 13096 37398 13124 38286
rect 13188 37942 13216 38830
rect 13464 38826 13492 39374
rect 13452 38820 13504 38826
rect 13452 38762 13504 38768
rect 13464 38554 13492 38762
rect 13452 38548 13504 38554
rect 13452 38490 13504 38496
rect 13176 37936 13228 37942
rect 13176 37878 13228 37884
rect 13176 37800 13228 37806
rect 13176 37742 13228 37748
rect 13084 37392 13136 37398
rect 13084 37334 13136 37340
rect 13096 36718 13124 37334
rect 13084 36712 13136 36718
rect 13084 36654 13136 36660
rect 13096 36242 13124 36654
rect 13084 36236 13136 36242
rect 13084 36178 13136 36184
rect 12992 35284 13044 35290
rect 12992 35226 13044 35232
rect 13188 35170 13216 37742
rect 13268 36576 13320 36582
rect 13268 36518 13320 36524
rect 13280 36242 13308 36518
rect 13268 36236 13320 36242
rect 13268 36178 13320 36184
rect 13728 36032 13780 36038
rect 13728 35974 13780 35980
rect 13452 35692 13504 35698
rect 13452 35634 13504 35640
rect 13004 35142 13216 35170
rect 12624 34672 12676 34678
rect 12624 34614 12676 34620
rect 13004 34474 13032 35142
rect 13360 34944 13412 34950
rect 13360 34886 13412 34892
rect 13372 34474 13400 34886
rect 13464 34626 13492 35634
rect 13544 35556 13596 35562
rect 13544 35498 13596 35504
rect 13556 34746 13584 35498
rect 13544 34740 13596 34746
rect 13544 34682 13596 34688
rect 13740 34678 13768 35974
rect 13728 34672 13780 34678
rect 13464 34598 13584 34626
rect 13728 34614 13780 34620
rect 12992 34468 13044 34474
rect 12992 34410 13044 34416
rect 13360 34468 13412 34474
rect 13360 34410 13412 34416
rect 13452 34468 13504 34474
rect 13452 34410 13504 34416
rect 12808 34128 12860 34134
rect 12808 34070 12860 34076
rect 12532 33040 12584 33046
rect 12532 32982 12584 32988
rect 12544 32842 12572 32982
rect 12716 32972 12768 32978
rect 12716 32914 12768 32920
rect 12532 32836 12584 32842
rect 12532 32778 12584 32784
rect 12544 31414 12572 32778
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12636 31890 12664 32302
rect 12624 31884 12676 31890
rect 12624 31826 12676 31832
rect 12532 31408 12584 31414
rect 12532 31350 12584 31356
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12348 30796 12400 30802
rect 12348 30738 12400 30744
rect 12360 29578 12388 30738
rect 12452 30734 12480 31214
rect 12544 31124 12572 31350
rect 12636 31278 12664 31826
rect 12728 31686 12756 32914
rect 12716 31680 12768 31686
rect 12716 31622 12768 31628
rect 12624 31272 12676 31278
rect 12624 31214 12676 31220
rect 12544 31096 12664 31124
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12440 30388 12492 30394
rect 12440 30330 12492 30336
rect 12348 29572 12400 29578
rect 12348 29514 12400 29520
rect 12360 29170 12388 29514
rect 12348 29164 12400 29170
rect 12348 29106 12400 29112
rect 12268 29022 12388 29050
rect 12256 28960 12308 28966
rect 12256 28902 12308 28908
rect 12268 28626 12296 28902
rect 12256 28620 12308 28626
rect 12256 28562 12308 28568
rect 12164 28552 12216 28558
rect 12164 28494 12216 28500
rect 12360 28490 12388 29022
rect 12348 28484 12400 28490
rect 12348 28426 12400 28432
rect 11992 28376 12296 28404
rect 11888 28358 11940 28364
rect 11808 27878 11836 28358
rect 11796 27872 11848 27878
rect 11796 27814 11848 27820
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 26518 11836 26862
rect 11900 26858 11928 28358
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11992 27130 12020 27474
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11796 26512 11848 26518
rect 11796 26454 11848 26460
rect 11900 26450 11928 26794
rect 11992 26450 12020 26862
rect 11888 26444 11940 26450
rect 11888 26386 11940 26392
rect 11980 26444 12032 26450
rect 11980 26386 12032 26392
rect 11520 26182 11572 26188
rect 11624 26206 11744 26234
rect 11253 25596 11561 25616
rect 11253 25594 11259 25596
rect 11315 25594 11339 25596
rect 11395 25594 11419 25596
rect 11475 25594 11499 25596
rect 11555 25594 11561 25596
rect 11315 25542 11317 25594
rect 11497 25542 11499 25594
rect 11253 25540 11259 25542
rect 11315 25540 11339 25542
rect 11395 25540 11419 25542
rect 11475 25540 11499 25542
rect 11555 25540 11561 25542
rect 11253 25520 11561 25540
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11348 24750 11376 24890
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11164 24410 11192 24686
rect 11253 24508 11561 24528
rect 11253 24506 11259 24508
rect 11315 24506 11339 24508
rect 11395 24506 11419 24508
rect 11475 24506 11499 24508
rect 11555 24506 11561 24508
rect 11315 24454 11317 24506
rect 11497 24454 11499 24506
rect 11253 24452 11259 24454
rect 11315 24452 11339 24454
rect 11395 24452 11419 24454
rect 11475 24452 11499 24454
rect 11555 24452 11561 24454
rect 11253 24432 11561 24452
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 11072 22642 11100 24006
rect 11532 23594 11560 24210
rect 11624 24138 11652 26206
rect 11992 25974 12020 26386
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 11980 25968 12032 25974
rect 11980 25910 12032 25916
rect 11992 25362 12020 25910
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 12084 25294 12112 26182
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 12084 24682 12112 25230
rect 12072 24676 12124 24682
rect 12072 24618 12124 24624
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11612 24132 11664 24138
rect 11612 24074 11664 24080
rect 11716 23662 11744 24550
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11253 23420 11561 23440
rect 11253 23418 11259 23420
rect 11315 23418 11339 23420
rect 11395 23418 11419 23420
rect 11475 23418 11499 23420
rect 11555 23418 11561 23420
rect 11315 23366 11317 23418
rect 11497 23366 11499 23418
rect 11253 23364 11259 23366
rect 11315 23364 11339 23366
rect 11395 23364 11419 23366
rect 11475 23364 11499 23366
rect 11555 23364 11561 23366
rect 11253 23344 11561 23364
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10796 21950 10916 21978
rect 10888 21486 10916 21950
rect 10980 21554 11008 22510
rect 11072 22234 11100 22578
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11253 22332 11561 22352
rect 11253 22330 11259 22332
rect 11315 22330 11339 22332
rect 11395 22330 11419 22332
rect 11475 22330 11499 22332
rect 11555 22330 11561 22332
rect 11315 22278 11317 22330
rect 11497 22278 11499 22330
rect 11253 22276 11259 22278
rect 11315 22276 11339 22278
rect 11395 22276 11419 22278
rect 11475 22276 11499 22278
rect 11555 22276 11561 22278
rect 11253 22256 11561 22276
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 11152 22160 11204 22166
rect 11152 22102 11204 22108
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10888 20806 10916 21422
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10888 19530 10916 20742
rect 10980 20534 11008 20946
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 11072 20398 11100 21966
rect 11164 21010 11192 22102
rect 11624 22098 11652 22510
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11253 21244 11561 21264
rect 11253 21242 11259 21244
rect 11315 21242 11339 21244
rect 11395 21242 11419 21244
rect 11475 21242 11499 21244
rect 11555 21242 11561 21244
rect 11315 21190 11317 21242
rect 11497 21190 11499 21242
rect 11253 21188 11259 21190
rect 11315 21188 11339 21190
rect 11395 21188 11419 21190
rect 11475 21188 11499 21190
rect 11555 21188 11561 21190
rect 11253 21168 11561 21188
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10612 16612 10732 16640
rect 10796 19502 10916 19530
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10336 13530 10364 15098
rect 10612 14618 10640 16612
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10704 15706 10732 16458
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10796 14890 10824 19502
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10888 18902 10916 19110
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10980 18834 11008 19994
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10888 17746 10916 18702
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10888 17202 10916 17546
rect 10980 17270 11008 18634
rect 11072 18426 11100 20334
rect 11164 19718 11192 20470
rect 11532 20398 11560 20946
rect 11716 20398 11744 21422
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11253 20156 11561 20176
rect 11253 20154 11259 20156
rect 11315 20154 11339 20156
rect 11395 20154 11419 20156
rect 11475 20154 11499 20156
rect 11555 20154 11561 20156
rect 11315 20102 11317 20154
rect 11497 20102 11499 20154
rect 11253 20100 11259 20102
rect 11315 20100 11339 20102
rect 11395 20100 11419 20102
rect 11475 20100 11499 20102
rect 11555 20100 11561 20102
rect 11253 20080 11561 20100
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11520 19304 11572 19310
rect 11624 19292 11652 20198
rect 11716 19446 11744 20334
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11572 19264 11652 19292
rect 11520 19246 11572 19252
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 18766 11192 19110
rect 11253 19068 11561 19088
rect 11253 19066 11259 19068
rect 11315 19066 11339 19068
rect 11395 19066 11419 19068
rect 11475 19066 11499 19068
rect 11555 19066 11561 19068
rect 11315 19014 11317 19066
rect 11497 19014 11499 19066
rect 11253 19012 11259 19014
rect 11315 19012 11339 19014
rect 11395 19012 11419 19014
rect 11475 19012 11499 19014
rect 11555 19012 11561 19014
rect 11253 18992 11561 19012
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 11256 18068 11284 18770
rect 11716 18222 11744 19382
rect 11808 19242 11836 24550
rect 11888 23656 11940 23662
rect 11888 23598 11940 23604
rect 11900 22574 11928 23598
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11900 20466 11928 21830
rect 11992 21622 12020 23462
rect 11980 21616 12032 21622
rect 11980 21558 12032 21564
rect 11992 20942 12020 21558
rect 12164 21412 12216 21418
rect 12164 21354 12216 21360
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11808 18086 11836 18838
rect 11164 18040 11284 18068
rect 11612 18080 11664 18086
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16726 11100 17070
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11072 16046 11100 16662
rect 11164 16164 11192 18040
rect 11612 18022 11664 18028
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11253 17980 11561 18000
rect 11253 17978 11259 17980
rect 11315 17978 11339 17980
rect 11395 17978 11419 17980
rect 11475 17978 11499 17980
rect 11555 17978 11561 17980
rect 11315 17926 11317 17978
rect 11497 17926 11499 17978
rect 11253 17924 11259 17926
rect 11315 17924 11339 17926
rect 11395 17924 11419 17926
rect 11475 17924 11499 17926
rect 11555 17924 11561 17926
rect 11253 17904 11561 17924
rect 11624 17882 11652 18022
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11624 17202 11652 17274
rect 11808 17218 11836 18022
rect 11900 17678 11928 20402
rect 11992 19922 12020 20742
rect 12072 20392 12124 20398
rect 12176 20380 12204 21354
rect 12124 20352 12204 20380
rect 12072 20334 12124 20340
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11716 17190 11836 17218
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11253 16892 11561 16912
rect 11253 16890 11259 16892
rect 11315 16890 11339 16892
rect 11395 16890 11419 16892
rect 11475 16890 11499 16892
rect 11555 16890 11561 16892
rect 11315 16838 11317 16890
rect 11497 16838 11499 16890
rect 11253 16836 11259 16838
rect 11315 16836 11339 16838
rect 11395 16836 11419 16838
rect 11475 16836 11499 16838
rect 11555 16836 11561 16838
rect 11253 16816 11561 16836
rect 11336 16176 11388 16182
rect 11164 16136 11336 16164
rect 11624 16130 11652 17138
rect 11716 16658 11744 17190
rect 11900 17116 11928 17206
rect 11992 17202 12020 19246
rect 12084 19242 12112 20334
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11808 17088 11928 17116
rect 12072 17128 12124 17134
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11808 16590 11836 17088
rect 12072 17070 12124 17076
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11336 16118 11388 16124
rect 11532 16102 11744 16130
rect 11808 16114 11836 16526
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11428 16040 11480 16046
rect 11532 16028 11560 16102
rect 11480 16000 11560 16028
rect 11428 15982 11480 15988
rect 11072 14958 11100 15982
rect 11253 15804 11561 15824
rect 11253 15802 11259 15804
rect 11315 15802 11339 15804
rect 11395 15802 11419 15804
rect 11475 15802 11499 15804
rect 11555 15802 11561 15804
rect 11315 15750 11317 15802
rect 11497 15750 11499 15802
rect 11253 15748 11259 15750
rect 11315 15748 11339 15750
rect 11395 15748 11419 15750
rect 11475 15748 11499 15750
rect 11555 15748 11561 15750
rect 11253 15728 11561 15748
rect 11716 15162 11744 16102
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11900 15638 11928 16934
rect 11992 16794 12020 16934
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10612 14074 10640 14554
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10336 12986 10364 13330
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10336 12646 10364 12922
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 12374 10364 12582
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10428 12306 10456 13670
rect 10612 13326 10640 14010
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10704 13394 10732 13874
rect 11072 13870 11100 14894
rect 11253 14716 11561 14736
rect 11253 14714 11259 14716
rect 11315 14714 11339 14716
rect 11395 14714 11419 14716
rect 11475 14714 11499 14716
rect 11555 14714 11561 14716
rect 11315 14662 11317 14714
rect 11497 14662 11499 14714
rect 11253 14660 11259 14662
rect 11315 14660 11339 14662
rect 11395 14660 11419 14662
rect 11475 14660 11499 14662
rect 11555 14660 11561 14662
rect 11253 14640 11561 14660
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11253 13628 11561 13648
rect 11253 13626 11259 13628
rect 11315 13626 11339 13628
rect 11395 13626 11419 13628
rect 11475 13626 11499 13628
rect 11555 13626 11561 13628
rect 11315 13574 11317 13626
rect 11497 13574 11499 13626
rect 11253 13572 11259 13574
rect 11315 13572 11339 13574
rect 11395 13572 11419 13574
rect 11475 13572 11499 13574
rect 11555 13572 11561 13574
rect 11253 13552 11561 13572
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 10600 13320 10652 13326
rect 10520 13268 10600 13274
rect 10520 13262 10652 13268
rect 10520 13246 10640 13262
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10336 11694 10364 12174
rect 10428 11762 10456 12242
rect 10520 12238 10548 13246
rect 10704 12782 10732 13330
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12782 11100 13262
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11164 12850 11192 13194
rect 11624 12986 11652 13330
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10692 12776 10744 12782
rect 10876 12776 10928 12782
rect 10692 12718 10744 12724
rect 10796 12736 10876 12764
rect 10704 12442 10732 12718
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10796 12306 10824 12736
rect 10876 12718 10928 12724
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10520 11914 10548 12174
rect 10520 11886 10640 11914
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10244 10810 10272 11562
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 9518 9352 10474
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9140 9110 9168 9454
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 8022 9168 8842
rect 9324 8022 9352 9454
rect 10152 9042 10180 10610
rect 10244 10266 10272 10746
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10336 9654 10364 11630
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10428 10742 10456 11086
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10428 10266 10456 10542
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10152 8634 10180 8978
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9600 8090 9628 8298
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9128 8016 9180 8022
rect 9312 8016 9364 8022
rect 9128 7958 9180 7964
rect 9232 7976 9312 8004
rect 9140 7342 9168 7958
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9232 7274 9260 7976
rect 9312 7958 9364 7964
rect 10048 7948 10100 7954
rect 10152 7936 10180 8570
rect 10244 8566 10272 8774
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10100 7908 10180 7936
rect 10048 7890 10100 7896
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 9324 7342 9352 7822
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7546 10272 7686
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9312 7336 9364 7342
rect 9496 7336 9548 7342
rect 9364 7296 9444 7324
rect 9312 7278 9364 7284
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9232 6458 9260 7210
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9232 6232 9260 6394
rect 9220 6226 9272 6232
rect 9416 6186 9444 7296
rect 9496 7278 9548 7284
rect 9508 7002 9536 7278
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9508 6254 9536 6938
rect 9600 6338 9628 7414
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6338 9720 6598
rect 9600 6310 9720 6338
rect 9876 6254 9904 6802
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9220 6168 9272 6174
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9140 4826 9168 5646
rect 9232 5166 9260 5850
rect 9416 5166 9444 6122
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9128 4820 9180 4826
rect 9180 4780 9260 4808
rect 9128 4762 9180 4768
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9140 4146 9168 4626
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9232 4078 9260 4780
rect 9416 4146 9444 5102
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 9600 2106 9628 5306
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9692 2650 9720 2926
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9588 2100 9640 2106
rect 9588 2042 9640 2048
rect 8392 2032 8444 2038
rect 8392 1974 8444 1980
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 9140 1562 9168 1974
rect 9692 1562 9720 2586
rect 9784 2514 9812 3606
rect 9876 3194 9904 5782
rect 9968 5778 9996 7210
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6254 10180 6598
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 10060 5710 10088 6122
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10244 5574 10272 6326
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4146 10272 4558
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9968 3602 9996 3946
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10060 3126 10088 4014
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3534 10180 3878
rect 10244 3602 10272 4082
rect 10336 4010 10364 7822
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10428 6254 10456 6394
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10244 3126 10272 3538
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10048 3120 10100 3126
rect 10232 3120 10284 3126
rect 10048 3062 10100 3068
rect 10152 3068 10232 3074
rect 10152 3062 10284 3068
rect 10152 3046 10272 3062
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10060 2038 10088 2926
rect 10152 2310 10180 3046
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10244 2446 10272 2926
rect 10336 2514 10364 3334
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 8392 1556 8444 1562
rect 8392 1498 8444 1504
rect 9128 1556 9180 1562
rect 9128 1498 9180 1504
rect 9680 1556 9732 1562
rect 9680 1498 9732 1504
rect 7380 1284 7432 1290
rect 7380 1226 7432 1232
rect 6102 1116 6410 1136
rect 6102 1114 6108 1116
rect 6164 1114 6188 1116
rect 6244 1114 6268 1116
rect 6324 1114 6348 1116
rect 6404 1114 6410 1116
rect 6164 1062 6166 1114
rect 6346 1062 6348 1114
rect 6102 1060 6108 1062
rect 6164 1060 6188 1062
rect 6244 1060 6268 1062
rect 6324 1060 6348 1062
rect 6404 1060 6410 1062
rect 6102 1040 6410 1060
rect 8404 1018 8432 1498
rect 10520 1340 10548 11766
rect 10612 11558 10640 11886
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10704 11150 10732 12174
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10796 10810 10824 12242
rect 11164 12238 11192 12786
rect 11253 12540 11561 12560
rect 11253 12538 11259 12540
rect 11315 12538 11339 12540
rect 11395 12538 11419 12540
rect 11475 12538 11499 12540
rect 11555 12538 11561 12540
rect 11315 12486 11317 12538
rect 11497 12486 11499 12538
rect 11253 12484 11259 12486
rect 11315 12484 11339 12486
rect 11395 12484 11419 12486
rect 11475 12484 11499 12486
rect 11555 12484 11561 12486
rect 11253 12464 11561 12484
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11253 11452 11561 11472
rect 11253 11450 11259 11452
rect 11315 11450 11339 11452
rect 11395 11450 11419 11452
rect 11475 11450 11499 11452
rect 11555 11450 11561 11452
rect 11315 11398 11317 11450
rect 11497 11398 11499 11450
rect 11253 11396 11259 11398
rect 11315 11396 11339 11398
rect 11395 11396 11419 11398
rect 11475 11396 11499 11398
rect 11555 11396 11561 11398
rect 11253 11376 11561 11396
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 11716 10606 11744 12038
rect 11808 11694 11836 12378
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 11218 11836 11494
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11900 10606 11928 13126
rect 11992 12434 12020 16594
rect 12084 16250 12112 17070
rect 12176 16658 12204 19110
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12072 16244 12124 16250
rect 12124 16204 12204 16232
rect 12072 16186 12124 16192
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 15570 12112 15982
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 14550 12112 15506
rect 12176 15366 12204 16204
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12268 14618 12296 28376
rect 12360 28014 12388 28426
rect 12348 28008 12400 28014
rect 12348 27950 12400 27956
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 12360 26382 12388 26794
rect 12452 26602 12480 30330
rect 12532 30116 12584 30122
rect 12532 30058 12584 30064
rect 12544 29306 12572 30058
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12636 28370 12664 31096
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 12728 29102 12756 29990
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12636 28342 12756 28370
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12452 26574 12572 26602
rect 12544 26518 12572 26574
rect 12532 26512 12584 26518
rect 12532 26454 12584 26460
rect 12348 26376 12400 26382
rect 12348 26318 12400 26324
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12452 25838 12480 26250
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12544 25650 12572 26250
rect 12452 25622 12572 25650
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12360 23798 12388 24686
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12360 18902 12388 23530
rect 12452 23186 12480 25622
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12544 24342 12572 24686
rect 12532 24336 12584 24342
rect 12532 24278 12584 24284
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12452 21010 12480 21830
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12452 20466 12480 20946
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12544 19530 12572 23666
rect 12636 20058 12664 27950
rect 12728 27826 12756 28342
rect 12820 27946 12848 34070
rect 13004 33862 13032 34410
rect 13464 34134 13492 34410
rect 13452 34128 13504 34134
rect 13452 34070 13504 34076
rect 13360 34060 13412 34066
rect 13360 34002 13412 34008
rect 12992 33856 13044 33862
rect 12992 33798 13044 33804
rect 13372 33658 13400 34002
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 13360 33652 13412 33658
rect 13360 33594 13412 33600
rect 12900 32836 12952 32842
rect 12900 32778 12952 32784
rect 12912 32502 12940 32778
rect 12992 32768 13044 32774
rect 12992 32710 13044 32716
rect 12900 32496 12952 32502
rect 12900 32438 12952 32444
rect 12912 31890 12940 32438
rect 12900 31884 12952 31890
rect 12900 31826 12952 31832
rect 13004 31754 13032 32710
rect 13188 32026 13216 33594
rect 13268 32904 13320 32910
rect 13268 32846 13320 32852
rect 13176 32020 13228 32026
rect 13176 31962 13228 31968
rect 12992 31748 13044 31754
rect 12992 31690 13044 31696
rect 13004 31362 13032 31690
rect 13188 31482 13216 31962
rect 13176 31476 13228 31482
rect 13176 31418 13228 31424
rect 12912 31334 13032 31362
rect 12912 30394 12940 31334
rect 12992 31204 13044 31210
rect 12992 31146 13044 31152
rect 12900 30388 12952 30394
rect 12900 30330 12952 30336
rect 12900 30184 12952 30190
rect 12900 30126 12952 30132
rect 12808 27940 12860 27946
rect 12808 27882 12860 27888
rect 12728 27798 12848 27826
rect 12716 26444 12768 26450
rect 12716 26386 12768 26392
rect 12728 25158 12756 26386
rect 12820 26042 12848 27798
rect 12912 27062 12940 30126
rect 13004 28762 13032 31146
rect 13188 31142 13216 31418
rect 13176 31136 13228 31142
rect 13176 31078 13228 31084
rect 13084 30660 13136 30666
rect 13084 30602 13136 30608
rect 13096 29714 13124 30602
rect 13280 29714 13308 32846
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13372 32434 13400 32710
rect 13360 32428 13412 32434
rect 13360 32370 13412 32376
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 13372 31634 13400 31826
rect 13556 31686 13584 34598
rect 13740 34066 13768 34614
rect 13728 34060 13780 34066
rect 13728 34002 13780 34008
rect 13636 33856 13688 33862
rect 13636 33798 13688 33804
rect 13452 31680 13504 31686
rect 13372 31628 13452 31634
rect 13372 31622 13504 31628
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 13372 31606 13492 31622
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 13372 30394 13400 30534
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 13084 29708 13136 29714
rect 13259 29708 13311 29714
rect 13136 29668 13216 29696
rect 13084 29650 13136 29656
rect 13084 29504 13136 29510
rect 13084 29446 13136 29452
rect 12992 28756 13044 28762
rect 12992 28698 13044 28704
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 13004 27946 13032 28494
rect 12992 27940 13044 27946
rect 12992 27882 13044 27888
rect 13004 27538 13032 27882
rect 12992 27532 13044 27538
rect 12992 27474 13044 27480
rect 12900 27056 12952 27062
rect 12900 26998 12952 27004
rect 12900 26444 12952 26450
rect 12900 26386 12952 26392
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 12912 25514 12940 26386
rect 13004 25838 13032 27474
rect 13096 26314 13124 29446
rect 13188 29102 13216 29668
rect 13259 29650 13311 29656
rect 13372 29646 13400 30330
rect 13464 30054 13492 31606
rect 13544 31136 13596 31142
rect 13544 31078 13596 31084
rect 13556 30666 13584 31078
rect 13544 30660 13596 30666
rect 13544 30602 13596 30608
rect 13452 30048 13504 30054
rect 13452 29990 13504 29996
rect 13452 29708 13504 29714
rect 13452 29650 13504 29656
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13176 29096 13228 29102
rect 13176 29038 13228 29044
rect 13176 28756 13228 28762
rect 13176 28698 13228 28704
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 12820 25486 12940 25514
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12820 24750 12848 25486
rect 12900 25424 12952 25430
rect 12900 25366 12952 25372
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12716 24336 12768 24342
rect 12716 24278 12768 24284
rect 12728 23866 12756 24278
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12728 22778 12756 23802
rect 12820 23730 12848 24686
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12912 22692 12940 25366
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 13004 24274 13032 24550
rect 12992 24268 13044 24274
rect 12992 24210 13044 24216
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13004 23186 13032 23258
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 12820 22664 12940 22692
rect 12820 22658 12848 22664
rect 12728 22630 12848 22658
rect 12728 20262 12756 22630
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12912 21146 12940 21422
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 13004 20992 13032 23122
rect 13096 21350 13124 25978
rect 13188 25430 13216 28698
rect 13280 28694 13308 29446
rect 13372 29170 13400 29582
rect 13464 29578 13492 29650
rect 13452 29572 13504 29578
rect 13452 29514 13504 29520
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13556 28994 13584 30602
rect 13372 28966 13584 28994
rect 13268 28688 13320 28694
rect 13268 28630 13320 28636
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13280 26926 13308 27270
rect 13268 26920 13320 26926
rect 13268 26862 13320 26868
rect 13280 26382 13308 26862
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13176 25424 13228 25430
rect 13176 25366 13228 25372
rect 13280 24342 13308 25638
rect 13268 24336 13320 24342
rect 13268 24278 13320 24284
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13188 23866 13216 24210
rect 13280 23866 13308 24278
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 13372 23798 13400 28966
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 13464 25362 13492 28018
rect 13648 26926 13676 33798
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13556 26450 13584 26862
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13636 26444 13688 26450
rect 13636 26386 13688 26392
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 13556 24750 13584 25774
rect 13648 25498 13676 26386
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13360 23792 13412 23798
rect 13360 23734 13412 23740
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 12912 20964 13032 20992
rect 13084 21004 13136 21010
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12912 19990 12940 20964
rect 13084 20946 13136 20952
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 13004 20398 13032 20810
rect 13096 20602 13124 20946
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13188 20482 13216 21626
rect 13280 21554 13308 23666
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13372 22438 13400 22714
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13372 22098 13400 22374
rect 13464 22098 13492 24686
rect 13556 23186 13584 24686
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13280 21010 13308 21286
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13372 20602 13400 21422
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13096 20454 13216 20482
rect 13360 20460 13412 20466
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12440 19508 12492 19514
rect 12544 19502 12848 19530
rect 12440 19450 12492 19456
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12360 18426 12388 18702
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12360 17746 12388 18362
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12452 17134 12480 19450
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12544 17338 12572 19314
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12636 17202 12664 19382
rect 12820 19334 12848 19502
rect 12912 19446 12940 19926
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 12728 19306 12848 19334
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12360 16794 12388 17070
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12072 14544 12124 14550
rect 12452 14498 12480 16730
rect 12728 16096 12756 19306
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18902 12940 19110
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12820 18086 12848 18294
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 13004 17882 13032 20334
rect 13096 19242 13124 20454
rect 13360 20402 13412 20408
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13084 19236 13136 19242
rect 13084 19178 13136 19184
rect 13096 18970 13124 19178
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16590 12848 17138
rect 13004 17134 13032 17818
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13096 17338 13124 17682
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12072 14486 12124 14492
rect 12176 14470 12480 14498
rect 12544 16068 12756 16096
rect 11992 12406 12112 12434
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11253 10364 11561 10384
rect 11253 10362 11259 10364
rect 11315 10362 11339 10364
rect 11395 10362 11419 10364
rect 11475 10362 11499 10364
rect 11555 10362 11561 10364
rect 11315 10310 11317 10362
rect 11497 10310 11499 10362
rect 11253 10308 11259 10310
rect 11315 10308 11339 10310
rect 11395 10308 11419 10310
rect 11475 10308 11499 10310
rect 11555 10308 11561 10310
rect 11253 10288 11561 10308
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8362 10732 8774
rect 10980 8498 11008 9318
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7342 10640 7686
rect 10704 7410 10732 8298
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7546 10824 7686
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10704 6934 10732 7346
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10612 5234 10640 6258
rect 10704 5778 10732 6870
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10796 5302 10824 7278
rect 10888 6866 10916 8366
rect 10980 7324 11008 8434
rect 11164 8430 11192 9862
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11253 9276 11561 9296
rect 11253 9274 11259 9276
rect 11315 9274 11339 9276
rect 11395 9274 11419 9276
rect 11475 9274 11499 9276
rect 11555 9274 11561 9276
rect 11315 9222 11317 9274
rect 11497 9222 11499 9274
rect 11253 9220 11259 9222
rect 11315 9220 11339 9222
rect 11395 9220 11419 9222
rect 11475 9220 11499 9222
rect 11555 9220 11561 9222
rect 11253 9200 11561 9220
rect 11624 9042 11652 9318
rect 11716 9178 11744 9862
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11072 8090 11100 8366
rect 11256 8276 11284 8910
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11164 8248 11284 8276
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11060 7336 11112 7342
rect 10980 7296 11060 7324
rect 11060 7278 11112 7284
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10704 4214 10732 5102
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3058 10640 3878
rect 10704 3602 10732 4150
rect 10888 3670 10916 6802
rect 11072 6798 11100 7278
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 5710 11100 6734
rect 11164 5896 11192 8248
rect 11253 8188 11561 8208
rect 11253 8186 11259 8188
rect 11315 8186 11339 8188
rect 11395 8186 11419 8188
rect 11475 8186 11499 8188
rect 11555 8186 11561 8188
rect 11315 8134 11317 8186
rect 11497 8134 11499 8186
rect 11253 8132 11259 8134
rect 11315 8132 11339 8134
rect 11395 8132 11419 8134
rect 11475 8132 11499 8134
rect 11555 8132 11561 8134
rect 11253 8112 11561 8132
rect 11624 7954 11652 8842
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11716 8090 11744 8230
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11808 7342 11836 9046
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11253 7100 11561 7120
rect 11253 7098 11259 7100
rect 11315 7098 11339 7100
rect 11395 7098 11419 7100
rect 11475 7098 11499 7100
rect 11555 7098 11561 7100
rect 11315 7046 11317 7098
rect 11497 7046 11499 7098
rect 11253 7044 11259 7046
rect 11315 7044 11339 7046
rect 11395 7044 11419 7046
rect 11475 7044 11499 7046
rect 11555 7044 11561 7046
rect 11253 7024 11561 7044
rect 11716 6866 11744 7142
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11253 6012 11561 6032
rect 11253 6010 11259 6012
rect 11315 6010 11339 6012
rect 11395 6010 11419 6012
rect 11475 6010 11499 6012
rect 11555 6010 11561 6012
rect 11315 5958 11317 6010
rect 11497 5958 11499 6010
rect 11253 5956 11259 5958
rect 11315 5956 11339 5958
rect 11395 5956 11419 5958
rect 11475 5956 11499 5958
rect 11555 5956 11561 5958
rect 11253 5936 11561 5956
rect 11164 5868 11284 5896
rect 11256 5778 11284 5868
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10980 5234 11008 5510
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10980 4078 11008 5034
rect 11072 4690 11100 5238
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10612 1494 10640 2790
rect 10704 2582 10732 3538
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10796 2514 10824 2926
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10704 2310 10732 2382
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 10888 1902 10916 3606
rect 10980 2854 11008 4014
rect 11072 3738 11100 4626
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11164 3194 11192 5714
rect 11256 5302 11284 5714
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11624 5098 11652 6394
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11253 4924 11561 4944
rect 11253 4922 11259 4924
rect 11315 4922 11339 4924
rect 11395 4922 11419 4924
rect 11475 4922 11499 4924
rect 11555 4922 11561 4924
rect 11315 4870 11317 4922
rect 11497 4870 11499 4922
rect 11253 4868 11259 4870
rect 11315 4868 11339 4870
rect 11395 4868 11419 4870
rect 11475 4868 11499 4870
rect 11555 4868 11561 4870
rect 11253 4848 11561 4868
rect 11253 3836 11561 3856
rect 11253 3834 11259 3836
rect 11315 3834 11339 3836
rect 11395 3834 11419 3836
rect 11475 3834 11499 3836
rect 11555 3834 11561 3836
rect 11315 3782 11317 3834
rect 11497 3782 11499 3834
rect 11253 3780 11259 3782
rect 11315 3780 11339 3782
rect 11395 3780 11419 3782
rect 11475 3780 11499 3782
rect 11555 3780 11561 3782
rect 11253 3760 11561 3780
rect 11808 3398 11836 6802
rect 11900 6458 11928 10134
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 5370 12020 11630
rect 12084 11218 12112 12406
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12084 5914 12112 8434
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4690 11928 4966
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11253 2748 11561 2768
rect 11253 2746 11259 2748
rect 11315 2746 11339 2748
rect 11395 2746 11419 2748
rect 11475 2746 11499 2748
rect 11555 2746 11561 2748
rect 11315 2694 11317 2746
rect 11497 2694 11499 2746
rect 11253 2692 11259 2694
rect 11315 2692 11339 2694
rect 11395 2692 11419 2694
rect 11475 2692 11499 2694
rect 11555 2692 11561 2694
rect 11253 2672 11561 2692
rect 11992 2514 12020 2858
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 10876 1896 10928 1902
rect 10876 1838 10928 1844
rect 10600 1488 10652 1494
rect 10600 1430 10652 1436
rect 10888 1426 10916 1838
rect 11253 1660 11561 1680
rect 11253 1658 11259 1660
rect 11315 1658 11339 1660
rect 11395 1658 11419 1660
rect 11475 1658 11499 1660
rect 11555 1658 11561 1660
rect 11315 1606 11317 1658
rect 11497 1606 11499 1658
rect 11253 1604 11259 1606
rect 11315 1604 11339 1606
rect 11395 1604 11419 1606
rect 11475 1604 11499 1606
rect 11555 1604 11561 1606
rect 11253 1584 11561 1604
rect 10876 1420 10928 1426
rect 10876 1362 10928 1368
rect 10520 1312 10640 1340
rect 10612 1222 10640 1312
rect 10600 1216 10652 1222
rect 10600 1158 10652 1164
rect 8392 1012 8444 1018
rect 8392 954 8444 960
rect 11716 950 11744 2450
rect 12084 2106 12112 3538
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 12176 1290 12204 14470
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12268 12102 12296 14214
rect 12544 12918 12572 16068
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12636 15722 12664 15914
rect 12636 15694 12756 15722
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12360 12442 12388 12718
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12268 11354 12296 11562
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12452 9654 12480 12310
rect 12636 11354 12664 14554
rect 12728 13734 12756 15694
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12820 13682 12848 16390
rect 12912 15910 12940 16594
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12912 13938 12940 15098
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13004 13870 13032 17070
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13096 16250 13124 16526
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 12820 13654 13032 13682
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 12850 12940 13194
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12728 12306 12756 12650
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12912 12102 12940 12786
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 8430 12296 8774
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12268 7342 12296 7958
rect 12360 7954 12388 8978
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12452 6866 12480 8910
rect 12544 7954 12572 10542
rect 12636 10198 12664 11290
rect 13004 10554 13032 13654
rect 13096 13394 13124 16186
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12808 10532 12860 10538
rect 13004 10526 13124 10554
rect 12808 10474 12860 10480
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 9160 12664 9862
rect 12728 9586 12756 10066
rect 12820 9926 12848 10474
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 13004 9586 13032 10406
rect 13096 10130 13124 10526
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13188 9654 13216 19790
rect 13280 18850 13308 20198
rect 13372 19922 13400 20402
rect 13464 20058 13492 20946
rect 13556 20942 13584 22714
rect 13648 21690 13676 25298
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13372 19514 13400 19858
rect 13556 19530 13584 20742
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13464 19502 13584 19530
rect 13372 18970 13400 19450
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13280 18822 13400 18850
rect 13464 18834 13492 19502
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13280 16454 13308 18294
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13372 16266 13400 18822
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13556 17678 13584 19382
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13556 16794 13584 17614
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13280 16238 13400 16266
rect 13280 15978 13308 16238
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13280 13802 13308 15574
rect 13372 15570 13400 15846
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13464 15162 13492 16594
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13556 14958 13584 15302
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13372 14074 13400 14418
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13280 12442 13308 12650
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13372 11898 13400 12310
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13464 10826 13492 13670
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13280 10798 13492 10826
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12636 9132 12756 9160
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12636 8634 12664 8978
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12728 7750 12756 9132
rect 12912 8634 12940 9454
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13096 8566 13124 8910
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13188 8430 13216 9590
rect 13176 8424 13228 8430
rect 13096 8384 13176 8412
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 13096 7546 13124 8384
rect 13176 8366 13228 8372
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13096 7342 13124 7482
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12268 6458 12296 6802
rect 12544 6662 12572 7278
rect 13188 7206 13216 7822
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13280 6984 13308 10798
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13004 6956 13308 6984
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12360 5710 12388 6258
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12360 5234 12388 5646
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12268 4554 12296 5034
rect 12360 4554 12388 5170
rect 12544 4758 12572 6598
rect 12728 6254 12756 6870
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12636 5166 12664 6122
rect 12728 5302 12756 6190
rect 12820 5574 12848 6190
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12728 4570 12756 5238
rect 12820 5166 12848 5510
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12820 4690 12848 5102
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12268 4078 12296 4490
rect 12360 4282 12388 4490
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12452 4078 12480 4558
rect 12728 4542 12848 4570
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12624 4208 12676 4214
rect 12544 4168 12624 4196
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12452 3194 12480 4014
rect 12544 4010 12572 4168
rect 12624 4150 12676 4156
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12728 2990 12756 4422
rect 12820 4282 12848 4542
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12728 2650 12756 2790
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 1834 12296 2246
rect 12256 1828 12308 1834
rect 12256 1770 12308 1776
rect 12164 1284 12216 1290
rect 12164 1226 12216 1232
rect 8300 944 8352 950
rect 8300 886 8352 892
rect 11704 944 11756 950
rect 11704 886 11756 892
rect 8312 800 8340 886
rect 12912 814 12940 3878
rect 13004 2106 13032 6956
rect 13372 6848 13400 10474
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8634 13492 9046
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13464 8022 13492 8570
rect 13556 8430 13584 13330
rect 13648 9042 13676 21354
rect 13740 10810 13768 34002
rect 13820 33380 13872 33386
rect 13820 33322 13872 33328
rect 13832 33114 13860 33322
rect 13820 33108 13872 33114
rect 13820 33050 13872 33056
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 13832 31958 13860 32914
rect 13820 31952 13872 31958
rect 13820 31894 13872 31900
rect 13924 31754 13952 44202
rect 14200 41750 14228 45494
rect 14292 44402 14320 45494
rect 14280 44396 14332 44402
rect 14280 44338 14332 44344
rect 14384 43246 14412 46446
rect 14648 46436 14700 46442
rect 14648 46378 14700 46384
rect 14660 46170 14688 46378
rect 15108 46368 15160 46374
rect 15108 46310 15160 46316
rect 14648 46164 14700 46170
rect 14648 46106 14700 46112
rect 15120 46034 15148 46310
rect 15396 46102 15424 47194
rect 15764 46170 15792 47466
rect 15856 47258 15884 48146
rect 15936 48000 15988 48006
rect 15936 47942 15988 47948
rect 16764 48000 16816 48006
rect 16764 47942 16816 47948
rect 20076 48000 20128 48006
rect 20076 47942 20128 47948
rect 15844 47252 15896 47258
rect 15844 47194 15896 47200
rect 15752 46164 15804 46170
rect 15752 46106 15804 46112
rect 15384 46096 15436 46102
rect 15384 46038 15436 46044
rect 14832 46028 14884 46034
rect 14832 45970 14884 45976
rect 15108 46028 15160 46034
rect 15108 45970 15160 45976
rect 14844 45422 14872 45970
rect 15292 45960 15344 45966
rect 15292 45902 15344 45908
rect 15304 45626 15332 45902
rect 15292 45620 15344 45626
rect 15292 45562 15344 45568
rect 15752 45484 15804 45490
rect 15752 45426 15804 45432
rect 14648 45416 14700 45422
rect 14648 45358 14700 45364
rect 14832 45416 14884 45422
rect 14832 45358 14884 45364
rect 14660 45098 14688 45358
rect 14568 45070 14688 45098
rect 14844 45082 14872 45358
rect 15108 45280 15160 45286
rect 15108 45222 15160 45228
rect 15568 45280 15620 45286
rect 15568 45222 15620 45228
rect 14832 45076 14884 45082
rect 14464 44396 14516 44402
rect 14464 44338 14516 44344
rect 14476 43790 14504 44338
rect 14568 43926 14596 45070
rect 14832 45018 14884 45024
rect 15120 45014 15148 45222
rect 15108 45008 15160 45014
rect 15108 44950 15160 44956
rect 14648 44940 14700 44946
rect 14648 44882 14700 44888
rect 15476 44940 15528 44946
rect 15476 44882 15528 44888
rect 14660 43994 14688 44882
rect 15488 44334 15516 44882
rect 15476 44328 15528 44334
rect 15476 44270 15528 44276
rect 14648 43988 14700 43994
rect 14648 43930 14700 43936
rect 14556 43920 14608 43926
rect 14556 43862 14608 43868
rect 15580 43858 15608 45222
rect 15764 45082 15792 45426
rect 15752 45076 15804 45082
rect 15752 45018 15804 45024
rect 15764 44946 15792 45018
rect 15948 44946 15976 47942
rect 16405 47900 16713 47920
rect 16405 47898 16411 47900
rect 16467 47898 16491 47900
rect 16547 47898 16571 47900
rect 16627 47898 16651 47900
rect 16707 47898 16713 47900
rect 16467 47846 16469 47898
rect 16649 47846 16651 47898
rect 16405 47844 16411 47846
rect 16467 47844 16491 47846
rect 16547 47844 16571 47846
rect 16627 47844 16651 47846
rect 16707 47844 16713 47846
rect 16405 47824 16713 47844
rect 16120 47456 16172 47462
rect 16120 47398 16172 47404
rect 16132 47122 16160 47398
rect 16120 47116 16172 47122
rect 16120 47058 16172 47064
rect 16028 46980 16080 46986
rect 16028 46922 16080 46928
rect 15752 44940 15804 44946
rect 15672 44900 15752 44928
rect 14924 43852 14976 43858
rect 14924 43794 14976 43800
rect 15568 43852 15620 43858
rect 15568 43794 15620 43800
rect 14464 43784 14516 43790
rect 14464 43726 14516 43732
rect 14464 43648 14516 43654
rect 14464 43590 14516 43596
rect 14476 43314 14504 43590
rect 14464 43308 14516 43314
rect 14464 43250 14516 43256
rect 14372 43240 14424 43246
rect 14372 43182 14424 43188
rect 14476 42702 14504 43250
rect 14936 42838 14964 43794
rect 15200 43784 15252 43790
rect 15200 43726 15252 43732
rect 15108 43104 15160 43110
rect 15212 43058 15240 43726
rect 15292 43648 15344 43654
rect 15292 43590 15344 43596
rect 15160 43052 15240 43058
rect 15108 43046 15240 43052
rect 15120 43030 15240 43046
rect 14924 42832 14976 42838
rect 14924 42774 14976 42780
rect 15212 42770 15240 43030
rect 14832 42764 14884 42770
rect 14832 42706 14884 42712
rect 15200 42764 15252 42770
rect 15200 42706 15252 42712
rect 14464 42696 14516 42702
rect 14464 42638 14516 42644
rect 14476 42140 14504 42638
rect 14556 42152 14608 42158
rect 14476 42112 14556 42140
rect 14556 42094 14608 42100
rect 14648 42152 14700 42158
rect 14648 42094 14700 42100
rect 14188 41744 14240 41750
rect 14188 41686 14240 41692
rect 14004 39976 14056 39982
rect 14004 39918 14056 39924
rect 14016 39846 14044 39918
rect 14004 39840 14056 39846
rect 14004 39782 14056 39788
rect 14016 37670 14044 39782
rect 14004 37664 14056 37670
rect 14004 37606 14056 37612
rect 13832 31726 13952 31754
rect 13832 30870 13860 31726
rect 13912 31680 13964 31686
rect 13912 31622 13964 31628
rect 13820 30864 13872 30870
rect 13820 30806 13872 30812
rect 13820 30728 13872 30734
rect 13820 30670 13872 30676
rect 13832 29646 13860 30670
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 13924 27946 13952 31622
rect 13912 27940 13964 27946
rect 13912 27882 13964 27888
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13832 24274 13860 26182
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13924 24954 13952 25230
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13832 23730 13860 24210
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13832 23186 13860 23462
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13832 14822 13860 19654
rect 13924 16726 13952 23802
rect 14016 18426 14044 37606
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 14108 36786 14136 37062
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 14108 36582 14136 36722
rect 14096 36576 14148 36582
rect 14096 36518 14148 36524
rect 14108 36038 14136 36518
rect 14096 36032 14148 36038
rect 14096 35974 14148 35980
rect 14096 35488 14148 35494
rect 14096 35430 14148 35436
rect 14108 34202 14136 35430
rect 14200 34474 14228 41686
rect 14280 41200 14332 41206
rect 14280 41142 14332 41148
rect 14292 39982 14320 41142
rect 14372 40996 14424 41002
rect 14372 40938 14424 40944
rect 14384 40050 14412 40938
rect 14568 40390 14596 42094
rect 14556 40384 14608 40390
rect 14556 40326 14608 40332
rect 14568 40118 14596 40326
rect 14556 40112 14608 40118
rect 14556 40054 14608 40060
rect 14372 40044 14424 40050
rect 14372 39986 14424 39992
rect 14280 39976 14332 39982
rect 14280 39918 14332 39924
rect 14660 38554 14688 42094
rect 14740 42084 14792 42090
rect 14740 42026 14792 42032
rect 14752 40934 14780 42026
rect 14844 41274 14872 42706
rect 15016 42696 15068 42702
rect 15016 42638 15068 42644
rect 15028 42226 15056 42638
rect 15016 42220 15068 42226
rect 15016 42162 15068 42168
rect 15200 41608 15252 41614
rect 15200 41550 15252 41556
rect 14832 41268 14884 41274
rect 14832 41210 14884 41216
rect 14740 40928 14792 40934
rect 14740 40870 14792 40876
rect 14752 40730 14780 40870
rect 14740 40724 14792 40730
rect 14740 40666 14792 40672
rect 14752 39982 14780 40666
rect 14740 39976 14792 39982
rect 14740 39918 14792 39924
rect 15212 39642 15240 41550
rect 15200 39636 15252 39642
rect 15200 39578 15252 39584
rect 15108 39500 15160 39506
rect 15108 39442 15160 39448
rect 14832 39364 14884 39370
rect 14832 39306 14884 39312
rect 14648 38548 14700 38554
rect 14648 38490 14700 38496
rect 14556 37800 14608 37806
rect 14556 37742 14608 37748
rect 14372 35624 14424 35630
rect 14372 35566 14424 35572
rect 14384 35494 14412 35566
rect 14372 35488 14424 35494
rect 14372 35430 14424 35436
rect 14384 34746 14412 35430
rect 14464 35148 14516 35154
rect 14464 35090 14516 35096
rect 14372 34740 14424 34746
rect 14372 34682 14424 34688
rect 14188 34468 14240 34474
rect 14188 34410 14240 34416
rect 14096 34196 14148 34202
rect 14096 34138 14148 34144
rect 14096 33448 14148 33454
rect 14096 33390 14148 33396
rect 14108 32570 14136 33390
rect 14384 32978 14412 34682
rect 14476 34542 14504 35090
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14372 32972 14424 32978
rect 14372 32914 14424 32920
rect 14476 32842 14504 34478
rect 14464 32836 14516 32842
rect 14464 32778 14516 32784
rect 14568 32570 14596 37742
rect 14740 36644 14792 36650
rect 14740 36586 14792 36592
rect 14752 35290 14780 36586
rect 14740 35284 14792 35290
rect 14740 35226 14792 35232
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14660 34950 14688 35022
rect 14648 34944 14700 34950
rect 14648 34886 14700 34892
rect 14660 34610 14688 34886
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14740 34400 14792 34406
rect 14740 34342 14792 34348
rect 14752 33930 14780 34342
rect 14844 34134 14872 39306
rect 15120 37806 15148 39442
rect 15200 39296 15252 39302
rect 15200 39238 15252 39244
rect 15212 38894 15240 39238
rect 15304 39030 15332 43590
rect 15672 43450 15700 44900
rect 15752 44882 15804 44888
rect 15936 44940 15988 44946
rect 15936 44882 15988 44888
rect 15844 44872 15896 44878
rect 15844 44814 15896 44820
rect 15752 44328 15804 44334
rect 15752 44270 15804 44276
rect 15764 43926 15792 44270
rect 15752 43920 15804 43926
rect 15752 43862 15804 43868
rect 15660 43444 15712 43450
rect 15660 43386 15712 43392
rect 15476 43240 15528 43246
rect 15476 43182 15528 43188
rect 15568 43240 15620 43246
rect 15568 43182 15620 43188
rect 15384 43172 15436 43178
rect 15384 43114 15436 43120
rect 15396 42906 15424 43114
rect 15384 42900 15436 42906
rect 15384 42842 15436 42848
rect 15384 42016 15436 42022
rect 15384 41958 15436 41964
rect 15396 39370 15424 41958
rect 15488 41478 15516 43182
rect 15580 42634 15608 43182
rect 15568 42628 15620 42634
rect 15568 42570 15620 42576
rect 15764 41750 15792 43862
rect 15856 42634 15884 44814
rect 15936 44736 15988 44742
rect 15936 44678 15988 44684
rect 15948 44180 15976 44678
rect 16040 44334 16068 46922
rect 16132 46102 16160 47058
rect 16405 46812 16713 46832
rect 16405 46810 16411 46812
rect 16467 46810 16491 46812
rect 16547 46810 16571 46812
rect 16627 46810 16651 46812
rect 16707 46810 16713 46812
rect 16467 46758 16469 46810
rect 16649 46758 16651 46810
rect 16405 46756 16411 46758
rect 16467 46756 16491 46758
rect 16547 46756 16571 46758
rect 16627 46756 16651 46758
rect 16707 46756 16713 46758
rect 16405 46736 16713 46756
rect 16672 46504 16724 46510
rect 16672 46446 16724 46452
rect 16304 46368 16356 46374
rect 16304 46310 16356 46316
rect 16120 46096 16172 46102
rect 16120 46038 16172 46044
rect 16212 45552 16264 45558
rect 16212 45494 16264 45500
rect 16120 44804 16172 44810
rect 16120 44746 16172 44752
rect 16028 44328 16080 44334
rect 16028 44270 16080 44276
rect 15948 44152 16068 44180
rect 15936 43716 15988 43722
rect 15936 43658 15988 43664
rect 15844 42628 15896 42634
rect 15844 42570 15896 42576
rect 15844 42016 15896 42022
rect 15844 41958 15896 41964
rect 15752 41744 15804 41750
rect 15752 41686 15804 41692
rect 15476 41472 15528 41478
rect 15476 41414 15528 41420
rect 15752 41472 15804 41478
rect 15752 41414 15804 41420
rect 15488 41070 15516 41414
rect 15476 41064 15528 41070
rect 15476 41006 15528 41012
rect 15568 39432 15620 39438
rect 15568 39374 15620 39380
rect 15384 39364 15436 39370
rect 15384 39306 15436 39312
rect 15292 39024 15344 39030
rect 15292 38966 15344 38972
rect 15580 38962 15608 39374
rect 15660 39296 15712 39302
rect 15660 39238 15712 39244
rect 15672 39098 15700 39238
rect 15660 39092 15712 39098
rect 15660 39034 15712 39040
rect 15568 38956 15620 38962
rect 15568 38898 15620 38904
rect 15200 38888 15252 38894
rect 15200 38830 15252 38836
rect 15384 38888 15436 38894
rect 15384 38830 15436 38836
rect 15476 38888 15528 38894
rect 15476 38830 15528 38836
rect 15292 38820 15344 38826
rect 15292 38762 15344 38768
rect 15304 38010 15332 38762
rect 15292 38004 15344 38010
rect 15292 37946 15344 37952
rect 15108 37800 15160 37806
rect 15108 37742 15160 37748
rect 15396 37738 15424 38830
rect 15488 37942 15516 38830
rect 15476 37936 15528 37942
rect 15476 37878 15528 37884
rect 15384 37732 15436 37738
rect 15384 37674 15436 37680
rect 15488 37398 15516 37878
rect 15476 37392 15528 37398
rect 15476 37334 15528 37340
rect 15672 37330 15700 39034
rect 15764 37874 15792 41414
rect 15752 37868 15804 37874
rect 15752 37810 15804 37816
rect 15856 37806 15884 41958
rect 15948 39506 15976 43658
rect 16040 40390 16068 44152
rect 16132 43858 16160 44746
rect 16224 44742 16252 45494
rect 16212 44736 16264 44742
rect 16212 44678 16264 44684
rect 16212 44396 16264 44402
rect 16212 44338 16264 44344
rect 16120 43852 16172 43858
rect 16120 43794 16172 43800
rect 16224 43790 16252 44338
rect 16316 43926 16344 46310
rect 16684 46034 16712 46446
rect 16672 46028 16724 46034
rect 16672 45970 16724 45976
rect 16405 45724 16713 45744
rect 16405 45722 16411 45724
rect 16467 45722 16491 45724
rect 16547 45722 16571 45724
rect 16627 45722 16651 45724
rect 16707 45722 16713 45724
rect 16467 45670 16469 45722
rect 16649 45670 16651 45722
rect 16405 45668 16411 45670
rect 16467 45668 16491 45670
rect 16547 45668 16571 45670
rect 16627 45668 16651 45670
rect 16707 45668 16713 45670
rect 16405 45648 16713 45668
rect 16672 45348 16724 45354
rect 16672 45290 16724 45296
rect 16684 44810 16712 45290
rect 16672 44804 16724 44810
rect 16672 44746 16724 44752
rect 16405 44636 16713 44656
rect 16405 44634 16411 44636
rect 16467 44634 16491 44636
rect 16547 44634 16571 44636
rect 16627 44634 16651 44636
rect 16707 44634 16713 44636
rect 16467 44582 16469 44634
rect 16649 44582 16651 44634
rect 16405 44580 16411 44582
rect 16467 44580 16491 44582
rect 16547 44580 16571 44582
rect 16627 44580 16651 44582
rect 16707 44580 16713 44582
rect 16405 44560 16713 44580
rect 16396 44192 16448 44198
rect 16396 44134 16448 44140
rect 16304 43920 16356 43926
rect 16304 43862 16356 43868
rect 16212 43784 16264 43790
rect 16212 43726 16264 43732
rect 16120 42560 16172 42566
rect 16120 42502 16172 42508
rect 16132 42226 16160 42502
rect 16120 42220 16172 42226
rect 16120 42162 16172 42168
rect 16224 42158 16252 43726
rect 16408 43722 16436 44134
rect 16396 43716 16448 43722
rect 16396 43658 16448 43664
rect 16405 43548 16713 43568
rect 16405 43546 16411 43548
rect 16467 43546 16491 43548
rect 16547 43546 16571 43548
rect 16627 43546 16651 43548
rect 16707 43546 16713 43548
rect 16467 43494 16469 43546
rect 16649 43494 16651 43546
rect 16405 43492 16411 43494
rect 16467 43492 16491 43494
rect 16547 43492 16571 43494
rect 16627 43492 16651 43494
rect 16707 43492 16713 43494
rect 16405 43472 16713 43492
rect 16405 42460 16713 42480
rect 16405 42458 16411 42460
rect 16467 42458 16491 42460
rect 16547 42458 16571 42460
rect 16627 42458 16651 42460
rect 16707 42458 16713 42460
rect 16467 42406 16469 42458
rect 16649 42406 16651 42458
rect 16405 42404 16411 42406
rect 16467 42404 16491 42406
rect 16547 42404 16571 42406
rect 16627 42404 16651 42406
rect 16707 42404 16713 42406
rect 16405 42384 16713 42404
rect 16396 42288 16448 42294
rect 16316 42236 16396 42242
rect 16316 42230 16448 42236
rect 16316 42214 16436 42230
rect 16212 42152 16264 42158
rect 16212 42094 16264 42100
rect 16224 42022 16252 42094
rect 16212 42016 16264 42022
rect 16212 41958 16264 41964
rect 16316 41750 16344 42214
rect 16304 41744 16356 41750
rect 16304 41686 16356 41692
rect 16212 41676 16264 41682
rect 16212 41618 16264 41624
rect 16120 41132 16172 41138
rect 16120 41074 16172 41080
rect 16132 40662 16160 41074
rect 16224 40934 16252 41618
rect 16212 40928 16264 40934
rect 16212 40870 16264 40876
rect 16120 40656 16172 40662
rect 16120 40598 16172 40604
rect 16028 40384 16080 40390
rect 16028 40326 16080 40332
rect 16212 40384 16264 40390
rect 16212 40326 16264 40332
rect 15936 39500 15988 39506
rect 15936 39442 15988 39448
rect 16224 38826 16252 40326
rect 16316 40186 16344 41686
rect 16405 41372 16713 41392
rect 16405 41370 16411 41372
rect 16467 41370 16491 41372
rect 16547 41370 16571 41372
rect 16627 41370 16651 41372
rect 16707 41370 16713 41372
rect 16467 41318 16469 41370
rect 16649 41318 16651 41370
rect 16405 41316 16411 41318
rect 16467 41316 16491 41318
rect 16547 41316 16571 41318
rect 16627 41316 16651 41318
rect 16707 41316 16713 41318
rect 16405 41296 16713 41316
rect 16405 40284 16713 40304
rect 16405 40282 16411 40284
rect 16467 40282 16491 40284
rect 16547 40282 16571 40284
rect 16627 40282 16651 40284
rect 16707 40282 16713 40284
rect 16467 40230 16469 40282
rect 16649 40230 16651 40282
rect 16405 40228 16411 40230
rect 16467 40228 16491 40230
rect 16547 40228 16571 40230
rect 16627 40228 16651 40230
rect 16707 40228 16713 40230
rect 16405 40208 16713 40228
rect 16304 40180 16356 40186
rect 16304 40122 16356 40128
rect 16405 39196 16713 39216
rect 16405 39194 16411 39196
rect 16467 39194 16491 39196
rect 16547 39194 16571 39196
rect 16627 39194 16651 39196
rect 16707 39194 16713 39196
rect 16467 39142 16469 39194
rect 16649 39142 16651 39194
rect 16405 39140 16411 39142
rect 16467 39140 16491 39142
rect 16547 39140 16571 39142
rect 16627 39140 16651 39142
rect 16707 39140 16713 39142
rect 16405 39120 16713 39140
rect 16212 38820 16264 38826
rect 16212 38762 16264 38768
rect 16672 38412 16724 38418
rect 16672 38354 16724 38360
rect 16684 38282 16712 38354
rect 16672 38276 16724 38282
rect 16672 38218 16724 38224
rect 16304 38208 16356 38214
rect 16304 38150 16356 38156
rect 15844 37800 15896 37806
rect 15844 37742 15896 37748
rect 15936 37800 15988 37806
rect 15936 37742 15988 37748
rect 15844 37664 15896 37670
rect 15844 37606 15896 37612
rect 15856 37346 15884 37606
rect 15948 37466 15976 37742
rect 16316 37466 16344 38150
rect 16405 38108 16713 38128
rect 16405 38106 16411 38108
rect 16467 38106 16491 38108
rect 16547 38106 16571 38108
rect 16627 38106 16651 38108
rect 16707 38106 16713 38108
rect 16467 38054 16469 38106
rect 16649 38054 16651 38106
rect 16405 38052 16411 38054
rect 16467 38052 16491 38054
rect 16547 38052 16571 38054
rect 16627 38052 16651 38054
rect 16707 38052 16713 38054
rect 16405 38032 16713 38052
rect 15936 37460 15988 37466
rect 15936 37402 15988 37408
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 15660 37324 15712 37330
rect 15856 37318 15976 37346
rect 15660 37266 15712 37272
rect 15568 36576 15620 36582
rect 15568 36518 15620 36524
rect 15016 36236 15068 36242
rect 15016 36178 15068 36184
rect 14924 35556 14976 35562
rect 14924 35498 14976 35504
rect 14936 35154 14964 35498
rect 14924 35148 14976 35154
rect 14924 35090 14976 35096
rect 15028 34746 15056 36178
rect 15476 36168 15528 36174
rect 15476 36110 15528 36116
rect 15108 35624 15160 35630
rect 15108 35566 15160 35572
rect 15016 34740 15068 34746
rect 15016 34682 15068 34688
rect 15016 34400 15068 34406
rect 15016 34342 15068 34348
rect 14832 34128 14884 34134
rect 14832 34070 14884 34076
rect 14844 33998 14872 34070
rect 14832 33992 14884 33998
rect 14832 33934 14884 33940
rect 14740 33924 14792 33930
rect 14740 33866 14792 33872
rect 14096 32564 14148 32570
rect 14096 32506 14148 32512
rect 14556 32564 14608 32570
rect 14556 32506 14608 32512
rect 14108 30802 14136 32506
rect 14280 32360 14332 32366
rect 14280 32302 14332 32308
rect 14292 32026 14320 32302
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14280 31272 14332 31278
rect 14280 31214 14332 31220
rect 14096 30796 14148 30802
rect 14096 30738 14148 30744
rect 14292 30734 14320 31214
rect 14752 31210 14780 33866
rect 14844 32366 14872 33934
rect 14924 33856 14976 33862
rect 14924 33798 14976 33804
rect 14936 33318 14964 33798
rect 14924 33312 14976 33318
rect 14924 33254 14976 33260
rect 15028 32978 15056 34342
rect 15120 33998 15148 35566
rect 15384 35556 15436 35562
rect 15384 35498 15436 35504
rect 15292 35284 15344 35290
rect 15292 35226 15344 35232
rect 15304 35018 15332 35226
rect 15292 35012 15344 35018
rect 15292 34954 15344 34960
rect 15396 34746 15424 35498
rect 15488 35290 15516 36110
rect 15476 35284 15528 35290
rect 15476 35226 15528 35232
rect 15476 35080 15528 35086
rect 15476 35022 15528 35028
rect 15488 34762 15516 35022
rect 15580 34950 15608 36518
rect 15568 34944 15620 34950
rect 15568 34886 15620 34892
rect 15384 34740 15436 34746
rect 15488 34734 15608 34762
rect 15384 34682 15436 34688
rect 15476 34672 15528 34678
rect 15476 34614 15528 34620
rect 15384 34604 15436 34610
rect 15384 34546 15436 34552
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15292 33992 15344 33998
rect 15292 33934 15344 33940
rect 15120 33522 15148 33934
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 15200 33312 15252 33318
rect 15200 33254 15252 33260
rect 15016 32972 15068 32978
rect 15016 32914 15068 32920
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 15120 32570 15148 32914
rect 15212 32842 15240 33254
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 14924 32564 14976 32570
rect 14924 32506 14976 32512
rect 15108 32564 15160 32570
rect 15108 32506 15160 32512
rect 14832 32360 14884 32366
rect 14832 32302 14884 32308
rect 14936 31890 14964 32506
rect 15304 32298 15332 33934
rect 15396 32978 15424 34546
rect 15488 32978 15516 34614
rect 15580 34542 15608 34734
rect 15568 34536 15620 34542
rect 15568 34478 15620 34484
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 15384 32972 15436 32978
rect 15384 32914 15436 32920
rect 15476 32972 15528 32978
rect 15476 32914 15528 32920
rect 15292 32292 15344 32298
rect 15292 32234 15344 32240
rect 14924 31884 14976 31890
rect 14924 31826 14976 31832
rect 15108 31816 15160 31822
rect 15108 31758 15160 31764
rect 15016 31680 15068 31686
rect 15016 31622 15068 31628
rect 14740 31204 14792 31210
rect 14740 31146 14792 31152
rect 14372 31136 14424 31142
rect 14372 31078 14424 31084
rect 14384 30938 14412 31078
rect 14372 30932 14424 30938
rect 14372 30874 14424 30880
rect 15028 30870 15056 31622
rect 15120 31278 15148 31758
rect 15108 31272 15160 31278
rect 15108 31214 15160 31220
rect 14464 30864 14516 30870
rect 14464 30806 14516 30812
rect 15016 30864 15068 30870
rect 15016 30806 15068 30812
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14476 29832 14504 30806
rect 14740 30796 14792 30802
rect 14740 30738 14792 30744
rect 14752 30190 14780 30738
rect 14740 30184 14792 30190
rect 14740 30126 14792 30132
rect 15016 30116 15068 30122
rect 15016 30058 15068 30064
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14384 29804 14504 29832
rect 14556 29844 14608 29850
rect 14280 29776 14332 29782
rect 14280 29718 14332 29724
rect 14292 29102 14320 29718
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 14096 29028 14148 29034
rect 14096 28970 14148 28976
rect 14108 28014 14136 28970
rect 14280 28756 14332 28762
rect 14280 28698 14332 28704
rect 14292 28014 14320 28698
rect 14096 28008 14148 28014
rect 14096 27950 14148 27956
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14108 27538 14136 27950
rect 14188 27940 14240 27946
rect 14188 27882 14240 27888
rect 14096 27532 14148 27538
rect 14096 27474 14148 27480
rect 14200 25362 14228 27882
rect 14292 27334 14320 27950
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14292 26042 14320 26862
rect 14384 26194 14412 29804
rect 14556 29786 14608 29792
rect 14464 29708 14516 29714
rect 14464 29650 14516 29656
rect 14476 29102 14504 29650
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 14476 28762 14504 29038
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14568 27520 14596 29786
rect 14844 29102 14872 29990
rect 15028 29102 15056 30058
rect 15120 29170 15148 31214
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15212 29510 15240 29582
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 14832 29096 14884 29102
rect 14832 29038 14884 29044
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 15016 28620 15068 28626
rect 15016 28562 15068 28568
rect 14832 28552 14884 28558
rect 14832 28494 14884 28500
rect 14648 28416 14700 28422
rect 14648 28358 14700 28364
rect 14660 28014 14688 28358
rect 14844 28218 14872 28494
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 14648 28008 14700 28014
rect 14648 27950 14700 27956
rect 14740 27872 14792 27878
rect 14740 27814 14792 27820
rect 14648 27532 14700 27538
rect 14568 27492 14648 27520
rect 14648 27474 14700 27480
rect 14660 26858 14688 27474
rect 14464 26852 14516 26858
rect 14464 26794 14516 26800
rect 14648 26852 14700 26858
rect 14648 26794 14700 26800
rect 14476 26382 14504 26794
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 14384 26166 14504 26194
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14372 26036 14424 26042
rect 14372 25978 14424 25984
rect 14384 25362 14412 25978
rect 14476 25702 14504 26166
rect 14648 25832 14700 25838
rect 14648 25774 14700 25780
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14188 25356 14240 25362
rect 14188 25298 14240 25304
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14108 24886 14136 25230
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 14200 24732 14228 25162
rect 14108 24704 14228 24732
rect 14108 18970 14136 24704
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 14200 22982 14228 24210
rect 14384 23662 14412 25298
rect 14476 25294 14504 25638
rect 14660 25294 14688 25774
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14752 24750 14780 27814
rect 15028 27674 15056 28562
rect 15016 27668 15068 27674
rect 15016 27610 15068 27616
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14936 25974 14964 26930
rect 15016 26852 15068 26858
rect 15016 26794 15068 26800
rect 14924 25968 14976 25974
rect 14924 25910 14976 25916
rect 15028 25770 15056 26794
rect 15016 25764 15068 25770
rect 15016 25706 15068 25712
rect 15212 24954 15240 29446
rect 15304 28994 15332 32234
rect 15396 31890 15424 32914
rect 15488 32502 15516 32914
rect 15672 32910 15700 34478
rect 15844 34400 15896 34406
rect 15844 34342 15896 34348
rect 15752 33380 15804 33386
rect 15752 33322 15804 33328
rect 15764 33114 15792 33322
rect 15752 33108 15804 33114
rect 15752 33050 15804 33056
rect 15752 32972 15804 32978
rect 15752 32914 15804 32920
rect 15660 32904 15712 32910
rect 15660 32846 15712 32852
rect 15476 32496 15528 32502
rect 15476 32438 15528 32444
rect 15384 31884 15436 31890
rect 15384 31826 15436 31832
rect 15672 31822 15700 32846
rect 15764 32502 15792 32914
rect 15752 32496 15804 32502
rect 15752 32438 15804 32444
rect 15856 31890 15884 34342
rect 15844 31884 15896 31890
rect 15844 31826 15896 31832
rect 15660 31816 15712 31822
rect 15660 31758 15712 31764
rect 15856 29714 15884 31826
rect 15844 29708 15896 29714
rect 15844 29650 15896 29656
rect 15568 29096 15620 29102
rect 15568 29038 15620 29044
rect 15304 28966 15424 28994
rect 15292 28008 15344 28014
rect 15292 27950 15344 27956
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14188 22976 14240 22982
rect 14188 22918 14240 22924
rect 14200 20058 14228 22918
rect 14384 21486 14412 23122
rect 14476 21690 14504 24618
rect 15120 24342 15148 24618
rect 15304 24562 15332 27950
rect 15396 26246 15424 28966
rect 15580 26450 15608 29038
rect 15844 29028 15896 29034
rect 15844 28970 15896 28976
rect 15660 27532 15712 27538
rect 15660 27474 15712 27480
rect 15672 26586 15700 27474
rect 15660 26580 15712 26586
rect 15660 26522 15712 26528
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15384 26240 15436 26246
rect 15384 26182 15436 26188
rect 15476 25968 15528 25974
rect 15476 25910 15528 25916
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 15396 25362 15424 25638
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15212 24534 15332 24562
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14660 23798 14688 24142
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14476 21010 14504 21286
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14292 19922 14320 20946
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14384 20330 14412 20742
rect 14372 20324 14424 20330
rect 14372 20266 14424 20272
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 14476 20210 14504 20266
rect 14384 20182 14504 20210
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14016 18222 14044 18362
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13740 10130 13768 10746
rect 13832 10130 13860 14758
rect 13924 14260 13952 15982
rect 14016 15366 14044 16594
rect 14108 15638 14136 18158
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14200 17746 14228 18090
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14292 17626 14320 19178
rect 14384 18834 14412 20182
rect 14660 19258 14688 23734
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14752 22982 14780 23598
rect 14844 23582 15056 23610
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14844 20330 14872 23582
rect 15028 23526 15056 23582
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 14936 22642 14964 23462
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14936 21554 14964 22578
rect 15120 22148 15148 22918
rect 15028 22120 15148 22148
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14936 21078 14964 21490
rect 15028 21486 15056 22120
rect 15212 22080 15240 24534
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15304 22574 15332 24346
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15396 23186 15424 23598
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15120 22052 15240 22080
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 15028 21078 15056 21422
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 14936 20584 14964 21014
rect 15120 20806 15148 22052
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 15016 20596 15068 20602
rect 14936 20556 15016 20584
rect 14832 20324 14884 20330
rect 14752 20284 14832 20312
rect 14752 19446 14780 20284
rect 14832 20266 14884 20272
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14844 19334 14872 19994
rect 14476 19230 14688 19258
rect 14752 19306 14872 19334
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14200 17598 14320 17626
rect 14200 16590 14228 17598
rect 14476 17542 14504 19230
rect 14556 19168 14608 19174
rect 14752 19122 14780 19306
rect 14936 19242 14964 20556
rect 15016 20538 15068 20544
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15120 19922 15148 20198
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15120 19446 15148 19858
rect 15304 19786 15332 22374
rect 15396 22250 15424 23122
rect 15488 22438 15516 25910
rect 15580 25378 15608 26386
rect 15672 25498 15700 26522
rect 15856 26450 15884 28970
rect 15948 28694 15976 37318
rect 16405 37020 16713 37040
rect 16405 37018 16411 37020
rect 16467 37018 16491 37020
rect 16547 37018 16571 37020
rect 16627 37018 16651 37020
rect 16707 37018 16713 37020
rect 16467 36966 16469 37018
rect 16649 36966 16651 37018
rect 16405 36964 16411 36966
rect 16467 36964 16491 36966
rect 16547 36964 16571 36966
rect 16627 36964 16651 36966
rect 16707 36964 16713 36966
rect 16405 36944 16713 36964
rect 16405 35932 16713 35952
rect 16405 35930 16411 35932
rect 16467 35930 16491 35932
rect 16547 35930 16571 35932
rect 16627 35930 16651 35932
rect 16707 35930 16713 35932
rect 16467 35878 16469 35930
rect 16649 35878 16651 35930
rect 16405 35876 16411 35878
rect 16467 35876 16491 35878
rect 16547 35876 16571 35878
rect 16627 35876 16651 35878
rect 16707 35876 16713 35878
rect 16405 35856 16713 35876
rect 16405 34844 16713 34864
rect 16405 34842 16411 34844
rect 16467 34842 16491 34844
rect 16547 34842 16571 34844
rect 16627 34842 16651 34844
rect 16707 34842 16713 34844
rect 16467 34790 16469 34842
rect 16649 34790 16651 34842
rect 16405 34788 16411 34790
rect 16467 34788 16491 34790
rect 16547 34788 16571 34790
rect 16627 34788 16651 34790
rect 16707 34788 16713 34790
rect 16405 34768 16713 34788
rect 16212 34672 16264 34678
rect 16212 34614 16264 34620
rect 16224 34066 16252 34614
rect 16776 34474 16804 47942
rect 18328 47796 18380 47802
rect 18328 47738 18380 47744
rect 18052 47592 18104 47598
rect 18052 47534 18104 47540
rect 17868 47524 17920 47530
rect 17868 47466 17920 47472
rect 17684 47456 17736 47462
rect 17684 47398 17736 47404
rect 17408 47116 17460 47122
rect 17408 47058 17460 47064
rect 17316 46912 17368 46918
rect 17316 46854 17368 46860
rect 17328 46510 17356 46854
rect 17132 46504 17184 46510
rect 17132 46446 17184 46452
rect 17316 46504 17368 46510
rect 17316 46446 17368 46452
rect 16856 45280 16908 45286
rect 16856 45222 16908 45228
rect 16868 42158 16896 45222
rect 17040 45076 17092 45082
rect 17040 45018 17092 45024
rect 16948 44736 17000 44742
rect 16948 44678 17000 44684
rect 16960 44266 16988 44678
rect 17052 44334 17080 45018
rect 17144 44946 17172 46446
rect 17328 46034 17356 46446
rect 17420 46170 17448 47058
rect 17696 46510 17724 47398
rect 17880 46714 17908 47466
rect 18064 47122 18092 47534
rect 18052 47116 18104 47122
rect 18052 47058 18104 47064
rect 18340 46714 18368 47738
rect 19708 47456 19760 47462
rect 19708 47398 19760 47404
rect 19720 47122 19748 47398
rect 18788 47116 18840 47122
rect 18788 47058 18840 47064
rect 19708 47116 19760 47122
rect 19708 47058 19760 47064
rect 17868 46708 17920 46714
rect 17868 46650 17920 46656
rect 18328 46708 18380 46714
rect 18328 46650 18380 46656
rect 18340 46510 18368 46650
rect 17684 46504 17736 46510
rect 17684 46446 17736 46452
rect 18328 46504 18380 46510
rect 18328 46446 18380 46452
rect 17592 46436 17644 46442
rect 17592 46378 17644 46384
rect 17500 46368 17552 46374
rect 17500 46310 17552 46316
rect 17408 46164 17460 46170
rect 17408 46106 17460 46112
rect 17512 46102 17540 46310
rect 17500 46096 17552 46102
rect 17500 46038 17552 46044
rect 17316 46028 17368 46034
rect 17316 45970 17368 45976
rect 17132 44940 17184 44946
rect 17132 44882 17184 44888
rect 17144 44470 17172 44882
rect 17512 44878 17540 46038
rect 17604 45966 17632 46378
rect 17592 45960 17644 45966
rect 17592 45902 17644 45908
rect 17604 44878 17632 45902
rect 17696 44946 17724 46446
rect 18052 45824 18104 45830
rect 18052 45766 18104 45772
rect 17960 45348 18012 45354
rect 17960 45290 18012 45296
rect 17972 45082 18000 45290
rect 17960 45076 18012 45082
rect 17960 45018 18012 45024
rect 17684 44940 17736 44946
rect 17868 44940 17920 44946
rect 17736 44900 17868 44928
rect 17684 44882 17736 44888
rect 17868 44882 17920 44888
rect 17500 44872 17552 44878
rect 17500 44814 17552 44820
rect 17592 44872 17644 44878
rect 17592 44814 17644 44820
rect 17696 44817 17724 44882
rect 17512 44690 17540 44814
rect 17236 44662 17540 44690
rect 17132 44464 17184 44470
rect 17132 44406 17184 44412
rect 17040 44328 17092 44334
rect 17040 44270 17092 44276
rect 16948 44260 17000 44266
rect 16948 44202 17000 44208
rect 17144 43314 17172 44406
rect 17236 44198 17264 44662
rect 17604 44402 17632 44814
rect 18064 44538 18092 45766
rect 18052 44532 18104 44538
rect 18052 44474 18104 44480
rect 17592 44396 17644 44402
rect 17592 44338 17644 44344
rect 17960 44328 18012 44334
rect 17960 44270 18012 44276
rect 17316 44260 17368 44266
rect 17316 44202 17368 44208
rect 17224 44192 17276 44198
rect 17224 44134 17276 44140
rect 17236 43994 17264 44134
rect 17224 43988 17276 43994
rect 17224 43930 17276 43936
rect 16948 43308 17000 43314
rect 16948 43250 17000 43256
rect 17132 43308 17184 43314
rect 17132 43250 17184 43256
rect 16960 42770 16988 43250
rect 16948 42764 17000 42770
rect 16948 42706 17000 42712
rect 17236 42702 17264 43930
rect 17224 42696 17276 42702
rect 17224 42638 17276 42644
rect 17328 42566 17356 44202
rect 17592 44192 17644 44198
rect 17592 44134 17644 44140
rect 17684 44192 17736 44198
rect 17684 44134 17736 44140
rect 17604 43926 17632 44134
rect 17592 43920 17644 43926
rect 17592 43862 17644 43868
rect 17408 43104 17460 43110
rect 17408 43046 17460 43052
rect 17420 42634 17448 43046
rect 17696 42770 17724 44134
rect 17972 43994 18000 44270
rect 17960 43988 18012 43994
rect 17960 43930 18012 43936
rect 17776 43444 17828 43450
rect 17776 43386 17828 43392
rect 17500 42764 17552 42770
rect 17500 42706 17552 42712
rect 17684 42764 17736 42770
rect 17684 42706 17736 42712
rect 17408 42628 17460 42634
rect 17408 42570 17460 42576
rect 17316 42560 17368 42566
rect 17316 42502 17368 42508
rect 16856 42152 16908 42158
rect 16856 42094 16908 42100
rect 16948 42016 17000 42022
rect 17132 42016 17184 42022
rect 17000 41976 17080 42004
rect 16948 41958 17000 41964
rect 17052 41614 17080 41976
rect 17132 41958 17184 41964
rect 17040 41608 17092 41614
rect 17040 41550 17092 41556
rect 17052 41274 17080 41550
rect 16856 41268 16908 41274
rect 16856 41210 16908 41216
rect 17040 41268 17092 41274
rect 17040 41210 17092 41216
rect 16868 41138 16896 41210
rect 16856 41132 16908 41138
rect 16856 41074 16908 41080
rect 16948 41064 17000 41070
rect 16948 41006 17000 41012
rect 16960 40934 16988 41006
rect 16948 40928 17000 40934
rect 16948 40870 17000 40876
rect 16856 40588 16908 40594
rect 16856 40530 16908 40536
rect 16868 38962 16896 40530
rect 16960 39982 16988 40870
rect 17144 40662 17172 41958
rect 17316 41744 17368 41750
rect 17316 41686 17368 41692
rect 17224 41268 17276 41274
rect 17224 41210 17276 41216
rect 17236 41070 17264 41210
rect 17224 41064 17276 41070
rect 17224 41006 17276 41012
rect 17236 40730 17264 41006
rect 17328 41002 17356 41686
rect 17316 40996 17368 41002
rect 17316 40938 17368 40944
rect 17420 40730 17448 42570
rect 17512 42022 17540 42706
rect 17684 42560 17736 42566
rect 17684 42502 17736 42508
rect 17696 42158 17724 42502
rect 17684 42152 17736 42158
rect 17684 42094 17736 42100
rect 17500 42016 17552 42022
rect 17500 41958 17552 41964
rect 17788 41206 17816 43386
rect 17972 42702 18000 43930
rect 17960 42696 18012 42702
rect 17960 42638 18012 42644
rect 17960 42084 18012 42090
rect 17960 42026 18012 42032
rect 17776 41200 17828 41206
rect 17776 41142 17828 41148
rect 17972 41002 18000 42026
rect 17684 40996 17736 41002
rect 17684 40938 17736 40944
rect 17960 40996 18012 41002
rect 17960 40938 18012 40944
rect 17224 40724 17276 40730
rect 17224 40666 17276 40672
rect 17408 40724 17460 40730
rect 17408 40666 17460 40672
rect 17132 40656 17184 40662
rect 17132 40598 17184 40604
rect 17316 40588 17368 40594
rect 17316 40530 17368 40536
rect 17328 40186 17356 40530
rect 17316 40180 17368 40186
rect 17316 40122 17368 40128
rect 16948 39976 17000 39982
rect 16948 39918 17000 39924
rect 17132 39568 17184 39574
rect 17132 39510 17184 39516
rect 16856 38956 16908 38962
rect 16856 38898 16908 38904
rect 16856 38752 16908 38758
rect 16856 38694 16908 38700
rect 16868 37330 16896 38694
rect 16948 38480 17000 38486
rect 17000 38428 17080 38434
rect 16948 38422 17080 38428
rect 16960 38406 17080 38422
rect 16948 38208 17000 38214
rect 16948 38150 17000 38156
rect 16960 37806 16988 38150
rect 16948 37800 17000 37806
rect 16948 37742 17000 37748
rect 16948 37664 17000 37670
rect 16948 37606 17000 37612
rect 16856 37324 16908 37330
rect 16856 37266 16908 37272
rect 16960 36718 16988 37606
rect 17052 37398 17080 38406
rect 17040 37392 17092 37398
rect 17040 37334 17092 37340
rect 16948 36712 17000 36718
rect 16948 36654 17000 36660
rect 16856 36032 16908 36038
rect 16856 35974 16908 35980
rect 16868 35630 16896 35974
rect 16856 35624 16908 35630
rect 16856 35566 16908 35572
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16856 35216 16908 35222
rect 16856 35158 16908 35164
rect 16764 34468 16816 34474
rect 16764 34410 16816 34416
rect 16304 34400 16356 34406
rect 16304 34342 16356 34348
rect 16316 34134 16344 34342
rect 16304 34128 16356 34134
rect 16304 34070 16356 34076
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16405 33756 16713 33776
rect 16405 33754 16411 33756
rect 16467 33754 16491 33756
rect 16547 33754 16571 33756
rect 16627 33754 16651 33756
rect 16707 33754 16713 33756
rect 16467 33702 16469 33754
rect 16649 33702 16651 33754
rect 16405 33700 16411 33702
rect 16467 33700 16491 33702
rect 16547 33700 16571 33702
rect 16627 33700 16651 33702
rect 16707 33700 16713 33702
rect 16405 33680 16713 33700
rect 16304 33380 16356 33386
rect 16304 33322 16356 33328
rect 16764 33380 16816 33386
rect 16764 33322 16816 33328
rect 16028 33040 16080 33046
rect 16028 32982 16080 32988
rect 16040 32570 16068 32982
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 16028 32564 16080 32570
rect 16028 32506 16080 32512
rect 16224 32366 16252 32846
rect 16316 32502 16344 33322
rect 16405 32668 16713 32688
rect 16405 32666 16411 32668
rect 16467 32666 16491 32668
rect 16547 32666 16571 32668
rect 16627 32666 16651 32668
rect 16707 32666 16713 32668
rect 16467 32614 16469 32666
rect 16649 32614 16651 32666
rect 16405 32612 16411 32614
rect 16467 32612 16491 32614
rect 16547 32612 16571 32614
rect 16627 32612 16651 32614
rect 16707 32612 16713 32614
rect 16405 32592 16713 32612
rect 16304 32496 16356 32502
rect 16304 32438 16356 32444
rect 16580 32496 16632 32502
rect 16580 32438 16632 32444
rect 16316 32366 16344 32438
rect 16592 32366 16620 32438
rect 16776 32366 16804 33322
rect 16028 32360 16080 32366
rect 16028 32302 16080 32308
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 16304 32360 16356 32366
rect 16304 32302 16356 32308
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16764 32360 16816 32366
rect 16764 32302 16816 32308
rect 16040 31822 16068 32302
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16028 31816 16080 31822
rect 16028 31758 16080 31764
rect 16132 30054 16160 31826
rect 16316 30938 16344 32302
rect 16488 32292 16540 32298
rect 16488 32234 16540 32240
rect 16500 31958 16528 32234
rect 16592 31958 16620 32302
rect 16488 31952 16540 31958
rect 16488 31894 16540 31900
rect 16580 31952 16632 31958
rect 16580 31894 16632 31900
rect 16764 31884 16816 31890
rect 16764 31826 16816 31832
rect 16405 31580 16713 31600
rect 16405 31578 16411 31580
rect 16467 31578 16491 31580
rect 16547 31578 16571 31580
rect 16627 31578 16651 31580
rect 16707 31578 16713 31580
rect 16467 31526 16469 31578
rect 16649 31526 16651 31578
rect 16405 31524 16411 31526
rect 16467 31524 16491 31526
rect 16547 31524 16571 31526
rect 16627 31524 16651 31526
rect 16707 31524 16713 31526
rect 16405 31504 16713 31524
rect 16776 31414 16804 31826
rect 16764 31408 16816 31414
rect 16764 31350 16816 31356
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16776 30870 16804 31350
rect 16764 30864 16816 30870
rect 16764 30806 16816 30812
rect 16405 30492 16713 30512
rect 16405 30490 16411 30492
rect 16467 30490 16491 30492
rect 16547 30490 16571 30492
rect 16627 30490 16651 30492
rect 16707 30490 16713 30492
rect 16467 30438 16469 30490
rect 16649 30438 16651 30490
rect 16405 30436 16411 30438
rect 16467 30436 16491 30438
rect 16547 30436 16571 30438
rect 16627 30436 16651 30438
rect 16707 30436 16713 30438
rect 16405 30416 16713 30436
rect 16580 30252 16632 30258
rect 16580 30194 16632 30200
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 16132 29850 16160 29990
rect 16120 29844 16172 29850
rect 16120 29786 16172 29792
rect 16592 29782 16620 30194
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 16580 29776 16632 29782
rect 16580 29718 16632 29724
rect 16684 29714 16712 30126
rect 16672 29708 16724 29714
rect 16724 29668 16804 29696
rect 16672 29650 16724 29656
rect 16405 29404 16713 29424
rect 16405 29402 16411 29404
rect 16467 29402 16491 29404
rect 16547 29402 16571 29404
rect 16627 29402 16651 29404
rect 16707 29402 16713 29404
rect 16467 29350 16469 29402
rect 16649 29350 16651 29402
rect 16405 29348 16411 29350
rect 16467 29348 16491 29350
rect 16547 29348 16571 29350
rect 16627 29348 16651 29350
rect 16707 29348 16713 29350
rect 16405 29328 16713 29348
rect 16304 29300 16356 29306
rect 16304 29242 16356 29248
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 15936 28688 15988 28694
rect 15936 28630 15988 28636
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15948 27878 15976 28494
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 15948 27470 15976 27814
rect 15936 27464 15988 27470
rect 15936 27406 15988 27412
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15660 25492 15712 25498
rect 15660 25434 15712 25440
rect 15580 25350 15700 25378
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15580 24614 15608 25230
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15580 23186 15608 24550
rect 15672 23526 15700 25350
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15764 23186 15792 23666
rect 15856 23662 15884 26386
rect 15948 25362 15976 27406
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 15936 25356 15988 25362
rect 15936 25298 15988 25304
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 15844 23656 15896 23662
rect 15844 23598 15896 23604
rect 15568 23180 15620 23186
rect 15752 23180 15804 23186
rect 15568 23122 15620 23128
rect 15672 23140 15752 23168
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15396 22222 15608 22250
rect 15580 22030 15608 22222
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15580 21554 15608 21966
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15396 21010 15424 21490
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15488 20398 15516 21422
rect 15672 21350 15700 23140
rect 15752 23122 15804 23128
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15752 22568 15804 22574
rect 15752 22510 15804 22516
rect 15764 21486 15792 22510
rect 15856 22506 15884 23122
rect 15844 22500 15896 22506
rect 15844 22442 15896 22448
rect 15948 22386 15976 25162
rect 16040 24410 16068 26726
rect 16132 26042 16160 29106
rect 16316 28966 16344 29242
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16304 28960 16356 28966
rect 16304 28902 16356 28908
rect 16316 28014 16344 28902
rect 16684 28490 16712 29038
rect 16672 28484 16724 28490
rect 16672 28426 16724 28432
rect 16405 28316 16713 28336
rect 16405 28314 16411 28316
rect 16467 28314 16491 28316
rect 16547 28314 16571 28316
rect 16627 28314 16651 28316
rect 16707 28314 16713 28316
rect 16467 28262 16469 28314
rect 16649 28262 16651 28314
rect 16405 28260 16411 28262
rect 16467 28260 16491 28262
rect 16547 28260 16571 28262
rect 16627 28260 16651 28262
rect 16707 28260 16713 28262
rect 16405 28240 16713 28260
rect 16776 28218 16804 29668
rect 16868 29170 16896 35158
rect 16960 35154 16988 35430
rect 17144 35290 17172 39510
rect 17328 38486 17356 40122
rect 17420 38554 17448 40666
rect 17592 39976 17644 39982
rect 17592 39918 17644 39924
rect 17500 38956 17552 38962
rect 17500 38898 17552 38904
rect 17408 38548 17460 38554
rect 17408 38490 17460 38496
rect 17316 38480 17368 38486
rect 17316 38422 17368 38428
rect 17224 38412 17276 38418
rect 17224 38354 17276 38360
rect 17236 36242 17264 38354
rect 17420 37942 17448 38490
rect 17512 38418 17540 38898
rect 17500 38412 17552 38418
rect 17500 38354 17552 38360
rect 17512 37942 17540 38354
rect 17408 37936 17460 37942
rect 17408 37878 17460 37884
rect 17500 37936 17552 37942
rect 17500 37878 17552 37884
rect 17316 36576 17368 36582
rect 17316 36518 17368 36524
rect 17224 36236 17276 36242
rect 17224 36178 17276 36184
rect 17236 35494 17264 36178
rect 17328 35630 17356 36518
rect 17420 36310 17448 37878
rect 17512 36718 17540 37878
rect 17500 36712 17552 36718
rect 17500 36654 17552 36660
rect 17408 36304 17460 36310
rect 17408 36246 17460 36252
rect 17512 36242 17540 36654
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 17500 35692 17552 35698
rect 17500 35634 17552 35640
rect 17316 35624 17368 35630
rect 17316 35566 17368 35572
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17132 35284 17184 35290
rect 17132 35226 17184 35232
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 17328 34950 17356 35566
rect 17040 34944 17092 34950
rect 17040 34886 17092 34892
rect 17316 34944 17368 34950
rect 17316 34886 17368 34892
rect 17052 34746 17080 34886
rect 17512 34746 17540 35634
rect 17040 34740 17092 34746
rect 17040 34682 17092 34688
rect 17500 34740 17552 34746
rect 17500 34682 17552 34688
rect 17040 34468 17092 34474
rect 17040 34410 17092 34416
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16960 31142 16988 32166
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16960 29850 16988 31078
rect 16948 29844 17000 29850
rect 16948 29786 17000 29792
rect 16948 29708 17000 29714
rect 16948 29650 17000 29656
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16960 28778 16988 29650
rect 17052 29102 17080 34410
rect 17224 33856 17276 33862
rect 17224 33798 17276 33804
rect 17236 33590 17264 33798
rect 17224 33584 17276 33590
rect 17224 33526 17276 33532
rect 17236 32978 17264 33526
rect 17316 33312 17368 33318
rect 17316 33254 17368 33260
rect 17224 32972 17276 32978
rect 17144 32932 17224 32960
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 16868 28762 16988 28778
rect 16856 28756 16988 28762
rect 16908 28750 16988 28756
rect 16856 28698 16908 28704
rect 17144 28642 17172 32932
rect 17224 32914 17276 32920
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 17236 32366 17264 32506
rect 17328 32434 17356 33254
rect 17408 32768 17460 32774
rect 17408 32710 17460 32716
rect 17420 32570 17448 32710
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17512 32450 17540 34682
rect 17604 33046 17632 39918
rect 17696 39914 17724 40938
rect 18052 40656 18104 40662
rect 18052 40598 18104 40604
rect 17776 40520 17828 40526
rect 17776 40462 17828 40468
rect 17684 39908 17736 39914
rect 17684 39850 17736 39856
rect 17696 36378 17724 39850
rect 17788 38350 17816 40462
rect 17960 40384 18012 40390
rect 17960 40326 18012 40332
rect 17972 39982 18000 40326
rect 17960 39976 18012 39982
rect 17960 39918 18012 39924
rect 18064 39098 18092 40598
rect 18340 39574 18368 46446
rect 18800 46170 18828 47058
rect 18972 46912 19024 46918
rect 18972 46854 19024 46860
rect 18788 46164 18840 46170
rect 18788 46106 18840 46112
rect 18984 46034 19012 46854
rect 20088 46442 20116 47942
rect 21916 47592 21968 47598
rect 21916 47534 21968 47540
rect 20996 47524 21048 47530
rect 20996 47466 21048 47472
rect 20720 47184 20772 47190
rect 20720 47126 20772 47132
rect 20168 47116 20220 47122
rect 20168 47058 20220 47064
rect 19616 46436 19668 46442
rect 19616 46378 19668 46384
rect 20076 46436 20128 46442
rect 20076 46378 20128 46384
rect 18972 46028 19024 46034
rect 18972 45970 19024 45976
rect 19340 46028 19392 46034
rect 19340 45970 19392 45976
rect 19352 45286 19380 45970
rect 19628 45626 19656 46378
rect 19984 46368 20036 46374
rect 19984 46310 20036 46316
rect 19616 45620 19668 45626
rect 19616 45562 19668 45568
rect 18512 45280 18564 45286
rect 18512 45222 18564 45228
rect 18696 45280 18748 45286
rect 18696 45222 18748 45228
rect 19340 45280 19392 45286
rect 19340 45222 19392 45228
rect 18524 45082 18552 45222
rect 18512 45076 18564 45082
rect 18512 45018 18564 45024
rect 18708 44878 18736 45222
rect 18696 44872 18748 44878
rect 18696 44814 18748 44820
rect 18420 44396 18472 44402
rect 18420 44338 18472 44344
rect 18432 43314 18460 44338
rect 19432 44192 19484 44198
rect 19432 44134 19484 44140
rect 18972 43852 19024 43858
rect 18972 43794 19024 43800
rect 18512 43648 18564 43654
rect 18512 43590 18564 43596
rect 18420 43308 18472 43314
rect 18420 43250 18472 43256
rect 18524 42770 18552 43590
rect 18512 42764 18564 42770
rect 18512 42706 18564 42712
rect 18524 42226 18552 42706
rect 18512 42220 18564 42226
rect 18512 42162 18564 42168
rect 18524 40594 18552 42162
rect 18604 42016 18656 42022
rect 18604 41958 18656 41964
rect 18616 41614 18644 41958
rect 18604 41608 18656 41614
rect 18604 41550 18656 41556
rect 18616 41274 18644 41550
rect 18984 41414 19012 43794
rect 19340 43240 19392 43246
rect 19340 43182 19392 43188
rect 19352 42770 19380 43182
rect 19248 42764 19300 42770
rect 19248 42706 19300 42712
rect 19340 42764 19392 42770
rect 19340 42706 19392 42712
rect 18984 41386 19104 41414
rect 18604 41268 18656 41274
rect 18604 41210 18656 41216
rect 18616 40934 18644 41210
rect 18604 40928 18656 40934
rect 18604 40870 18656 40876
rect 18512 40588 18564 40594
rect 18512 40530 18564 40536
rect 18328 39568 18380 39574
rect 18328 39510 18380 39516
rect 18236 39500 18288 39506
rect 18236 39442 18288 39448
rect 18144 39296 18196 39302
rect 18144 39238 18196 39244
rect 18052 39092 18104 39098
rect 18052 39034 18104 39040
rect 17868 38820 17920 38826
rect 17868 38762 17920 38768
rect 17880 38554 17908 38762
rect 17868 38548 17920 38554
rect 17868 38490 17920 38496
rect 18156 38418 18184 39238
rect 18248 38554 18276 39442
rect 18512 39296 18564 39302
rect 18512 39238 18564 39244
rect 18524 38894 18552 39238
rect 18512 38888 18564 38894
rect 18512 38830 18564 38836
rect 18236 38548 18288 38554
rect 18236 38490 18288 38496
rect 18144 38412 18196 38418
rect 18064 38372 18144 38400
rect 17776 38344 17828 38350
rect 17776 38286 17828 38292
rect 17788 37874 17816 38286
rect 17776 37868 17828 37874
rect 17776 37810 17828 37816
rect 17788 36854 17816 37810
rect 17960 37732 18012 37738
rect 17960 37674 18012 37680
rect 17868 37664 17920 37670
rect 17868 37606 17920 37612
rect 17776 36848 17828 36854
rect 17776 36790 17828 36796
rect 17684 36372 17736 36378
rect 17684 36314 17736 36320
rect 17788 36242 17816 36790
rect 17880 36582 17908 37606
rect 17868 36576 17920 36582
rect 17868 36518 17920 36524
rect 17868 36304 17920 36310
rect 17868 36246 17920 36252
rect 17776 36236 17828 36242
rect 17776 36178 17828 36184
rect 17880 36174 17908 36246
rect 17972 36242 18000 37674
rect 17960 36236 18012 36242
rect 17960 36178 18012 36184
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 17972 35834 18000 36178
rect 18064 36106 18092 38372
rect 18144 38354 18196 38360
rect 18524 37806 18552 38830
rect 19076 38554 19104 41386
rect 19260 41274 19288 42706
rect 19352 41682 19380 42706
rect 19444 42362 19472 44134
rect 19524 42560 19576 42566
rect 19524 42502 19576 42508
rect 19432 42356 19484 42362
rect 19432 42298 19484 42304
rect 19536 42242 19564 42502
rect 19444 42214 19564 42242
rect 19340 41676 19392 41682
rect 19340 41618 19392 41624
rect 19340 41472 19392 41478
rect 19340 41414 19392 41420
rect 19248 41268 19300 41274
rect 19248 41210 19300 41216
rect 19248 41132 19300 41138
rect 19248 41074 19300 41080
rect 19260 40730 19288 41074
rect 19352 41002 19380 41414
rect 19444 41070 19472 42214
rect 19524 42016 19576 42022
rect 19524 41958 19576 41964
rect 19536 41206 19564 41958
rect 19524 41200 19576 41206
rect 19524 41142 19576 41148
rect 19432 41064 19484 41070
rect 19432 41006 19484 41012
rect 19340 40996 19392 41002
rect 19340 40938 19392 40944
rect 19248 40724 19300 40730
rect 19248 40666 19300 40672
rect 19260 39098 19288 40666
rect 19432 40588 19484 40594
rect 19484 40548 19564 40576
rect 19432 40530 19484 40536
rect 19536 39982 19564 40548
rect 19524 39976 19576 39982
rect 19524 39918 19576 39924
rect 19340 39908 19392 39914
rect 19340 39850 19392 39856
rect 19248 39092 19300 39098
rect 19248 39034 19300 39040
rect 19064 38548 19116 38554
rect 19064 38490 19116 38496
rect 18696 38412 18748 38418
rect 18696 38354 18748 38360
rect 18708 38010 18736 38354
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18512 37800 18564 37806
rect 18512 37742 18564 37748
rect 19064 37732 19116 37738
rect 19064 37674 19116 37680
rect 18236 37324 18288 37330
rect 18236 37266 18288 37272
rect 18144 36576 18196 36582
rect 18144 36518 18196 36524
rect 18052 36100 18104 36106
rect 18052 36042 18104 36048
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 17868 35760 17920 35766
rect 17868 35702 17920 35708
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17788 33318 17816 33934
rect 17776 33312 17828 33318
rect 17776 33254 17828 33260
rect 17592 33040 17644 33046
rect 17592 32982 17644 32988
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17420 32422 17540 32450
rect 17224 32360 17276 32366
rect 17224 32302 17276 32308
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17224 31816 17276 31822
rect 17224 31758 17276 31764
rect 16960 28614 17172 28642
rect 16856 28416 16908 28422
rect 16856 28358 16908 28364
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16304 28008 16356 28014
rect 16304 27950 16356 27956
rect 16212 27396 16264 27402
rect 16212 27338 16264 27344
rect 16224 26518 16252 27338
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16316 26858 16344 27270
rect 16405 27228 16713 27248
rect 16405 27226 16411 27228
rect 16467 27226 16491 27228
rect 16547 27226 16571 27228
rect 16627 27226 16651 27228
rect 16707 27226 16713 27228
rect 16467 27174 16469 27226
rect 16649 27174 16651 27226
rect 16405 27172 16411 27174
rect 16467 27172 16491 27174
rect 16547 27172 16571 27174
rect 16627 27172 16651 27174
rect 16707 27172 16713 27174
rect 16405 27152 16713 27172
rect 16776 26926 16804 28154
rect 16868 27538 16896 28358
rect 16856 27532 16908 27538
rect 16856 27474 16908 27480
rect 16868 27130 16896 27474
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16304 26852 16356 26858
rect 16304 26794 16356 26800
rect 16580 26852 16632 26858
rect 16580 26794 16632 26800
rect 16592 26518 16620 26794
rect 16212 26512 16264 26518
rect 16212 26454 16264 26460
rect 16580 26512 16632 26518
rect 16580 26454 16632 26460
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 16316 26246 16344 26318
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 16120 26036 16172 26042
rect 16120 25978 16172 25984
rect 16224 24954 16252 26182
rect 16405 26140 16713 26160
rect 16405 26138 16411 26140
rect 16467 26138 16491 26140
rect 16547 26138 16571 26140
rect 16627 26138 16651 26140
rect 16707 26138 16713 26140
rect 16467 26086 16469 26138
rect 16649 26086 16651 26138
rect 16405 26084 16411 26086
rect 16467 26084 16491 26086
rect 16547 26084 16571 26086
rect 16627 26084 16651 26086
rect 16707 26084 16713 26086
rect 16405 26064 16713 26084
rect 16776 25362 16804 26862
rect 16960 26466 16988 28614
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 16868 26450 16988 26466
rect 16856 26444 16988 26450
rect 16908 26438 16988 26444
rect 16856 26386 16908 26392
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16405 25052 16713 25072
rect 16405 25050 16411 25052
rect 16467 25050 16491 25052
rect 16547 25050 16571 25052
rect 16627 25050 16651 25052
rect 16707 25050 16713 25052
rect 16467 24998 16469 25050
rect 16649 24998 16651 25050
rect 16405 24996 16411 24998
rect 16467 24996 16491 24998
rect 16547 24996 16571 24998
rect 16627 24996 16651 24998
rect 16707 24996 16713 24998
rect 16405 24976 16713 24996
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 16040 23186 16068 24346
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 16040 22574 16068 22918
rect 16028 22568 16080 22574
rect 16028 22510 16080 22516
rect 15948 22358 16068 22386
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15672 20942 15700 21286
rect 15856 21026 15884 22170
rect 15764 20998 15884 21026
rect 15936 21004 15988 21010
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15396 19922 15424 20266
rect 15384 19916 15436 19922
rect 15436 19876 15516 19904
rect 15384 19858 15436 19864
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 15304 19122 15332 19722
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 14556 19110 14608 19116
rect 14568 18834 14596 19110
rect 14660 19094 14780 19122
rect 15212 19094 15332 19122
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14660 18408 14688 19094
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14660 18380 14872 18408
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14096 15632 14148 15638
rect 14096 15574 14148 15580
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 14004 14272 14056 14278
rect 13924 14232 14004 14260
rect 13924 13530 13952 14232
rect 14004 14214 14056 14220
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 14016 12306 14044 13874
rect 14108 13870 14136 14282
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14200 13716 14228 16526
rect 14108 13688 14228 13716
rect 14108 12628 14136 13688
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12782 14228 13126
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14108 12600 14228 12628
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13924 11830 13952 12106
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 14016 11150 14044 12242
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14108 10606 14136 12174
rect 14200 11014 14228 12600
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 8498 13676 8774
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13280 6820 13400 6848
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4690 13124 4966
rect 13188 4758 13216 5102
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13188 2582 13216 4014
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13280 2106 13308 6820
rect 13556 6746 13584 8366
rect 13648 8022 13676 8434
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13740 7546 13768 7890
rect 13924 7818 13952 10542
rect 14200 10538 14228 10950
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14016 9382 14044 10066
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13372 6718 13584 6746
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13004 1222 13032 2042
rect 13372 1562 13400 6718
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6254 13584 6598
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13464 4690 13492 6122
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13648 4146 13676 7142
rect 13832 4282 13860 7686
rect 13924 7274 13952 7754
rect 14016 7478 14044 8978
rect 14108 8634 14136 9930
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14016 6458 14044 6802
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14016 4826 14044 5714
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 14108 4078 14136 4150
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14200 3670 14228 8978
rect 14292 8906 14320 17206
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14384 16794 14412 17070
rect 14476 17066 14504 17478
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14568 16810 14596 18022
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14476 16782 14596 16810
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14384 16250 14412 16526
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14476 15162 14504 16782
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14384 14074 14412 14486
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12374 14412 12582
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14384 10266 14412 10474
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14384 8514 14412 9998
rect 14292 8486 14412 8514
rect 14292 6882 14320 8486
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14384 7546 14412 8298
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14292 6854 14412 6882
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 5710 14320 6734
rect 14384 6254 14412 6854
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14292 5166 14320 5646
rect 14384 5302 14412 6190
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13832 3058 13860 3470
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13832 1970 13860 2994
rect 14292 2650 14320 3946
rect 14384 3670 14412 4966
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13820 1964 13872 1970
rect 13820 1906 13872 1912
rect 13360 1556 13412 1562
rect 13360 1498 13412 1504
rect 13832 1494 13860 1906
rect 14372 1896 14424 1902
rect 14372 1838 14424 1844
rect 14384 1562 14412 1838
rect 14372 1556 14424 1562
rect 14372 1498 14424 1504
rect 13820 1488 13872 1494
rect 13820 1430 13872 1436
rect 14004 1420 14056 1426
rect 14004 1362 14056 1368
rect 13176 1352 13228 1358
rect 13176 1294 13228 1300
rect 12992 1216 13044 1222
rect 12992 1158 13044 1164
rect 13188 882 13216 1294
rect 14016 950 14044 1362
rect 14476 1018 14504 14894
rect 14568 11898 14596 16662
rect 14660 15570 14688 18226
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14660 14482 14688 15506
rect 14752 15434 14780 17002
rect 14844 16046 14872 18380
rect 14936 18290 14964 18770
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14924 18148 14976 18154
rect 14924 18090 14976 18096
rect 14936 16658 14964 18090
rect 15212 17954 15240 19094
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15304 18766 15332 18906
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15028 17926 15240 17954
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 13938 14688 14418
rect 14936 14278 14964 15914
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13462 14688 13738
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14660 12646 14688 13398
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14844 12782 14872 13330
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 15028 12458 15056 17926
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 15910 15148 17682
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15212 16250 15240 16594
rect 15304 16590 15332 17274
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15120 15366 15148 15574
rect 15212 15570 15240 16186
rect 15396 16096 15424 19450
rect 15488 18970 15516 19876
rect 15580 19360 15608 20878
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15580 19306 15617 19360
rect 15580 19224 15608 19306
rect 15580 19196 15617 19224
rect 15589 19156 15617 19196
rect 15580 19128 15617 19156
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15488 18290 15516 18906
rect 15580 18358 15608 19128
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15488 17202 15516 17614
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16250 15516 17002
rect 15580 16794 15608 18294
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15304 16068 15424 16096
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15304 15502 15332 16068
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15396 15706 15424 15914
rect 15580 15706 15608 16594
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15212 14550 15240 15098
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15304 14482 15332 15438
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15120 14056 15148 14418
rect 15120 14028 15240 14056
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15120 13190 15148 13874
rect 15212 13870 15240 14028
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15304 13394 15332 14418
rect 15396 14414 15424 15302
rect 15488 14482 15516 15370
rect 15672 15162 15700 20742
rect 15764 19258 15792 20998
rect 15936 20946 15988 20952
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15856 20330 15884 20878
rect 15948 20398 15976 20946
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15844 19916 15896 19922
rect 15896 19876 15976 19904
rect 15844 19858 15896 19864
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15856 19378 15884 19722
rect 15948 19446 15976 19876
rect 15936 19440 15988 19446
rect 15936 19382 15988 19388
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15764 19230 15884 19258
rect 15856 18850 15884 19230
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15764 18822 15884 18850
rect 15948 18834 15976 19110
rect 15936 18828 15988 18834
rect 15764 18086 15792 18822
rect 15936 18770 15988 18776
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15764 16998 15792 17750
rect 15856 17066 15884 18702
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15672 14890 15700 15098
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12782 15148 13126
rect 15304 12918 15332 13330
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15396 12850 15424 14350
rect 15488 13530 15516 14418
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 14660 12430 15056 12458
rect 15488 12442 15516 12650
rect 15476 12436 15528 12442
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14568 11218 14596 11834
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14568 10130 14596 10474
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14568 6458 14596 10066
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 4146 14596 5510
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14464 1012 14516 1018
rect 14464 954 14516 960
rect 14004 944 14056 950
rect 13176 876 13228 882
rect 13176 818 13228 824
rect 13832 870 13952 898
rect 14004 886 14056 892
rect 12900 808 12952 814
rect 2778 0 2834 800
rect 8298 0 8354 800
rect 13832 800 13860 870
rect 13924 814 13952 870
rect 13912 808 13964 814
rect 12900 750 12952 756
rect 9496 672 9548 678
rect 9496 614 9548 620
rect 9508 474 9536 614
rect 11253 572 11561 592
rect 11253 570 11259 572
rect 11315 570 11339 572
rect 11395 570 11419 572
rect 11475 570 11499 572
rect 11555 570 11561 572
rect 11315 518 11317 570
rect 11497 518 11499 570
rect 11253 516 11259 518
rect 11315 516 11339 518
rect 11395 516 11419 518
rect 11475 516 11499 518
rect 11555 516 11561 518
rect 11253 496 11561 516
rect 9496 468 9548 474
rect 9496 410 9548 416
rect 13818 0 13874 800
rect 13912 750 13964 756
rect 14660 678 14688 12430
rect 15476 12378 15528 12384
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 10062 14780 10542
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14844 9722 14872 10066
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14936 8786 14964 11154
rect 15028 9654 15056 11494
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 14752 8758 14964 8786
rect 14752 6934 14780 8758
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14844 7342 14872 8570
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 7546 14964 8298
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 15028 6866 15056 7890
rect 15120 7546 15148 10406
rect 15212 9496 15240 11698
rect 15200 9490 15252 9496
rect 15200 9432 15252 9438
rect 15292 9444 15344 9450
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15212 7392 15240 9432
rect 15292 9386 15344 9392
rect 15304 8294 15332 9386
rect 15488 8906 15516 12174
rect 15580 11608 15608 14826
rect 15764 14822 15792 16934
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15856 16590 15884 16730
rect 15948 16658 15976 18362
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15672 13462 15700 14554
rect 15764 13870 15792 14554
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15764 11778 15792 13806
rect 15856 11898 15884 16526
rect 15948 15570 15976 16594
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15948 12442 15976 14826
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15948 12170 15976 12378
rect 16040 12238 16068 22358
rect 16224 22098 16252 24142
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16316 23798 16344 24006
rect 16405 23964 16713 23984
rect 16405 23962 16411 23964
rect 16467 23962 16491 23964
rect 16547 23962 16571 23964
rect 16627 23962 16651 23964
rect 16707 23962 16713 23964
rect 16467 23910 16469 23962
rect 16649 23910 16651 23962
rect 16405 23908 16411 23910
rect 16467 23908 16491 23910
rect 16547 23908 16571 23910
rect 16627 23908 16651 23910
rect 16707 23908 16713 23910
rect 16405 23888 16713 23908
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16304 23588 16356 23594
rect 16304 23530 16356 23536
rect 16316 22760 16344 23530
rect 16405 22876 16713 22896
rect 16405 22874 16411 22876
rect 16467 22874 16491 22876
rect 16547 22874 16571 22876
rect 16627 22874 16651 22876
rect 16707 22874 16713 22876
rect 16467 22822 16469 22874
rect 16649 22822 16651 22874
rect 16405 22820 16411 22822
rect 16467 22820 16491 22822
rect 16547 22820 16571 22822
rect 16627 22820 16651 22822
rect 16707 22820 16713 22822
rect 16405 22800 16713 22820
rect 16316 22732 16528 22760
rect 16304 22500 16356 22506
rect 16304 22442 16356 22448
rect 16316 22166 16344 22442
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 16224 20942 16252 22034
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16132 19990 16160 20878
rect 16316 20534 16344 22102
rect 16500 22030 16528 22732
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16405 21788 16713 21808
rect 16405 21786 16411 21788
rect 16467 21786 16491 21788
rect 16547 21786 16571 21788
rect 16627 21786 16651 21788
rect 16707 21786 16713 21788
rect 16467 21734 16469 21786
rect 16649 21734 16651 21786
rect 16405 21732 16411 21734
rect 16467 21732 16491 21734
rect 16547 21732 16571 21734
rect 16627 21732 16651 21734
rect 16707 21732 16713 21734
rect 16405 21712 16713 21732
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16408 20874 16436 21422
rect 16592 21146 16620 21422
rect 16776 21146 16804 25094
rect 16868 23746 16896 26386
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16960 26042 16988 26318
rect 16948 26036 17000 26042
rect 16948 25978 17000 25984
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16960 24274 16988 25094
rect 17052 24682 17080 28426
rect 17144 28014 17172 28494
rect 17132 28008 17184 28014
rect 17132 27950 17184 27956
rect 17144 27538 17172 27950
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 17236 27418 17264 31758
rect 17328 31142 17356 32166
rect 17420 31822 17448 32422
rect 17880 32416 17908 35702
rect 18052 35624 18104 35630
rect 18052 35566 18104 35572
rect 18064 34542 18092 35566
rect 18052 34536 18104 34542
rect 18052 34478 18104 34484
rect 17960 34468 18012 34474
rect 17960 34410 18012 34416
rect 17972 32774 18000 34410
rect 17960 32768 18012 32774
rect 17960 32710 18012 32716
rect 18052 32496 18104 32502
rect 18052 32438 18104 32444
rect 17880 32388 18000 32416
rect 17972 32298 18000 32388
rect 17868 32292 17920 32298
rect 17868 32234 17920 32240
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 17500 31884 17552 31890
rect 17500 31826 17552 31832
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17316 31136 17368 31142
rect 17316 31078 17368 31084
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17328 28626 17356 30534
rect 17316 28620 17368 28626
rect 17316 28562 17368 28568
rect 17420 27962 17448 31758
rect 17512 31278 17540 31826
rect 17880 31362 17908 32234
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 17604 31334 17908 31362
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17500 31136 17552 31142
rect 17500 31078 17552 31084
rect 17512 30274 17540 31078
rect 17604 30394 17632 31334
rect 17684 31272 17736 31278
rect 17868 31272 17920 31278
rect 17736 31232 17816 31260
rect 17684 31214 17736 31220
rect 17684 30728 17736 30734
rect 17684 30670 17736 30676
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17512 30246 17632 30274
rect 17500 29776 17552 29782
rect 17500 29718 17552 29724
rect 17512 29034 17540 29718
rect 17500 29028 17552 29034
rect 17500 28970 17552 28976
rect 17512 28082 17540 28970
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 17420 27934 17540 27962
rect 17316 27532 17368 27538
rect 17316 27474 17368 27480
rect 17144 27390 17264 27418
rect 17144 26738 17172 27390
rect 17328 27334 17356 27474
rect 17316 27328 17368 27334
rect 17316 27270 17368 27276
rect 17512 27146 17540 27934
rect 17328 27118 17540 27146
rect 17144 26710 17264 26738
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 17144 26450 17172 26522
rect 17132 26444 17184 26450
rect 17132 26386 17184 26392
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16868 23718 16988 23746
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16868 22098 16896 23598
rect 16960 23322 16988 23718
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16868 21978 16896 22034
rect 16868 21950 16988 21978
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16396 20868 16448 20874
rect 16396 20810 16448 20816
rect 16405 20700 16713 20720
rect 16405 20698 16411 20700
rect 16467 20698 16491 20700
rect 16547 20698 16571 20700
rect 16627 20698 16651 20700
rect 16707 20698 16713 20700
rect 16467 20646 16469 20698
rect 16649 20646 16651 20698
rect 16405 20644 16411 20646
rect 16467 20644 16491 20646
rect 16547 20644 16571 20646
rect 16627 20644 16651 20646
rect 16707 20644 16713 20646
rect 16405 20624 16713 20644
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16120 19984 16172 19990
rect 16120 19926 16172 19932
rect 16132 19310 16160 19926
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16132 17814 16160 18566
rect 16224 18426 16252 19858
rect 16500 19700 16528 20470
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16592 19922 16620 20334
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16684 19854 16712 20198
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16316 19672 16528 19700
rect 16316 18834 16344 19672
rect 16405 19612 16713 19632
rect 16405 19610 16411 19612
rect 16467 19610 16491 19612
rect 16547 19610 16571 19612
rect 16627 19610 16651 19612
rect 16707 19610 16713 19612
rect 16467 19558 16469 19610
rect 16649 19558 16651 19610
rect 16405 19556 16411 19558
rect 16467 19556 16491 19558
rect 16547 19556 16571 19558
rect 16627 19556 16651 19558
rect 16707 19556 16713 19558
rect 16405 19536 16713 19556
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16408 18612 16436 19110
rect 16592 18698 16620 19178
rect 16684 18970 16712 19246
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16776 18714 16804 20946
rect 16868 20602 16896 21354
rect 16960 21350 16988 21950
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16868 18834 16896 19722
rect 17052 19666 17080 24618
rect 17144 23662 17172 25434
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17144 21434 17172 23462
rect 17236 22098 17264 26710
rect 17328 22522 17356 27118
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17420 24274 17448 26522
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17604 23594 17632 30246
rect 17696 29170 17724 30670
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17696 28694 17724 29106
rect 17684 28688 17736 28694
rect 17684 28630 17736 28636
rect 17696 27606 17724 28630
rect 17788 28558 17816 31232
rect 17972 31260 18000 31758
rect 17920 31232 18000 31260
rect 17868 31214 17920 31220
rect 18064 30938 18092 32438
rect 18156 31278 18184 36518
rect 18248 36378 18276 37266
rect 19076 37194 19104 37674
rect 19064 37188 19116 37194
rect 19064 37130 19116 37136
rect 18328 37120 18380 37126
rect 18328 37062 18380 37068
rect 18236 36372 18288 36378
rect 18236 36314 18288 36320
rect 18340 35766 18368 37062
rect 18880 36100 18932 36106
rect 18880 36042 18932 36048
rect 18328 35760 18380 35766
rect 18328 35702 18380 35708
rect 18340 34542 18368 35702
rect 18696 35080 18748 35086
rect 18696 35022 18748 35028
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18524 34610 18552 34886
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18328 34536 18380 34542
rect 18328 34478 18380 34484
rect 18340 34048 18368 34478
rect 18512 34128 18564 34134
rect 18512 34070 18564 34076
rect 18248 34020 18368 34048
rect 18248 31872 18276 34020
rect 18524 33454 18552 34070
rect 18604 33924 18656 33930
rect 18604 33866 18656 33872
rect 18512 33448 18564 33454
rect 18512 33390 18564 33396
rect 18524 33114 18552 33390
rect 18512 33108 18564 33114
rect 18512 33050 18564 33056
rect 18328 33040 18380 33046
rect 18328 32982 18380 32988
rect 18340 32230 18368 32982
rect 18524 32978 18552 33050
rect 18512 32972 18564 32978
rect 18512 32914 18564 32920
rect 18328 32224 18380 32230
rect 18328 32166 18380 32172
rect 18616 31958 18644 33866
rect 18604 31952 18656 31958
rect 18604 31894 18656 31900
rect 18248 31844 18368 31872
rect 18144 31272 18196 31278
rect 18144 31214 18196 31220
rect 18052 30932 18104 30938
rect 18052 30874 18104 30880
rect 18144 30864 18196 30870
rect 18144 30806 18196 30812
rect 18052 30796 18104 30802
rect 18052 30738 18104 30744
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17788 28218 17816 28358
rect 17776 28212 17828 28218
rect 17776 28154 17828 28160
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 17696 27470 17724 27542
rect 17788 27538 17816 28018
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17696 26994 17724 27406
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17788 26874 17816 27474
rect 17696 26846 17816 26874
rect 17696 26790 17724 26846
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17696 26586 17724 26726
rect 17779 26602 17807 26726
rect 17684 26580 17736 26586
rect 17779 26574 17816 26602
rect 17684 26522 17736 26528
rect 17788 25430 17816 26574
rect 17880 26450 17908 29446
rect 17972 28626 18000 30534
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 18064 28422 18092 30738
rect 18156 29850 18184 30806
rect 18144 29844 18196 29850
rect 18144 29786 18196 29792
rect 18156 28762 18184 29786
rect 18144 28756 18196 28762
rect 18144 28698 18196 28704
rect 18236 28688 18288 28694
rect 18236 28630 18288 28636
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 17972 28082 18000 28154
rect 18064 28082 18092 28358
rect 18248 28218 18276 28630
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17972 26450 18000 27882
rect 18064 27538 18092 28018
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18052 27532 18104 27538
rect 18052 27474 18104 27480
rect 18156 27470 18184 27950
rect 18144 27464 18196 27470
rect 18196 27424 18276 27452
rect 18144 27406 18196 27412
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 18052 26784 18104 26790
rect 18052 26726 18104 26732
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 17960 26444 18012 26450
rect 17960 26386 18012 26392
rect 18064 25974 18092 26726
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 18156 25838 18184 26862
rect 18248 26858 18276 27424
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18156 25498 18184 25774
rect 18144 25492 18196 25498
rect 18144 25434 18196 25440
rect 17776 25424 17828 25430
rect 17776 25366 17828 25372
rect 17684 24744 17736 24750
rect 17684 24686 17736 24692
rect 17592 23588 17644 23594
rect 17592 23530 17644 23536
rect 17500 22568 17552 22574
rect 17328 22494 17448 22522
rect 17500 22510 17552 22516
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17328 22098 17356 22374
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17236 21944 17264 22034
rect 17236 21916 17356 21944
rect 17144 21406 17264 21434
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17144 19922 17172 21286
rect 17236 20534 17264 21406
rect 17328 21078 17356 21916
rect 17316 21072 17368 21078
rect 17316 21014 17368 21020
rect 17328 20806 17356 21014
rect 17420 21010 17448 22494
rect 17512 22098 17540 22510
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 17604 21978 17632 23530
rect 17696 23526 17724 24686
rect 18156 24274 18184 25434
rect 18248 24274 18276 26794
rect 18340 24936 18368 31844
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18420 30660 18472 30666
rect 18420 30602 18472 30608
rect 18432 29238 18460 30602
rect 18420 29232 18472 29238
rect 18420 29174 18472 29180
rect 18524 28966 18552 31214
rect 18604 30116 18656 30122
rect 18604 30058 18656 30064
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 18432 26382 18460 26726
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18432 25838 18460 26318
rect 18524 25974 18552 28154
rect 18616 27606 18644 30058
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18340 24908 18460 24936
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18236 24268 18288 24274
rect 18236 24210 18288 24216
rect 18340 24206 18368 24754
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17512 21950 17632 21978
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 16960 19638 17080 19666
rect 16856 18828 16908 18834
rect 16960 18816 16988 19638
rect 17132 19440 17184 19446
rect 17236 19428 17264 20334
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17184 19400 17264 19428
rect 17316 19440 17368 19446
rect 17132 19382 17184 19388
rect 17316 19382 17368 19388
rect 17040 19304 17092 19310
rect 17328 19292 17356 19382
rect 17092 19264 17356 19292
rect 17040 19246 17092 19252
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18834 17356 19110
rect 17224 18828 17276 18834
rect 16960 18788 17080 18816
rect 16856 18770 16908 18776
rect 16580 18692 16632 18698
rect 16776 18686 16896 18714
rect 16580 18634 16632 18640
rect 16316 18584 16436 18612
rect 16764 18624 16816 18630
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16316 18154 16344 18584
rect 16764 18566 16816 18572
rect 16405 18524 16713 18544
rect 16405 18522 16411 18524
rect 16467 18522 16491 18524
rect 16547 18522 16571 18524
rect 16627 18522 16651 18524
rect 16707 18522 16713 18524
rect 16467 18470 16469 18522
rect 16649 18470 16651 18522
rect 16405 18468 16411 18470
rect 16467 18468 16491 18470
rect 16547 18468 16571 18470
rect 16627 18468 16651 18470
rect 16707 18468 16713 18470
rect 16405 18448 16713 18468
rect 16776 18222 16804 18566
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16132 16114 16160 17750
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 14074 16160 16050
rect 16224 16046 16252 18022
rect 16316 17134 16344 18090
rect 16684 18068 16712 18158
rect 16684 18040 16804 18068
rect 16405 17436 16713 17456
rect 16405 17434 16411 17436
rect 16467 17434 16491 17436
rect 16547 17434 16571 17436
rect 16627 17434 16651 17436
rect 16707 17434 16713 17436
rect 16467 17382 16469 17434
rect 16649 17382 16651 17434
rect 16405 17380 16411 17382
rect 16467 17380 16491 17382
rect 16547 17380 16571 17382
rect 16627 17380 16651 17382
rect 16707 17380 16713 17382
rect 16405 17360 16713 17380
rect 16776 17338 16804 18040
rect 16868 17610 16896 18686
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16960 17882 16988 18634
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16304 16448 16356 16454
rect 16408 16436 16436 17138
rect 16408 16408 16804 16436
rect 16304 16390 16356 16396
rect 16316 16114 16344 16390
rect 16405 16348 16713 16368
rect 16405 16346 16411 16348
rect 16467 16346 16491 16348
rect 16547 16346 16571 16348
rect 16627 16346 16651 16348
rect 16707 16346 16713 16348
rect 16467 16294 16469 16346
rect 16649 16294 16651 16346
rect 16405 16292 16411 16294
rect 16467 16292 16491 16294
rect 16547 16292 16571 16294
rect 16627 16292 16651 16294
rect 16707 16292 16713 16294
rect 16405 16272 16713 16292
rect 16776 16182 16804 16408
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15094 16252 15846
rect 16408 15706 16436 16118
rect 16672 15972 16724 15978
rect 16776 15960 16804 16118
rect 16868 16114 16896 17546
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16658 16988 16934
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16856 15972 16908 15978
rect 16776 15932 16856 15960
rect 16672 15914 16724 15920
rect 16856 15914 16908 15920
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16684 15570 16712 15914
rect 16672 15564 16724 15570
rect 16724 15524 16804 15552
rect 16672 15506 16724 15512
rect 16405 15260 16713 15280
rect 16405 15258 16411 15260
rect 16467 15258 16491 15260
rect 16547 15258 16571 15260
rect 16627 15258 16651 15260
rect 16707 15258 16713 15260
rect 16467 15206 16469 15258
rect 16649 15206 16651 15258
rect 16405 15204 16411 15206
rect 16467 15204 16491 15206
rect 16547 15204 16571 15206
rect 16627 15204 16651 15206
rect 16707 15204 16713 15206
rect 16405 15184 16713 15204
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16132 13394 16160 14010
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 16132 12986 16160 13194
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15764 11750 15884 11778
rect 15752 11620 15804 11626
rect 15580 11580 15752 11608
rect 15752 11562 15804 11568
rect 15856 11014 15884 11750
rect 15948 11218 15976 12106
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16040 11558 16068 12038
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 11354 16068 11494
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 16132 11098 16160 11834
rect 15948 11070 16160 11098
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15580 8634 15608 9590
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15304 8266 15424 8294
rect 15292 7404 15344 7410
rect 15212 7364 15292 7392
rect 15292 7346 15344 7352
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 6866 15148 7142
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15108 6860 15160 6866
rect 15304 6848 15332 7346
rect 15396 7342 15424 8266
rect 15672 7342 15700 9454
rect 15764 8838 15792 9862
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15764 8430 15792 8774
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15764 7886 15792 8366
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15384 7336 15436 7342
rect 15660 7336 15712 7342
rect 15436 7296 15516 7324
rect 15384 7278 15436 7284
rect 15384 6860 15436 6866
rect 15304 6820 15384 6848
rect 15108 6802 15160 6808
rect 15384 6802 15436 6808
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5846 15332 6054
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15396 5710 15424 6802
rect 15488 6798 15516 7296
rect 15660 7278 15712 7284
rect 15672 7002 15700 7278
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 5778 15516 6734
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15580 5778 15608 6598
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15028 5098 15056 5510
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 15212 3738 15240 4694
rect 15396 4146 15424 5646
rect 15580 4826 15608 5714
rect 15672 5642 15700 6802
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15672 5030 15700 5578
rect 15764 5166 15792 7822
rect 15948 6934 15976 11070
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 9518 16068 9998
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9586 16160 9862
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16132 9382 16160 9522
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16224 9110 16252 15030
rect 16776 14890 16804 15524
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 9382 16344 14758
rect 16868 14550 16896 15302
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16405 14172 16713 14192
rect 16405 14170 16411 14172
rect 16467 14170 16491 14172
rect 16547 14170 16571 14172
rect 16627 14170 16651 14172
rect 16707 14170 16713 14172
rect 16467 14118 16469 14170
rect 16649 14118 16651 14170
rect 16405 14116 16411 14118
rect 16467 14116 16491 14118
rect 16547 14116 16571 14118
rect 16627 14116 16651 14118
rect 16707 14116 16713 14118
rect 16405 14096 16713 14116
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16408 13394 16436 13874
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16500 13462 16528 13738
rect 16592 13530 16620 13942
rect 16672 13932 16724 13938
rect 16776 13920 16804 14350
rect 16868 14278 16896 14486
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16868 13938 16896 14010
rect 16960 13954 16988 15982
rect 17052 14958 17080 18788
rect 17224 18770 17276 18776
rect 17316 18828 17368 18834
rect 17420 18816 17448 19654
rect 17512 19174 17540 21950
rect 17696 21554 17724 23462
rect 17972 22574 18000 23802
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 18064 22030 18092 23054
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17592 20324 17644 20330
rect 17592 20266 17644 20272
rect 17604 19242 17632 20266
rect 17696 19990 17724 20470
rect 17972 20466 18000 21898
rect 18156 21690 18184 23598
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17684 19984 17736 19990
rect 18156 19938 18184 21082
rect 17684 19926 17736 19932
rect 18064 19910 18184 19938
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17592 19236 17644 19242
rect 17592 19178 17644 19184
rect 17880 19174 17908 19314
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17420 18788 17540 18816
rect 17316 18770 17368 18776
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17144 18340 17172 18702
rect 17236 18698 17264 18770
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17328 18426 17356 18566
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17224 18352 17276 18358
rect 17144 18312 17224 18340
rect 17224 18294 17276 18300
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17132 17808 17184 17814
rect 17132 17750 17184 17756
rect 17144 17134 17172 17750
rect 17236 17338 17264 18158
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17144 14362 17172 16934
rect 17420 16794 17448 18566
rect 17512 18340 17540 18788
rect 17696 18748 17724 18906
rect 17604 18720 17724 18748
rect 17604 18630 17632 18720
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17512 18312 17632 18340
rect 17604 18086 17632 18312
rect 17788 18306 17816 19110
rect 17696 18278 17816 18306
rect 17696 18222 17724 18278
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17604 17746 17632 18022
rect 17788 17814 17816 18158
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17604 17338 17632 17682
rect 17880 17660 17908 19110
rect 17696 17632 17908 17660
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17328 16114 17356 16186
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17052 14334 17172 14362
rect 17052 14056 17080 14334
rect 17132 14272 17184 14278
rect 17184 14232 17264 14260
rect 17132 14214 17184 14220
rect 17052 14028 17172 14056
rect 16724 13892 16804 13920
rect 16856 13932 16908 13938
rect 16672 13874 16724 13880
rect 16960 13926 17080 13954
rect 16856 13874 16908 13880
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16488 13456 16540 13462
rect 16488 13398 16540 13404
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16408 13258 16436 13330
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16405 13084 16713 13104
rect 16405 13082 16411 13084
rect 16467 13082 16491 13084
rect 16547 13082 16571 13084
rect 16627 13082 16651 13084
rect 16707 13082 16713 13084
rect 16467 13030 16469 13082
rect 16649 13030 16651 13082
rect 16405 13028 16411 13030
rect 16467 13028 16491 13030
rect 16547 13028 16571 13030
rect 16627 13028 16651 13030
rect 16707 13028 16713 13030
rect 16405 13008 16713 13028
rect 16776 12782 16804 13126
rect 16960 12782 16988 13398
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16405 11996 16713 12016
rect 16405 11994 16411 11996
rect 16467 11994 16491 11996
rect 16547 11994 16571 11996
rect 16627 11994 16651 11996
rect 16707 11994 16713 11996
rect 16467 11942 16469 11994
rect 16649 11942 16651 11994
rect 16405 11940 16411 11942
rect 16467 11940 16491 11942
rect 16547 11940 16571 11942
rect 16627 11940 16651 11942
rect 16707 11940 16713 11942
rect 16405 11920 16713 11940
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16868 11354 16896 11562
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16960 11286 16988 11494
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16405 10908 16713 10928
rect 16405 10906 16411 10908
rect 16467 10906 16491 10908
rect 16547 10906 16571 10908
rect 16627 10906 16651 10908
rect 16707 10906 16713 10908
rect 16467 10854 16469 10906
rect 16649 10854 16651 10906
rect 16405 10852 16411 10854
rect 16467 10852 16491 10854
rect 16547 10852 16571 10854
rect 16627 10852 16651 10854
rect 16707 10852 16713 10854
rect 16405 10832 16713 10852
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16405 9820 16713 9840
rect 16405 9818 16411 9820
rect 16467 9818 16491 9820
rect 16547 9818 16571 9820
rect 16627 9818 16651 9820
rect 16707 9818 16713 9820
rect 16467 9766 16469 9818
rect 16649 9766 16651 9818
rect 16405 9764 16411 9766
rect 16467 9764 16491 9766
rect 16547 9764 16571 9766
rect 16627 9764 16651 9766
rect 16707 9764 16713 9766
rect 16405 9744 16713 9764
rect 16776 9654 16804 10474
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16224 8430 16252 8842
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 7206 16160 7686
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15856 5778 15884 6802
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15948 5658 15976 6870
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16132 6458 16160 6734
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 15856 5630 15976 5658
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15488 4282 15516 4626
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15580 4078 15608 4762
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15672 2774 15700 4966
rect 15764 4690 15792 5102
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15672 2746 15792 2774
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14752 1970 14780 2382
rect 14740 1964 14792 1970
rect 14740 1906 14792 1912
rect 15396 1358 15424 2450
rect 15764 1902 15792 2746
rect 15752 1896 15804 1902
rect 15752 1838 15804 1844
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15856 1018 15884 5630
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16040 3194 16068 4014
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16040 2774 16068 3130
rect 15948 2746 16068 2774
rect 15948 2582 15976 2746
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15948 1562 15976 2314
rect 15936 1556 15988 1562
rect 15936 1498 15988 1504
rect 15844 1012 15896 1018
rect 15844 954 15896 960
rect 15948 814 15976 1498
rect 16040 1358 16068 2382
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 16040 882 16068 1294
rect 16132 1018 16160 3878
rect 16224 1766 16252 8366
rect 16316 7528 16344 9114
rect 16868 8922 16896 9862
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16776 8894 16896 8922
rect 16405 8732 16713 8752
rect 16405 8730 16411 8732
rect 16467 8730 16491 8732
rect 16547 8730 16571 8732
rect 16627 8730 16651 8732
rect 16707 8730 16713 8732
rect 16467 8678 16469 8730
rect 16649 8678 16651 8730
rect 16405 8676 16411 8678
rect 16467 8676 16491 8678
rect 16547 8676 16571 8678
rect 16627 8676 16651 8678
rect 16707 8676 16713 8678
rect 16405 8656 16713 8676
rect 16776 8072 16804 8894
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16684 8044 16804 8072
rect 16684 7818 16712 8044
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16405 7644 16713 7664
rect 16405 7642 16411 7644
rect 16467 7642 16491 7644
rect 16547 7642 16571 7644
rect 16627 7642 16651 7644
rect 16707 7642 16713 7644
rect 16467 7590 16469 7642
rect 16649 7590 16651 7642
rect 16405 7588 16411 7590
rect 16467 7588 16491 7590
rect 16547 7588 16571 7590
rect 16627 7588 16651 7590
rect 16707 7588 16713 7590
rect 16405 7568 16713 7588
rect 16776 7546 16804 7890
rect 16764 7540 16816 7546
rect 16316 7500 16436 7528
rect 16408 7410 16436 7500
rect 16764 7482 16816 7488
rect 16868 7478 16896 8774
rect 16960 8566 16988 9318
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17052 8362 17080 13926
rect 17144 12594 17172 14028
rect 17236 13802 17264 14232
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17236 13394 17264 13738
rect 17236 13388 17288 13394
rect 17236 13330 17288 13336
rect 17236 12782 17264 13330
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17144 12566 17264 12594
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 10674 17172 11630
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17144 9450 17172 10610
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 17236 9042 17264 12566
rect 17328 9178 17356 16050
rect 17420 16046 17448 16594
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17420 13258 17448 14282
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17420 12374 17448 12718
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11150 17448 12038
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17316 8900 17368 8906
rect 17316 8842 17368 8848
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16960 7954 16988 8230
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16960 7410 16988 7890
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16316 6730 16344 7346
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16405 6556 16713 6576
rect 16405 6554 16411 6556
rect 16467 6554 16491 6556
rect 16547 6554 16571 6556
rect 16627 6554 16651 6556
rect 16707 6554 16713 6556
rect 16467 6502 16469 6554
rect 16649 6502 16651 6554
rect 16405 6500 16411 6502
rect 16467 6500 16491 6502
rect 16547 6500 16571 6502
rect 16627 6500 16651 6502
rect 16707 6500 16713 6502
rect 16405 6480 16713 6500
rect 16776 6186 16804 7278
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16868 6458 16896 6802
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16868 6254 16896 6394
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16684 5914 16712 6054
rect 16960 5930 16988 7210
rect 17052 6866 17080 8298
rect 17144 7546 17172 8502
rect 17328 8362 17356 8842
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17052 6458 17080 6802
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16868 5914 16988 5930
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16856 5908 16988 5914
rect 16908 5902 16988 5908
rect 16856 5850 16908 5856
rect 16405 5468 16713 5488
rect 16405 5466 16411 5468
rect 16467 5466 16491 5468
rect 16547 5466 16571 5468
rect 16627 5466 16651 5468
rect 16707 5466 16713 5468
rect 16467 5414 16469 5466
rect 16649 5414 16651 5466
rect 16405 5412 16411 5414
rect 16467 5412 16491 5414
rect 16547 5412 16571 5414
rect 16627 5412 16651 5414
rect 16707 5412 16713 5414
rect 16405 5392 16713 5412
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16316 4078 16344 4558
rect 16405 4380 16713 4400
rect 16405 4378 16411 4380
rect 16467 4378 16491 4380
rect 16547 4378 16571 4380
rect 16627 4378 16651 4380
rect 16707 4378 16713 4380
rect 16467 4326 16469 4378
rect 16649 4326 16651 4378
rect 16405 4324 16411 4326
rect 16467 4324 16491 4326
rect 16547 4324 16571 4326
rect 16627 4324 16651 4326
rect 16707 4324 16713 4326
rect 16405 4304 16713 4324
rect 16776 4146 16804 4966
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16405 3292 16713 3312
rect 16405 3290 16411 3292
rect 16467 3290 16491 3292
rect 16547 3290 16571 3292
rect 16627 3290 16651 3292
rect 16707 3290 16713 3292
rect 16467 3238 16469 3290
rect 16649 3238 16651 3290
rect 16405 3236 16411 3238
rect 16467 3236 16491 3238
rect 16547 3236 16571 3238
rect 16627 3236 16651 3238
rect 16707 3236 16713 3238
rect 16405 3216 16713 3236
rect 16776 3194 16804 3538
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16684 2650 16712 2858
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16405 2204 16713 2224
rect 16405 2202 16411 2204
rect 16467 2202 16491 2204
rect 16547 2202 16571 2204
rect 16627 2202 16651 2204
rect 16707 2202 16713 2204
rect 16467 2150 16469 2202
rect 16649 2150 16651 2202
rect 16405 2148 16411 2150
rect 16467 2148 16491 2150
rect 16547 2148 16571 2150
rect 16627 2148 16651 2150
rect 16707 2148 16713 2150
rect 16405 2128 16713 2148
rect 16868 2106 16896 4966
rect 16960 4078 16988 5902
rect 17144 5302 17172 7346
rect 17236 7002 17264 7754
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17144 4196 17172 5238
rect 17236 5234 17264 6938
rect 17328 6390 17356 8298
rect 17420 7342 17448 10950
rect 17512 10742 17540 17274
rect 17604 17134 17632 17274
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17604 16046 17632 16730
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17604 13462 17632 15370
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17696 12434 17724 17632
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17788 16028 17816 16934
rect 17880 16794 17908 17138
rect 17972 17134 18000 19450
rect 18064 18154 18092 19910
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18156 18834 18184 19790
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17972 16658 18000 17070
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 18064 16250 18092 17614
rect 18156 16726 18184 18770
rect 18248 17814 18276 23258
rect 18340 21690 18368 24142
rect 18432 22710 18460 24908
rect 18524 23118 18552 25910
rect 18616 25838 18644 27270
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18616 25226 18644 25774
rect 18604 25220 18656 25226
rect 18604 25162 18656 25168
rect 18616 24274 18644 25162
rect 18708 24750 18736 35022
rect 18788 34944 18840 34950
rect 18788 34886 18840 34892
rect 18800 33658 18828 34886
rect 18788 33652 18840 33658
rect 18788 33594 18840 33600
rect 18788 33312 18840 33318
rect 18788 33254 18840 33260
rect 18800 32230 18828 33254
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 18800 27674 18828 31894
rect 18892 31346 18920 36042
rect 18972 35556 19024 35562
rect 18972 35498 19024 35504
rect 18984 34678 19012 35498
rect 19076 35154 19104 37130
rect 19156 36032 19208 36038
rect 19156 35974 19208 35980
rect 19064 35148 19116 35154
rect 19064 35090 19116 35096
rect 18972 34672 19024 34678
rect 18972 34614 19024 34620
rect 19168 34184 19196 35974
rect 19352 35894 19380 39850
rect 19536 39794 19564 39918
rect 19628 39914 19656 45562
rect 19800 45280 19852 45286
rect 19800 45222 19852 45228
rect 19812 44946 19840 45222
rect 19800 44940 19852 44946
rect 19800 44882 19852 44888
rect 19996 41414 20024 46310
rect 20180 46034 20208 47058
rect 20628 46980 20680 46986
rect 20628 46922 20680 46928
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 20180 45286 20208 45970
rect 20352 45960 20404 45966
rect 20352 45902 20404 45908
rect 20364 45830 20392 45902
rect 20352 45824 20404 45830
rect 20352 45766 20404 45772
rect 20168 45280 20220 45286
rect 20168 45222 20220 45228
rect 20364 43994 20392 45766
rect 20640 44198 20668 46922
rect 20732 46374 20760 47126
rect 20812 46436 20864 46442
rect 20812 46378 20864 46384
rect 20720 46368 20772 46374
rect 20720 46310 20772 46316
rect 20732 45422 20760 46310
rect 20824 46170 20852 46378
rect 20812 46164 20864 46170
rect 20812 46106 20864 46112
rect 20812 46028 20864 46034
rect 20812 45970 20864 45976
rect 20720 45416 20772 45422
rect 20720 45358 20772 45364
rect 20824 45370 20852 45970
rect 20904 45824 20956 45830
rect 20904 45766 20956 45772
rect 20916 45490 20944 45766
rect 21008 45558 21036 47466
rect 21557 47356 21865 47376
rect 21557 47354 21563 47356
rect 21619 47354 21643 47356
rect 21699 47354 21723 47356
rect 21779 47354 21803 47356
rect 21859 47354 21865 47356
rect 21619 47302 21621 47354
rect 21801 47302 21803 47354
rect 21557 47300 21563 47302
rect 21619 47300 21643 47302
rect 21699 47300 21723 47302
rect 21779 47300 21803 47302
rect 21859 47300 21865 47302
rect 21557 47280 21865 47300
rect 21456 47116 21508 47122
rect 21456 47058 21508 47064
rect 21272 47048 21324 47054
rect 21272 46990 21324 46996
rect 21088 46912 21140 46918
rect 21088 46854 21140 46860
rect 21100 45830 21128 46854
rect 21284 45966 21312 46990
rect 21364 46980 21416 46986
rect 21364 46922 21416 46928
rect 21272 45960 21324 45966
rect 21272 45902 21324 45908
rect 21088 45824 21140 45830
rect 21088 45766 21140 45772
rect 20996 45552 21048 45558
rect 20996 45494 21048 45500
rect 20904 45484 20956 45490
rect 20904 45426 20956 45432
rect 20628 44192 20680 44198
rect 20628 44134 20680 44140
rect 20352 43988 20404 43994
rect 20352 43930 20404 43936
rect 20260 43852 20312 43858
rect 20260 43794 20312 43800
rect 20168 43648 20220 43654
rect 20168 43590 20220 43596
rect 20076 42560 20128 42566
rect 20076 42502 20128 42508
rect 20088 41562 20116 42502
rect 20180 42090 20208 43590
rect 20168 42084 20220 42090
rect 20168 42026 20220 42032
rect 20272 41682 20300 43794
rect 20364 43246 20392 43930
rect 20536 43852 20588 43858
rect 20536 43794 20588 43800
rect 20444 43784 20496 43790
rect 20444 43726 20496 43732
rect 20352 43240 20404 43246
rect 20352 43182 20404 43188
rect 20260 41676 20312 41682
rect 20312 41636 20392 41664
rect 20260 41618 20312 41624
rect 20088 41534 20300 41562
rect 19996 41386 20208 41414
rect 20076 41132 20128 41138
rect 20076 41074 20128 41080
rect 19708 40928 19760 40934
rect 19708 40870 19760 40876
rect 19616 39908 19668 39914
rect 19616 39850 19668 39856
rect 19536 39766 19656 39794
rect 19628 39438 19656 39766
rect 19720 39574 19748 40870
rect 20088 40390 20116 41074
rect 20076 40384 20128 40390
rect 20076 40326 20128 40332
rect 19708 39568 19760 39574
rect 19708 39510 19760 39516
rect 19616 39432 19668 39438
rect 19616 39374 19668 39380
rect 19628 39302 19656 39374
rect 19616 39296 19668 39302
rect 19616 39238 19668 39244
rect 19432 38888 19484 38894
rect 19432 38830 19484 38836
rect 19444 37806 19472 38830
rect 19628 38350 19656 39238
rect 19800 39024 19852 39030
rect 19800 38966 19852 38972
rect 19708 38752 19760 38758
rect 19708 38694 19760 38700
rect 19616 38344 19668 38350
rect 19616 38286 19668 38292
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19628 37330 19656 38286
rect 19720 37806 19748 38694
rect 19812 37874 19840 38966
rect 19984 38888 20036 38894
rect 20088 38876 20116 40326
rect 20036 38848 20116 38876
rect 19984 38830 20036 38836
rect 20076 38412 20128 38418
rect 20076 38354 20128 38360
rect 20088 38010 20116 38354
rect 20076 38004 20128 38010
rect 20076 37946 20128 37952
rect 19800 37868 19852 37874
rect 19800 37810 19852 37816
rect 19708 37800 19760 37806
rect 19708 37742 19760 37748
rect 19616 37324 19668 37330
rect 19616 37266 19668 37272
rect 19524 36916 19576 36922
rect 19524 36858 19576 36864
rect 19260 35866 19380 35894
rect 19260 35834 19288 35866
rect 19536 35834 19564 36858
rect 19248 35828 19300 35834
rect 19248 35770 19300 35776
rect 19524 35828 19576 35834
rect 19524 35770 19576 35776
rect 19248 35624 19300 35630
rect 19248 35566 19300 35572
rect 19260 34542 19288 35566
rect 19524 35556 19576 35562
rect 19524 35498 19576 35504
rect 19340 35216 19392 35222
rect 19340 35158 19392 35164
rect 19248 34536 19300 34542
rect 19248 34478 19300 34484
rect 18984 34156 19288 34184
rect 18984 32570 19012 34156
rect 19156 34060 19208 34066
rect 19156 34002 19208 34008
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 19076 32892 19104 33866
rect 19168 33454 19196 34002
rect 19260 33522 19288 34156
rect 19352 33998 19380 35158
rect 19536 34202 19564 35498
rect 19628 34610 19656 37266
rect 19720 36854 19748 37742
rect 19800 37732 19852 37738
rect 19800 37674 19852 37680
rect 19708 36848 19760 36854
rect 19708 36790 19760 36796
rect 19812 36718 19840 37674
rect 19892 37324 19944 37330
rect 19892 37266 19944 37272
rect 19904 36922 19932 37266
rect 19892 36916 19944 36922
rect 19892 36858 19944 36864
rect 19800 36712 19852 36718
rect 19800 36654 19852 36660
rect 20180 36174 20208 41386
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 19800 35488 19852 35494
rect 19800 35430 19852 35436
rect 19812 35154 19840 35430
rect 19800 35148 19852 35154
rect 19800 35090 19852 35096
rect 19708 35080 19760 35086
rect 19708 35022 19760 35028
rect 19616 34604 19668 34610
rect 19616 34546 19668 34552
rect 19524 34196 19576 34202
rect 19524 34138 19576 34144
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 19720 33862 19748 35022
rect 19812 34066 19840 35090
rect 19984 35080 20036 35086
rect 19904 35040 19984 35068
rect 19904 34134 19932 35040
rect 19984 35022 20036 35028
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 19892 34128 19944 34134
rect 19892 34070 19944 34076
rect 19800 34060 19852 34066
rect 19800 34002 19852 34008
rect 19708 33856 19760 33862
rect 19708 33798 19760 33804
rect 19812 33658 19840 34002
rect 19904 33930 19932 34070
rect 19892 33924 19944 33930
rect 19892 33866 19944 33872
rect 19800 33652 19852 33658
rect 19800 33594 19852 33600
rect 19248 33516 19300 33522
rect 19248 33458 19300 33464
rect 19156 33448 19208 33454
rect 19432 33448 19484 33454
rect 19156 33390 19208 33396
rect 19352 33408 19432 33436
rect 19352 32978 19380 33408
rect 19800 33448 19852 33454
rect 19628 33408 19800 33436
rect 19628 33402 19656 33408
rect 19432 33390 19484 33396
rect 19536 33374 19656 33402
rect 19800 33390 19852 33396
rect 19536 33318 19564 33374
rect 19524 33312 19576 33318
rect 19524 33254 19576 33260
rect 19708 33312 19760 33318
rect 19708 33254 19760 33260
rect 19616 33040 19668 33046
rect 19616 32982 19668 32988
rect 19340 32972 19392 32978
rect 19340 32914 19392 32920
rect 19156 32904 19208 32910
rect 19076 32864 19156 32892
rect 19156 32846 19208 32852
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19248 32836 19300 32842
rect 19248 32778 19300 32784
rect 19156 32768 19208 32774
rect 19076 32728 19156 32756
rect 18972 32564 19024 32570
rect 18972 32506 19024 32512
rect 18972 32224 19024 32230
rect 19076 32212 19104 32728
rect 19156 32710 19208 32716
rect 19156 32292 19208 32298
rect 19156 32234 19208 32240
rect 19024 32184 19104 32212
rect 18972 32166 19024 32172
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18984 31210 19012 31758
rect 18972 31204 19024 31210
rect 18972 31146 19024 31152
rect 18984 30258 19012 31146
rect 19168 30870 19196 32234
rect 19260 31346 19288 32778
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19156 30864 19208 30870
rect 19156 30806 19208 30812
rect 19260 30598 19288 31282
rect 19444 30666 19472 32846
rect 19628 32774 19656 32982
rect 19720 32978 19748 33254
rect 19708 32972 19760 32978
rect 19708 32914 19760 32920
rect 19800 32972 19852 32978
rect 19904 32960 19932 33866
rect 19996 33522 20024 34614
rect 20076 34060 20128 34066
rect 20128 34020 20208 34048
rect 20076 34002 20128 34008
rect 20180 33862 20208 34020
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 19984 33516 20036 33522
rect 19984 33458 20036 33464
rect 20076 33448 20128 33454
rect 20076 33390 20128 33396
rect 19852 32932 19932 32960
rect 19800 32914 19852 32920
rect 19616 32768 19668 32774
rect 19812 32756 19840 32914
rect 19984 32768 20036 32774
rect 19812 32728 19932 32756
rect 19616 32710 19668 32716
rect 19708 32564 19760 32570
rect 19708 32506 19760 32512
rect 19720 32366 19748 32506
rect 19708 32360 19760 32366
rect 19708 32302 19760 32308
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19720 31278 19748 31826
rect 19708 31272 19760 31278
rect 19708 31214 19760 31220
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19064 30320 19116 30326
rect 19064 30262 19116 30268
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 18880 29844 18932 29850
rect 18880 29786 18932 29792
rect 18788 27668 18840 27674
rect 18788 27610 18840 27616
rect 18892 26858 18920 29786
rect 18984 29646 19012 30194
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18984 29170 19012 29582
rect 18972 29164 19024 29170
rect 18972 29106 19024 29112
rect 18972 27600 19024 27606
rect 18972 27542 19024 27548
rect 18880 26852 18932 26858
rect 18880 26794 18932 26800
rect 18880 25764 18932 25770
rect 18880 25706 18932 25712
rect 18788 25356 18840 25362
rect 18788 25298 18840 25304
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18432 22574 18460 22646
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18616 22522 18644 22918
rect 18708 22642 18736 24686
rect 18800 24410 18828 25298
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18340 18970 18368 21490
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 18340 18426 18368 18634
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18248 16640 18276 17478
rect 18340 17270 18368 18158
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18248 16612 18368 16640
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18156 16114 18184 16526
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 17868 16040 17920 16046
rect 17788 16000 17868 16028
rect 18052 16040 18104 16046
rect 17868 15982 17920 15988
rect 17972 16000 18052 16028
rect 17972 15570 18000 16000
rect 18052 15982 18104 15988
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 18064 14550 18092 15846
rect 18248 15570 18276 16458
rect 18340 16114 18368 16612
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18156 15162 18184 15506
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18144 14952 18196 14958
rect 18248 14940 18276 15506
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18340 14958 18368 15030
rect 18196 14912 18276 14940
rect 18328 14952 18380 14958
rect 18144 14894 18196 14900
rect 18328 14894 18380 14900
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 17776 14408 17828 14414
rect 17828 14356 18092 14362
rect 17776 14350 18092 14356
rect 17788 14334 18092 14350
rect 17788 12986 17816 14334
rect 18064 14278 18092 14334
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17972 13870 18000 14214
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13258 18092 13806
rect 18156 13530 18184 14894
rect 18432 14890 18460 22510
rect 18616 22494 18736 22522
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18616 21486 18644 22034
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18524 20942 18552 21354
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18524 20534 18552 20878
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18524 20398 18552 20470
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18524 19378 18552 20334
rect 18616 19922 18644 20946
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18616 19514 18644 19858
rect 18708 19786 18736 22494
rect 18800 22094 18828 24074
rect 18892 23322 18920 25706
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18800 22066 18920 22094
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18800 21554 18828 21966
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18800 21010 18828 21490
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18892 20534 18920 22066
rect 18880 20528 18932 20534
rect 18880 20470 18932 20476
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 18892 19904 18920 20266
rect 18984 20058 19012 27542
rect 19076 27538 19104 30262
rect 19260 30190 19288 30534
rect 19248 30184 19300 30190
rect 19248 30126 19300 30132
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19352 29714 19380 29990
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19352 29306 19380 29650
rect 19812 29306 19840 31962
rect 19904 31822 19932 32728
rect 19984 32710 20036 32716
rect 19892 31816 19944 31822
rect 19892 31758 19944 31764
rect 19996 30326 20024 32710
rect 20088 32434 20116 33390
rect 20180 32978 20208 33798
rect 20168 32972 20220 32978
rect 20168 32914 20220 32920
rect 20168 32768 20220 32774
rect 20168 32710 20220 32716
rect 20180 32502 20208 32710
rect 20168 32496 20220 32502
rect 20168 32438 20220 32444
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 20168 31884 20220 31890
rect 20168 31826 20220 31832
rect 20180 31482 20208 31826
rect 20168 31476 20220 31482
rect 20168 31418 20220 31424
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 20076 30320 20128 30326
rect 20076 30262 20128 30268
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 19812 28626 19840 29242
rect 19984 29028 20036 29034
rect 19984 28970 20036 28976
rect 19892 28960 19944 28966
rect 19892 28902 19944 28908
rect 19800 28620 19852 28626
rect 19800 28562 19852 28568
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19168 27606 19196 28358
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19156 27600 19208 27606
rect 19156 27542 19208 27548
rect 19064 27532 19116 27538
rect 19064 27474 19116 27480
rect 19076 27062 19104 27474
rect 19168 27130 19196 27542
rect 19260 27538 19288 27814
rect 19248 27532 19300 27538
rect 19248 27474 19300 27480
rect 19444 27470 19472 28086
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19800 28008 19852 28014
rect 19800 27950 19852 27956
rect 19628 27674 19656 27950
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19616 27668 19668 27674
rect 19616 27610 19668 27616
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19156 27124 19208 27130
rect 19156 27066 19208 27072
rect 19064 27056 19116 27062
rect 19064 26998 19116 27004
rect 19536 26858 19564 27610
rect 19812 27130 19840 27950
rect 19800 27124 19852 27130
rect 19800 27066 19852 27072
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 19524 26852 19576 26858
rect 19524 26794 19576 26800
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18972 19916 19024 19922
rect 18892 19876 18972 19904
rect 18972 19858 19024 19864
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18616 18834 18644 19178
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18708 18408 18736 19722
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18708 18380 18828 18408
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18524 17542 18552 18090
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18616 17542 18644 17818
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18524 15042 18552 17002
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18616 16046 18644 16594
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18616 15162 18644 15982
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18524 15014 18644 15042
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18248 13734 18276 14758
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 17880 12714 18000 12730
rect 17880 12708 18012 12714
rect 17880 12702 17960 12708
rect 17880 12434 17908 12702
rect 17960 12650 18012 12656
rect 18064 12646 18092 12922
rect 18156 12782 18184 13126
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 17696 12406 17908 12434
rect 18144 12436 18196 12442
rect 17696 11558 17724 12406
rect 18144 12378 18196 12384
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17880 11694 17908 12242
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17972 10606 18000 12310
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10266 17540 10406
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17512 9518 17540 10202
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17500 9376 17552 9382
rect 17604 9364 17632 9998
rect 17972 9654 18000 10542
rect 18064 10266 18092 12242
rect 18156 11014 18184 12378
rect 18248 11626 18276 12582
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18156 10606 18184 10950
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17552 9336 17632 9364
rect 17500 9318 17552 9324
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17512 7206 17540 9318
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17604 8022 17632 9114
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17696 7698 17724 8978
rect 17868 8968 17920 8974
rect 17788 8928 17868 8956
rect 17788 8566 17816 8928
rect 17868 8910 17920 8916
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17604 7670 17724 7698
rect 17604 7426 17632 7670
rect 17788 7478 17816 8366
rect 17880 7698 17908 8774
rect 17972 8430 18000 8774
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17880 7670 17917 7698
rect 17889 7528 17917 7670
rect 17880 7500 17917 7528
rect 17776 7472 17828 7478
rect 17604 7398 17724 7426
rect 17776 7414 17828 7420
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17316 6384 17368 6390
rect 17316 6326 17368 6332
rect 17328 5778 17356 6326
rect 17420 5914 17448 7142
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17420 5166 17448 5646
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17512 4690 17540 7142
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17604 6458 17632 6666
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17224 4208 17276 4214
rect 17144 4168 17224 4196
rect 17224 4150 17276 4156
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16960 3670 16988 4014
rect 17040 4004 17092 4010
rect 17040 3946 17092 3952
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 17052 2310 17080 3946
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 16856 2100 16908 2106
rect 16856 2042 16908 2048
rect 16212 1760 16264 1766
rect 16212 1702 16264 1708
rect 16948 1760 17000 1766
rect 16948 1702 17000 1708
rect 16764 1420 16816 1426
rect 16764 1362 16816 1368
rect 16405 1116 16713 1136
rect 16405 1114 16411 1116
rect 16467 1114 16491 1116
rect 16547 1114 16571 1116
rect 16627 1114 16651 1116
rect 16707 1114 16713 1116
rect 16467 1062 16469 1114
rect 16649 1062 16651 1114
rect 16405 1060 16411 1062
rect 16467 1060 16491 1062
rect 16547 1060 16571 1062
rect 16627 1060 16651 1062
rect 16707 1060 16713 1062
rect 16405 1040 16713 1060
rect 16120 1012 16172 1018
rect 16120 954 16172 960
rect 16028 876 16080 882
rect 16028 818 16080 824
rect 16776 814 16804 1362
rect 16960 814 16988 1702
rect 17132 1284 17184 1290
rect 17236 1272 17264 2586
rect 17328 1766 17356 2926
rect 17420 2514 17448 4558
rect 17512 3942 17540 4626
rect 17604 4146 17632 6394
rect 17696 5370 17724 7398
rect 17880 6798 17908 7500
rect 17972 7342 18000 8230
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5778 17816 6122
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17604 3534 17632 4082
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17696 3738 17724 4014
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17880 3398 17908 5850
rect 17972 5794 18000 7278
rect 18064 6848 18092 8298
rect 18156 8294 18184 8978
rect 18248 8566 18276 10678
rect 18340 8906 18368 13874
rect 18432 13802 18460 14826
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18432 12434 18460 13738
rect 18432 12406 18552 12434
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18432 12238 18460 12310
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18432 11558 18460 12174
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 10606 18460 11494
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18524 8906 18552 12406
rect 18616 11830 18644 15014
rect 18708 12374 18736 18226
rect 18800 17134 18828 18380
rect 18892 18154 18920 18770
rect 18880 18148 18932 18154
rect 18880 18090 18932 18096
rect 18984 18034 19012 19858
rect 18892 18006 19012 18034
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18800 16590 18828 17070
rect 18892 16998 18920 18006
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18892 16658 18920 16934
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18800 13462 18828 16186
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18892 12434 18920 16050
rect 18984 15570 19012 17818
rect 19076 17066 19104 26794
rect 19708 26444 19760 26450
rect 19708 26386 19760 26392
rect 19340 26308 19392 26314
rect 19340 26250 19392 26256
rect 19352 24834 19380 26250
rect 19720 26042 19748 26386
rect 19708 26036 19760 26042
rect 19760 25996 19840 26024
rect 19708 25978 19760 25984
rect 19260 24806 19380 24834
rect 19260 24290 19288 24806
rect 19812 24750 19840 25996
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19352 24410 19380 24686
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19524 24404 19576 24410
rect 19524 24346 19576 24352
rect 19260 24262 19380 24290
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19168 23866 19196 24142
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 19352 23746 19380 24262
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19444 23866 19472 24210
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19352 23718 19472 23746
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19352 22250 19380 23462
rect 19444 22658 19472 23718
rect 19536 22778 19564 24346
rect 19628 24206 19656 24686
rect 19904 24274 19932 28902
rect 19996 28762 20024 28970
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 20088 28150 20116 30262
rect 20168 29640 20220 29646
rect 20168 29582 20220 29588
rect 20180 29102 20208 29582
rect 20168 29096 20220 29102
rect 20168 29038 20220 29044
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 19996 27470 20024 27542
rect 20180 27538 20208 28562
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 19996 26382 20024 27406
rect 20088 27130 20116 27406
rect 20076 27124 20128 27130
rect 20076 27066 20128 27072
rect 20088 26908 20116 27066
rect 20180 27062 20208 27474
rect 20168 27056 20220 27062
rect 20168 26998 20220 27004
rect 20088 26880 20208 26908
rect 20180 26382 20208 26880
rect 20272 26568 20300 41534
rect 20364 41070 20392 41636
rect 20456 41206 20484 43726
rect 20548 42634 20576 43794
rect 20536 42628 20588 42634
rect 20536 42570 20588 42576
rect 20548 41818 20576 42570
rect 20732 42158 20760 45358
rect 20824 45342 20944 45370
rect 20812 44192 20864 44198
rect 20812 44134 20864 44140
rect 20720 42152 20772 42158
rect 20720 42094 20772 42100
rect 20536 41812 20588 41818
rect 20536 41754 20588 41760
rect 20444 41200 20496 41206
rect 20444 41142 20496 41148
rect 20456 41070 20484 41142
rect 20352 41064 20404 41070
rect 20352 41006 20404 41012
rect 20444 41064 20496 41070
rect 20444 41006 20496 41012
rect 20364 38826 20392 41006
rect 20456 39030 20484 41006
rect 20720 39908 20772 39914
rect 20720 39850 20772 39856
rect 20628 39840 20680 39846
rect 20628 39782 20680 39788
rect 20536 39500 20588 39506
rect 20536 39442 20588 39448
rect 20548 39098 20576 39442
rect 20640 39302 20668 39782
rect 20628 39296 20680 39302
rect 20628 39238 20680 39244
rect 20536 39092 20588 39098
rect 20536 39034 20588 39040
rect 20444 39024 20496 39030
rect 20444 38966 20496 38972
rect 20536 38888 20588 38894
rect 20536 38830 20588 38836
rect 20352 38820 20404 38826
rect 20352 38762 20404 38768
rect 20352 38548 20404 38554
rect 20352 38490 20404 38496
rect 20364 32314 20392 38490
rect 20548 38010 20576 38830
rect 20536 38004 20588 38010
rect 20536 37946 20588 37952
rect 20732 37942 20760 39850
rect 20824 38570 20852 44134
rect 20916 42838 20944 45342
rect 21180 45348 21232 45354
rect 21180 45290 21232 45296
rect 21192 45082 21220 45290
rect 21180 45076 21232 45082
rect 21180 45018 21232 45024
rect 21284 45014 21312 45902
rect 21272 45008 21324 45014
rect 21272 44950 21324 44956
rect 21088 44872 21140 44878
rect 21088 44814 21140 44820
rect 21100 43790 21128 44814
rect 21272 44328 21324 44334
rect 21272 44270 21324 44276
rect 21284 43858 21312 44270
rect 21376 43858 21404 46922
rect 21468 45898 21496 47058
rect 21928 46986 21956 47534
rect 22560 47524 22612 47530
rect 22560 47466 22612 47472
rect 22376 47456 22428 47462
rect 22376 47398 22428 47404
rect 22388 47122 22416 47398
rect 22572 47258 22600 47466
rect 24492 47456 24544 47462
rect 24492 47398 24544 47404
rect 22560 47252 22612 47258
rect 22560 47194 22612 47200
rect 23848 47184 23900 47190
rect 23848 47126 23900 47132
rect 22008 47116 22060 47122
rect 22008 47058 22060 47064
rect 22376 47116 22428 47122
rect 22376 47058 22428 47064
rect 21916 46980 21968 46986
rect 21916 46922 21968 46928
rect 21928 46578 21956 46922
rect 21916 46572 21968 46578
rect 21916 46514 21968 46520
rect 21928 46374 21956 46514
rect 22020 46374 22048 47058
rect 22560 47048 22612 47054
rect 22560 46990 22612 46996
rect 21916 46368 21968 46374
rect 21916 46310 21968 46316
rect 22008 46368 22060 46374
rect 22008 46310 22060 46316
rect 21557 46268 21865 46288
rect 21557 46266 21563 46268
rect 21619 46266 21643 46268
rect 21699 46266 21723 46268
rect 21779 46266 21803 46268
rect 21859 46266 21865 46268
rect 21619 46214 21621 46266
rect 21801 46214 21803 46266
rect 21557 46212 21563 46214
rect 21619 46212 21643 46214
rect 21699 46212 21723 46214
rect 21779 46212 21803 46214
rect 21859 46212 21865 46214
rect 21557 46192 21865 46212
rect 21928 45966 21956 46310
rect 22020 46170 22048 46310
rect 22008 46164 22060 46170
rect 22008 46106 22060 46112
rect 22284 46096 22336 46102
rect 22284 46038 22336 46044
rect 22100 46028 22152 46034
rect 22100 45970 22152 45976
rect 21548 45960 21600 45966
rect 21548 45902 21600 45908
rect 21916 45960 21968 45966
rect 21916 45902 21968 45908
rect 21456 45892 21508 45898
rect 21456 45834 21508 45840
rect 21468 45558 21496 45834
rect 21456 45552 21508 45558
rect 21456 45494 21508 45500
rect 21468 44946 21496 45494
rect 21560 45400 21588 45902
rect 21640 45824 21692 45830
rect 21640 45766 21692 45772
rect 21916 45824 21968 45830
rect 21916 45766 21968 45772
rect 21652 45422 21680 45766
rect 21640 45416 21692 45422
rect 21548 45394 21600 45400
rect 21640 45358 21692 45364
rect 21548 45336 21600 45342
rect 21557 45180 21865 45200
rect 21557 45178 21563 45180
rect 21619 45178 21643 45180
rect 21699 45178 21723 45180
rect 21779 45178 21803 45180
rect 21859 45178 21865 45180
rect 21619 45126 21621 45178
rect 21801 45126 21803 45178
rect 21557 45124 21563 45126
rect 21619 45124 21643 45126
rect 21699 45124 21723 45126
rect 21779 45124 21803 45126
rect 21859 45124 21865 45126
rect 21557 45104 21865 45124
rect 21456 44940 21508 44946
rect 21456 44882 21508 44888
rect 21468 44470 21496 44882
rect 21456 44464 21508 44470
rect 21456 44406 21508 44412
rect 21456 44192 21508 44198
rect 21456 44134 21508 44140
rect 21272 43852 21324 43858
rect 21272 43794 21324 43800
rect 21364 43852 21416 43858
rect 21364 43794 21416 43800
rect 21088 43784 21140 43790
rect 21088 43726 21140 43732
rect 21100 43382 21128 43726
rect 21088 43376 21140 43382
rect 21088 43318 21140 43324
rect 20904 42832 20956 42838
rect 20904 42774 20956 42780
rect 20996 42696 21048 42702
rect 20996 42638 21048 42644
rect 21008 41274 21036 42638
rect 20996 41268 21048 41274
rect 20996 41210 21048 41216
rect 21008 39114 21036 41210
rect 21100 41206 21128 43318
rect 21284 42362 21312 43794
rect 21364 42832 21416 42838
rect 21364 42774 21416 42780
rect 21272 42356 21324 42362
rect 21272 42298 21324 42304
rect 21272 41676 21324 41682
rect 21272 41618 21324 41624
rect 21284 41274 21312 41618
rect 21272 41268 21324 41274
rect 21272 41210 21324 41216
rect 21088 41200 21140 41206
rect 21088 41142 21140 41148
rect 21180 40724 21232 40730
rect 21180 40666 21232 40672
rect 21192 40390 21220 40666
rect 21180 40384 21232 40390
rect 21180 40326 21232 40332
rect 21192 39982 21220 40326
rect 21180 39976 21232 39982
rect 21180 39918 21232 39924
rect 20916 39086 21036 39114
rect 20916 38962 20944 39086
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 20916 38758 20944 38898
rect 21180 38888 21232 38894
rect 21180 38830 21232 38836
rect 20904 38752 20956 38758
rect 20904 38694 20956 38700
rect 20824 38542 20944 38570
rect 20720 37936 20772 37942
rect 20720 37878 20772 37884
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20628 35148 20680 35154
rect 20628 35090 20680 35096
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20456 34474 20484 34886
rect 20444 34468 20496 34474
rect 20444 34410 20496 34416
rect 20640 34406 20668 35090
rect 20720 34468 20772 34474
rect 20720 34410 20772 34416
rect 20536 34400 20588 34406
rect 20536 34342 20588 34348
rect 20628 34400 20680 34406
rect 20628 34342 20680 34348
rect 20548 33930 20576 34342
rect 20640 34134 20668 34342
rect 20732 34202 20760 34410
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20628 34128 20680 34134
rect 20628 34070 20680 34076
rect 20536 33924 20588 33930
rect 20536 33866 20588 33872
rect 20536 33652 20588 33658
rect 20536 33594 20588 33600
rect 20548 33386 20576 33594
rect 20640 33522 20668 34070
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20536 33380 20588 33386
rect 20536 33322 20588 33328
rect 20824 33318 20852 35974
rect 20916 33454 20944 38542
rect 21192 38214 21220 38830
rect 21180 38208 21232 38214
rect 21180 38150 21232 38156
rect 21192 37874 21220 38150
rect 21180 37868 21232 37874
rect 21180 37810 21232 37816
rect 21088 37800 21140 37806
rect 21088 37742 21140 37748
rect 20996 37664 21048 37670
rect 20996 37606 21048 37612
rect 21008 37466 21036 37606
rect 21100 37466 21128 37742
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 21088 37460 21140 37466
rect 21088 37402 21140 37408
rect 21192 37398 21220 37810
rect 21180 37392 21232 37398
rect 21180 37334 21232 37340
rect 21088 36848 21140 36854
rect 21088 36790 21140 36796
rect 20996 35556 21048 35562
rect 20996 35498 21048 35504
rect 20904 33448 20956 33454
rect 20904 33390 20956 33396
rect 20628 33312 20680 33318
rect 20812 33312 20864 33318
rect 20680 33260 20760 33266
rect 20628 33254 20760 33260
rect 20812 33254 20864 33260
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 20640 33238 20760 33254
rect 20732 32978 20760 33238
rect 20536 32972 20588 32978
rect 20536 32914 20588 32920
rect 20720 32972 20772 32978
rect 20720 32914 20772 32920
rect 20444 32836 20496 32842
rect 20444 32778 20496 32784
rect 20456 32434 20484 32778
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20364 32298 20484 32314
rect 20364 32292 20496 32298
rect 20364 32286 20444 32292
rect 20444 32234 20496 32240
rect 20456 31754 20484 32234
rect 20548 32026 20576 32914
rect 20824 32774 20852 33254
rect 20916 32978 20944 33254
rect 20904 32972 20956 32978
rect 20904 32914 20956 32920
rect 20812 32768 20864 32774
rect 20812 32710 20864 32716
rect 20628 32496 20680 32502
rect 21008 32450 21036 35498
rect 20628 32438 20680 32444
rect 20640 32298 20668 32438
rect 20916 32422 21036 32450
rect 20628 32292 20680 32298
rect 20628 32234 20680 32240
rect 20536 32020 20588 32026
rect 20536 31962 20588 31968
rect 20640 31890 20668 32234
rect 20720 32020 20772 32026
rect 20720 31962 20772 31968
rect 20628 31884 20680 31890
rect 20628 31826 20680 31832
rect 20732 31770 20760 31962
rect 20640 31754 20760 31770
rect 20456 31726 20576 31754
rect 20444 31680 20496 31686
rect 20444 31622 20496 31628
rect 20456 31278 20484 31622
rect 20444 31272 20496 31278
rect 20444 31214 20496 31220
rect 20352 30184 20404 30190
rect 20352 30126 20404 30132
rect 20364 28558 20392 30126
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20456 28626 20484 29582
rect 20444 28620 20496 28626
rect 20444 28562 20496 28568
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20548 28218 20576 31726
rect 20628 31748 20760 31754
rect 20680 31742 20760 31748
rect 20628 31690 20680 31696
rect 20640 30802 20668 31690
rect 20628 30796 20680 30802
rect 20628 30738 20680 30744
rect 20720 30660 20772 30666
rect 20720 30602 20772 30608
rect 20732 30190 20760 30602
rect 20720 30184 20772 30190
rect 20720 30126 20772 30132
rect 20732 29578 20760 30126
rect 20720 29572 20772 29578
rect 20720 29514 20772 29520
rect 20628 28688 20680 28694
rect 20628 28630 20680 28636
rect 20536 28212 20588 28218
rect 20536 28154 20588 28160
rect 20640 27538 20668 28630
rect 20628 27532 20680 27538
rect 20628 27474 20680 27480
rect 20640 27130 20668 27474
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20732 26858 20760 26930
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 20272 26540 20576 26568
rect 20548 26450 20576 26540
rect 20732 26518 20760 26794
rect 20824 26586 20852 27406
rect 20916 26858 20944 32422
rect 20996 32360 21048 32366
rect 20996 32302 21048 32308
rect 21008 32026 21036 32302
rect 20996 32020 21048 32026
rect 20996 31962 21048 31968
rect 21008 31890 21036 31962
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 21100 29510 21128 36790
rect 21284 36650 21312 41210
rect 21376 39030 21404 42774
rect 21468 42226 21496 44134
rect 21557 44092 21865 44112
rect 21557 44090 21563 44092
rect 21619 44090 21643 44092
rect 21699 44090 21723 44092
rect 21779 44090 21803 44092
rect 21859 44090 21865 44092
rect 21619 44038 21621 44090
rect 21801 44038 21803 44090
rect 21557 44036 21563 44038
rect 21619 44036 21643 44038
rect 21699 44036 21723 44038
rect 21779 44036 21803 44038
rect 21859 44036 21865 44038
rect 21557 44016 21865 44036
rect 21557 43004 21865 43024
rect 21557 43002 21563 43004
rect 21619 43002 21643 43004
rect 21699 43002 21723 43004
rect 21779 43002 21803 43004
rect 21859 43002 21865 43004
rect 21619 42950 21621 43002
rect 21801 42950 21803 43002
rect 21557 42948 21563 42950
rect 21619 42948 21643 42950
rect 21699 42948 21723 42950
rect 21779 42948 21803 42950
rect 21859 42948 21865 42950
rect 21557 42928 21865 42948
rect 21456 42220 21508 42226
rect 21456 42162 21508 42168
rect 21824 42152 21876 42158
rect 21928 42140 21956 45766
rect 22112 45014 22140 45970
rect 22296 45558 22324 46038
rect 22376 46028 22428 46034
rect 22376 45970 22428 45976
rect 22284 45552 22336 45558
rect 22284 45494 22336 45500
rect 22192 45280 22244 45286
rect 22192 45222 22244 45228
rect 22100 45008 22152 45014
rect 22100 44950 22152 44956
rect 22204 44946 22232 45222
rect 22008 44940 22060 44946
rect 22008 44882 22060 44888
rect 22192 44940 22244 44946
rect 22192 44882 22244 44888
rect 22020 44334 22048 44882
rect 22388 44742 22416 45970
rect 22376 44736 22428 44742
rect 22376 44678 22428 44684
rect 22572 44538 22600 46990
rect 23756 46640 23808 46646
rect 23756 46582 23808 46588
rect 23480 46572 23532 46578
rect 23480 46514 23532 46520
rect 23112 46436 23164 46442
rect 23112 46378 23164 46384
rect 23124 45422 23152 46378
rect 23492 45558 23520 46514
rect 23664 46368 23716 46374
rect 23664 46310 23716 46316
rect 23480 45552 23532 45558
rect 23480 45494 23532 45500
rect 23112 45416 23164 45422
rect 23112 45358 23164 45364
rect 23296 45416 23348 45422
rect 23296 45358 23348 45364
rect 23124 44946 23152 45358
rect 23112 44940 23164 44946
rect 23112 44882 23164 44888
rect 22560 44532 22612 44538
rect 22560 44474 22612 44480
rect 22100 44396 22152 44402
rect 22100 44338 22152 44344
rect 22192 44396 22244 44402
rect 22192 44338 22244 44344
rect 22008 44328 22060 44334
rect 22008 44270 22060 44276
rect 22112 43722 22140 44338
rect 22204 43790 22232 44338
rect 22284 44192 22336 44198
rect 22284 44134 22336 44140
rect 22376 44192 22428 44198
rect 22376 44134 22428 44140
rect 22192 43784 22244 43790
rect 22192 43726 22244 43732
rect 22100 43716 22152 43722
rect 22100 43658 22152 43664
rect 21876 42112 21956 42140
rect 21824 42094 21876 42100
rect 21557 41916 21865 41936
rect 21557 41914 21563 41916
rect 21619 41914 21643 41916
rect 21699 41914 21723 41916
rect 21779 41914 21803 41916
rect 21859 41914 21865 41916
rect 21619 41862 21621 41914
rect 21801 41862 21803 41914
rect 21557 41860 21563 41862
rect 21619 41860 21643 41862
rect 21699 41860 21723 41862
rect 21779 41860 21803 41862
rect 21859 41860 21865 41862
rect 21557 41840 21865 41860
rect 22112 41834 22140 43658
rect 22204 42226 22232 43726
rect 22296 42786 22324 44134
rect 22388 43858 22416 44134
rect 22376 43852 22428 43858
rect 22376 43794 22428 43800
rect 22468 43172 22520 43178
rect 22468 43114 22520 43120
rect 22296 42758 22416 42786
rect 22480 42770 22508 43114
rect 22572 43110 22600 44474
rect 22836 44464 22888 44470
rect 22836 44406 22888 44412
rect 22744 44328 22796 44334
rect 22744 44270 22796 44276
rect 22756 43790 22784 44270
rect 22744 43784 22796 43790
rect 22744 43726 22796 43732
rect 22848 43466 22876 44406
rect 23020 44328 23072 44334
rect 23020 44270 23072 44276
rect 22928 43784 22980 43790
rect 22928 43726 22980 43732
rect 22756 43438 22876 43466
rect 22560 43104 22612 43110
rect 22560 43046 22612 43052
rect 22652 43104 22704 43110
rect 22652 43046 22704 43052
rect 22572 42906 22600 43046
rect 22560 42900 22612 42906
rect 22560 42842 22612 42848
rect 22192 42220 22244 42226
rect 22192 42162 22244 42168
rect 22192 42016 22244 42022
rect 22192 41958 22244 41964
rect 22020 41806 22140 41834
rect 22020 41546 22048 41806
rect 22100 41676 22152 41682
rect 22100 41618 22152 41624
rect 22008 41540 22060 41546
rect 22008 41482 22060 41488
rect 21916 40928 21968 40934
rect 21916 40870 21968 40876
rect 21557 40828 21865 40848
rect 21557 40826 21563 40828
rect 21619 40826 21643 40828
rect 21699 40826 21723 40828
rect 21779 40826 21803 40828
rect 21859 40826 21865 40828
rect 21619 40774 21621 40826
rect 21801 40774 21803 40826
rect 21557 40772 21563 40774
rect 21619 40772 21643 40774
rect 21699 40772 21723 40774
rect 21779 40772 21803 40774
rect 21859 40772 21865 40774
rect 21557 40752 21865 40772
rect 21456 40112 21508 40118
rect 21456 40054 21508 40060
rect 21364 39024 21416 39030
rect 21364 38966 21416 38972
rect 21364 37732 21416 37738
rect 21364 37674 21416 37680
rect 21376 36854 21404 37674
rect 21468 37448 21496 40054
rect 21928 39982 21956 40870
rect 22112 40746 22140 41618
rect 22020 40718 22140 40746
rect 22020 40594 22048 40718
rect 22100 40656 22152 40662
rect 22100 40598 22152 40604
rect 22008 40588 22060 40594
rect 22008 40530 22060 40536
rect 22020 40390 22048 40530
rect 22008 40384 22060 40390
rect 22008 40326 22060 40332
rect 21916 39976 21968 39982
rect 21916 39918 21968 39924
rect 22008 39840 22060 39846
rect 22008 39782 22060 39788
rect 21557 39740 21865 39760
rect 21557 39738 21563 39740
rect 21619 39738 21643 39740
rect 21699 39738 21723 39740
rect 21779 39738 21803 39740
rect 21859 39738 21865 39740
rect 21619 39686 21621 39738
rect 21801 39686 21803 39738
rect 21557 39684 21563 39686
rect 21619 39684 21643 39686
rect 21699 39684 21723 39686
rect 21779 39684 21803 39686
rect 21859 39684 21865 39686
rect 21557 39664 21865 39684
rect 22020 38758 22048 39782
rect 22008 38752 22060 38758
rect 22008 38694 22060 38700
rect 21557 38652 21865 38672
rect 21557 38650 21563 38652
rect 21619 38650 21643 38652
rect 21699 38650 21723 38652
rect 21779 38650 21803 38652
rect 21859 38650 21865 38652
rect 21619 38598 21621 38650
rect 21801 38598 21803 38650
rect 21557 38596 21563 38598
rect 21619 38596 21643 38598
rect 21699 38596 21723 38598
rect 21779 38596 21803 38598
rect 21859 38596 21865 38598
rect 21557 38576 21865 38596
rect 22008 38548 22060 38554
rect 22008 38490 22060 38496
rect 21916 37868 21968 37874
rect 21916 37810 21968 37816
rect 21557 37564 21865 37584
rect 21557 37562 21563 37564
rect 21619 37562 21643 37564
rect 21699 37562 21723 37564
rect 21779 37562 21803 37564
rect 21859 37562 21865 37564
rect 21619 37510 21621 37562
rect 21801 37510 21803 37562
rect 21557 37508 21563 37510
rect 21619 37508 21643 37510
rect 21699 37508 21723 37510
rect 21779 37508 21803 37510
rect 21859 37508 21865 37510
rect 21557 37488 21865 37508
rect 21928 37466 21956 37810
rect 21916 37460 21968 37466
rect 21468 37420 21864 37448
rect 21364 36848 21416 36854
rect 21364 36790 21416 36796
rect 21364 36712 21416 36718
rect 21364 36654 21416 36660
rect 21272 36644 21324 36650
rect 21272 36586 21324 36592
rect 21180 36168 21232 36174
rect 21180 36110 21232 36116
rect 21192 35630 21220 36110
rect 21284 35834 21312 36586
rect 21376 36242 21404 36654
rect 21836 36650 21864 37420
rect 21916 37402 21968 37408
rect 21928 36922 21956 37402
rect 21916 36916 21968 36922
rect 21916 36858 21968 36864
rect 21456 36644 21508 36650
rect 21456 36586 21508 36592
rect 21824 36644 21876 36650
rect 21824 36586 21876 36592
rect 21468 36378 21496 36586
rect 21557 36476 21865 36496
rect 21557 36474 21563 36476
rect 21619 36474 21643 36476
rect 21699 36474 21723 36476
rect 21779 36474 21803 36476
rect 21859 36474 21865 36476
rect 21619 36422 21621 36474
rect 21801 36422 21803 36474
rect 21557 36420 21563 36422
rect 21619 36420 21643 36422
rect 21699 36420 21723 36422
rect 21779 36420 21803 36422
rect 21859 36420 21865 36422
rect 21557 36400 21865 36420
rect 21456 36372 21508 36378
rect 21456 36314 21508 36320
rect 21364 36236 21416 36242
rect 21364 36178 21416 36184
rect 21456 36236 21508 36242
rect 21456 36178 21508 36184
rect 21272 35828 21324 35834
rect 21272 35770 21324 35776
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21192 33318 21220 35566
rect 21180 33312 21232 33318
rect 21180 33254 21232 33260
rect 21272 33040 21324 33046
rect 21272 32982 21324 32988
rect 21284 32502 21312 32982
rect 21272 32496 21324 32502
rect 21272 32438 21324 32444
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21180 31884 21232 31890
rect 21180 31826 21232 31832
rect 21192 31754 21220 31826
rect 21180 31748 21232 31754
rect 21180 31690 21232 31696
rect 21180 30864 21232 30870
rect 21180 30806 21232 30812
rect 21192 29850 21220 30806
rect 21284 30190 21312 32302
rect 21376 30870 21404 36178
rect 21468 35630 21496 36178
rect 22020 36106 22048 38490
rect 22112 38418 22140 40598
rect 22204 40594 22232 41958
rect 22284 41608 22336 41614
rect 22284 41550 22336 41556
rect 22296 41070 22324 41550
rect 22284 41064 22336 41070
rect 22284 41006 22336 41012
rect 22284 40928 22336 40934
rect 22284 40870 22336 40876
rect 22296 40594 22324 40870
rect 22192 40588 22244 40594
rect 22192 40530 22244 40536
rect 22284 40588 22336 40594
rect 22284 40530 22336 40536
rect 22284 40384 22336 40390
rect 22284 40326 22336 40332
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 22100 38412 22152 38418
rect 22100 38354 22152 38360
rect 22100 38208 22152 38214
rect 22100 38150 22152 38156
rect 22112 37806 22140 38150
rect 22204 37874 22232 39918
rect 22296 39098 22324 40326
rect 22388 39506 22416 42758
rect 22468 42764 22520 42770
rect 22468 42706 22520 42712
rect 22664 42702 22692 43046
rect 22652 42696 22704 42702
rect 22652 42638 22704 42644
rect 22756 42566 22784 43438
rect 22744 42560 22796 42566
rect 22744 42502 22796 42508
rect 22940 42226 22968 43726
rect 23032 42362 23060 44270
rect 23124 43858 23152 44882
rect 23112 43852 23164 43858
rect 23112 43794 23164 43800
rect 23124 42770 23152 43794
rect 23308 43790 23336 45358
rect 23388 45076 23440 45082
rect 23388 45018 23440 45024
rect 23296 43784 23348 43790
rect 23296 43726 23348 43732
rect 23204 43648 23256 43654
rect 23204 43590 23256 43596
rect 23112 42764 23164 42770
rect 23112 42706 23164 42712
rect 23112 42560 23164 42566
rect 23112 42502 23164 42508
rect 23020 42356 23072 42362
rect 23020 42298 23072 42304
rect 22836 42220 22888 42226
rect 22836 42162 22888 42168
rect 22928 42220 22980 42226
rect 22928 42162 22980 42168
rect 22560 42016 22612 42022
rect 22560 41958 22612 41964
rect 22468 41064 22520 41070
rect 22468 41006 22520 41012
rect 22480 40730 22508 41006
rect 22468 40724 22520 40730
rect 22468 40666 22520 40672
rect 22468 40588 22520 40594
rect 22468 40530 22520 40536
rect 22480 39642 22508 40530
rect 22572 40050 22600 41958
rect 22744 41472 22796 41478
rect 22744 41414 22796 41420
rect 22652 40724 22704 40730
rect 22652 40666 22704 40672
rect 22560 40044 22612 40050
rect 22560 39986 22612 39992
rect 22560 39840 22612 39846
rect 22560 39782 22612 39788
rect 22468 39636 22520 39642
rect 22468 39578 22520 39584
rect 22572 39506 22600 39782
rect 22664 39642 22692 40666
rect 22652 39636 22704 39642
rect 22652 39578 22704 39584
rect 22376 39500 22428 39506
rect 22376 39442 22428 39448
rect 22560 39500 22612 39506
rect 22560 39442 22612 39448
rect 22560 39364 22612 39370
rect 22560 39306 22612 39312
rect 22468 39296 22520 39302
rect 22388 39244 22468 39250
rect 22388 39238 22520 39244
rect 22388 39222 22508 39238
rect 22284 39092 22336 39098
rect 22284 39034 22336 39040
rect 22388 38894 22416 39222
rect 22376 38888 22428 38894
rect 22376 38830 22428 38836
rect 22284 38752 22336 38758
rect 22284 38694 22336 38700
rect 22192 37868 22244 37874
rect 22192 37810 22244 37816
rect 22100 37800 22152 37806
rect 22100 37742 22152 37748
rect 22192 37460 22244 37466
rect 22192 37402 22244 37408
rect 22100 37324 22152 37330
rect 22100 37266 22152 37272
rect 22112 36922 22140 37266
rect 22100 36916 22152 36922
rect 22100 36858 22152 36864
rect 22112 36310 22140 36858
rect 22204 36786 22232 37402
rect 22192 36780 22244 36786
rect 22192 36722 22244 36728
rect 22192 36576 22244 36582
rect 22192 36518 22244 36524
rect 22100 36304 22152 36310
rect 22100 36246 22152 36252
rect 22008 36100 22060 36106
rect 22008 36042 22060 36048
rect 21548 35828 21600 35834
rect 21548 35770 21600 35776
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 21468 33658 21496 35566
rect 21560 35562 21588 35770
rect 22204 35630 22232 36518
rect 22296 36310 22324 38694
rect 22388 37194 22416 38830
rect 22468 38004 22520 38010
rect 22468 37946 22520 37952
rect 22480 37466 22508 37946
rect 22468 37460 22520 37466
rect 22468 37402 22520 37408
rect 22376 37188 22428 37194
rect 22376 37130 22428 37136
rect 22572 36786 22600 39306
rect 22560 36780 22612 36786
rect 22560 36722 22612 36728
rect 22664 36718 22692 39578
rect 22756 39506 22784 41414
rect 22848 39846 22876 42162
rect 22940 39914 22968 42162
rect 23124 42158 23152 42502
rect 23112 42152 23164 42158
rect 23112 42094 23164 42100
rect 23216 41414 23244 43590
rect 23400 42786 23428 45018
rect 23492 45014 23520 45494
rect 23480 45008 23532 45014
rect 23480 44950 23532 44956
rect 23492 43314 23520 44950
rect 23676 44334 23704 46310
rect 23768 45490 23796 46582
rect 23756 45484 23808 45490
rect 23756 45426 23808 45432
rect 23768 44878 23796 45426
rect 23756 44872 23808 44878
rect 23756 44814 23808 44820
rect 23768 44538 23796 44814
rect 23756 44532 23808 44538
rect 23756 44474 23808 44480
rect 23664 44328 23716 44334
rect 23664 44270 23716 44276
rect 23480 43308 23532 43314
rect 23480 43250 23532 43256
rect 23756 43308 23808 43314
rect 23756 43250 23808 43256
rect 23492 42906 23520 43250
rect 23480 42900 23532 42906
rect 23480 42842 23532 42848
rect 23308 42758 23428 42786
rect 23768 42770 23796 43250
rect 23756 42764 23808 42770
rect 23308 42158 23336 42758
rect 23756 42706 23808 42712
rect 23572 42628 23624 42634
rect 23572 42570 23624 42576
rect 23388 42288 23440 42294
rect 23388 42230 23440 42236
rect 23296 42152 23348 42158
rect 23296 42094 23348 42100
rect 23308 41750 23336 42094
rect 23400 42022 23428 42230
rect 23388 42016 23440 42022
rect 23388 41958 23440 41964
rect 23296 41744 23348 41750
rect 23296 41686 23348 41692
rect 23480 41676 23532 41682
rect 23480 41618 23532 41624
rect 23388 41540 23440 41546
rect 23388 41482 23440 41488
rect 23124 41386 23244 41414
rect 23020 41132 23072 41138
rect 23020 41074 23072 41080
rect 22928 39908 22980 39914
rect 22928 39850 22980 39856
rect 22836 39840 22888 39846
rect 22836 39782 22888 39788
rect 22744 39500 22796 39506
rect 22744 39442 22796 39448
rect 23032 39302 23060 41074
rect 23124 41070 23152 41386
rect 23112 41064 23164 41070
rect 23112 41006 23164 41012
rect 23400 41018 23428 41482
rect 23492 41274 23520 41618
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23480 41064 23532 41070
rect 23400 41012 23480 41018
rect 23400 41006 23532 41012
rect 23400 40990 23520 41006
rect 23112 40588 23164 40594
rect 23112 40530 23164 40536
rect 23124 40186 23152 40530
rect 23204 40520 23256 40526
rect 23204 40462 23256 40468
rect 23112 40180 23164 40186
rect 23112 40122 23164 40128
rect 23112 39976 23164 39982
rect 23112 39918 23164 39924
rect 23124 39370 23152 39918
rect 23216 39438 23244 40462
rect 23296 40384 23348 40390
rect 23296 40326 23348 40332
rect 23308 39982 23336 40326
rect 23296 39976 23348 39982
rect 23296 39918 23348 39924
rect 23204 39432 23256 39438
rect 23204 39374 23256 39380
rect 23112 39364 23164 39370
rect 23112 39306 23164 39312
rect 23020 39296 23072 39302
rect 23020 39238 23072 39244
rect 23204 38956 23256 38962
rect 23204 38898 23256 38904
rect 23112 38888 23164 38894
rect 23112 38830 23164 38836
rect 23124 38554 23152 38830
rect 23112 38548 23164 38554
rect 23112 38490 23164 38496
rect 22744 38480 22796 38486
rect 22744 38422 22796 38428
rect 22756 37126 22784 38422
rect 23020 38004 23072 38010
rect 23020 37946 23072 37952
rect 23032 37262 23060 37946
rect 23124 37806 23152 38490
rect 23216 37874 23244 38898
rect 23308 38894 23336 39918
rect 23400 39574 23428 40990
rect 23480 40656 23532 40662
rect 23480 40598 23532 40604
rect 23492 39574 23520 40598
rect 23584 40118 23612 42570
rect 23664 42016 23716 42022
rect 23664 41958 23716 41964
rect 23572 40112 23624 40118
rect 23572 40054 23624 40060
rect 23388 39568 23440 39574
rect 23388 39510 23440 39516
rect 23480 39568 23532 39574
rect 23480 39510 23532 39516
rect 23584 39250 23612 40054
rect 23676 39982 23704 41958
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23664 39500 23716 39506
rect 23664 39442 23716 39448
rect 23492 39222 23612 39250
rect 23388 39092 23440 39098
rect 23388 39034 23440 39040
rect 23400 38962 23428 39034
rect 23492 38962 23520 39222
rect 23388 38956 23440 38962
rect 23388 38898 23440 38904
rect 23480 38956 23532 38962
rect 23480 38898 23532 38904
rect 23296 38888 23348 38894
rect 23296 38830 23348 38836
rect 23204 37868 23256 37874
rect 23204 37810 23256 37816
rect 23112 37800 23164 37806
rect 23112 37742 23164 37748
rect 23308 37398 23336 38830
rect 23492 37806 23520 38898
rect 23572 38888 23624 38894
rect 23572 38830 23624 38836
rect 23676 38842 23704 39442
rect 23860 38978 23888 47126
rect 24504 46510 24532 47398
rect 24780 47258 24808 48146
rect 24872 48074 24900 48160
rect 31300 48146 31352 48152
rect 24860 48068 24912 48074
rect 24860 48010 24912 48016
rect 26709 47900 27017 47920
rect 26709 47898 26715 47900
rect 26771 47898 26795 47900
rect 26851 47898 26875 47900
rect 26931 47898 26955 47900
rect 27011 47898 27017 47900
rect 26771 47846 26773 47898
rect 26953 47846 26955 47898
rect 26709 47844 26715 47846
rect 26771 47844 26795 47846
rect 26851 47844 26875 47846
rect 26931 47844 26955 47846
rect 27011 47844 27017 47846
rect 26709 47824 27017 47844
rect 31312 47258 31340 48146
rect 24768 47252 24820 47258
rect 24768 47194 24820 47200
rect 31300 47252 31352 47258
rect 31300 47194 31352 47200
rect 30656 47116 30708 47122
rect 30656 47058 30708 47064
rect 30668 46918 30696 47058
rect 30656 46912 30708 46918
rect 30656 46854 30708 46860
rect 26709 46812 27017 46832
rect 26709 46810 26715 46812
rect 26771 46810 26795 46812
rect 26851 46810 26875 46812
rect 26931 46810 26955 46812
rect 27011 46810 27017 46812
rect 26771 46758 26773 46810
rect 26953 46758 26955 46810
rect 26709 46756 26715 46758
rect 26771 46756 26795 46758
rect 26851 46756 26875 46758
rect 26931 46756 26955 46758
rect 27011 46756 27017 46758
rect 26709 46736 27017 46756
rect 24216 46504 24268 46510
rect 24216 46446 24268 46452
rect 24492 46504 24544 46510
rect 24544 46464 24624 46492
rect 24492 46446 24544 46452
rect 24032 46028 24084 46034
rect 24032 45970 24084 45976
rect 24124 46028 24176 46034
rect 24124 45970 24176 45976
rect 23940 45280 23992 45286
rect 23940 45222 23992 45228
rect 23952 43110 23980 45222
rect 24044 44742 24072 45970
rect 24136 45082 24164 45970
rect 24228 45898 24256 46446
rect 24308 46368 24360 46374
rect 24308 46310 24360 46316
rect 24216 45892 24268 45898
rect 24216 45834 24268 45840
rect 24320 45830 24348 46310
rect 24308 45824 24360 45830
rect 24308 45766 24360 45772
rect 24400 45824 24452 45830
rect 24400 45766 24452 45772
rect 24124 45076 24176 45082
rect 24124 45018 24176 45024
rect 24216 44872 24268 44878
rect 24216 44814 24268 44820
rect 24032 44736 24084 44742
rect 24032 44678 24084 44684
rect 23940 43104 23992 43110
rect 23940 43046 23992 43052
rect 24044 42294 24072 44678
rect 24124 44532 24176 44538
rect 24124 44474 24176 44480
rect 24032 42288 24084 42294
rect 24032 42230 24084 42236
rect 23940 42084 23992 42090
rect 23940 42026 23992 42032
rect 23952 41818 23980 42026
rect 23940 41812 23992 41818
rect 23940 41754 23992 41760
rect 23940 40044 23992 40050
rect 23940 39986 23992 39992
rect 23952 39642 23980 39986
rect 23940 39636 23992 39642
rect 23940 39578 23992 39584
rect 23860 38950 24072 38978
rect 23584 38214 23612 38830
rect 23676 38814 23980 38842
rect 23664 38752 23716 38758
rect 23664 38694 23716 38700
rect 23848 38752 23900 38758
rect 23848 38694 23900 38700
rect 23676 38486 23704 38694
rect 23860 38486 23888 38694
rect 23664 38480 23716 38486
rect 23664 38422 23716 38428
rect 23848 38480 23900 38486
rect 23848 38422 23900 38428
rect 23572 38208 23624 38214
rect 23572 38150 23624 38156
rect 23848 38208 23900 38214
rect 23848 38150 23900 38156
rect 23480 37800 23532 37806
rect 23480 37742 23532 37748
rect 23584 37738 23612 38150
rect 23664 37800 23716 37806
rect 23664 37742 23716 37748
rect 23572 37732 23624 37738
rect 23572 37674 23624 37680
rect 23296 37392 23348 37398
rect 23296 37334 23348 37340
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 22928 37188 22980 37194
rect 22928 37130 22980 37136
rect 22744 37120 22796 37126
rect 22744 37062 22796 37068
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22560 36644 22612 36650
rect 22560 36586 22612 36592
rect 22284 36304 22336 36310
rect 22284 36246 22336 36252
rect 22192 35624 22244 35630
rect 22192 35566 22244 35572
rect 21548 35556 21600 35562
rect 21548 35498 21600 35504
rect 22192 35488 22244 35494
rect 22192 35430 22244 35436
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 21557 35388 21865 35408
rect 21557 35386 21563 35388
rect 21619 35386 21643 35388
rect 21699 35386 21723 35388
rect 21779 35386 21803 35388
rect 21859 35386 21865 35388
rect 21619 35334 21621 35386
rect 21801 35334 21803 35386
rect 21557 35332 21563 35334
rect 21619 35332 21643 35334
rect 21699 35332 21723 35334
rect 21779 35332 21803 35334
rect 21859 35332 21865 35334
rect 21557 35312 21865 35332
rect 21824 35148 21876 35154
rect 21824 35090 21876 35096
rect 22008 35148 22060 35154
rect 22008 35090 22060 35096
rect 21836 34388 21864 35090
rect 22020 34406 22048 35090
rect 22008 34400 22060 34406
rect 21836 34360 21956 34388
rect 21557 34300 21865 34320
rect 21557 34298 21563 34300
rect 21619 34298 21643 34300
rect 21699 34298 21723 34300
rect 21779 34298 21803 34300
rect 21859 34298 21865 34300
rect 21619 34246 21621 34298
rect 21801 34246 21803 34298
rect 21557 34244 21563 34246
rect 21619 34244 21643 34246
rect 21699 34244 21723 34246
rect 21779 34244 21803 34246
rect 21859 34244 21865 34246
rect 21557 34224 21865 34244
rect 21928 34082 21956 34360
rect 22008 34342 22060 34348
rect 21836 34054 21956 34082
rect 21456 33652 21508 33658
rect 21456 33594 21508 33600
rect 21836 33454 21864 34054
rect 21916 33992 21968 33998
rect 22020 33980 22048 34342
rect 21968 33952 22048 33980
rect 21916 33934 21968 33940
rect 21916 33856 21968 33862
rect 21916 33798 21968 33804
rect 21928 33522 21956 33798
rect 21916 33516 21968 33522
rect 21916 33458 21968 33464
rect 21824 33448 21876 33454
rect 21824 33390 21876 33396
rect 21456 33312 21508 33318
rect 21456 33254 21508 33260
rect 21916 33312 21968 33318
rect 21916 33254 21968 33260
rect 21364 30864 21416 30870
rect 21364 30806 21416 30812
rect 21272 30184 21324 30190
rect 21272 30126 21324 30132
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 21284 29714 21312 30126
rect 21272 29708 21324 29714
rect 21272 29650 21324 29656
rect 21088 29504 21140 29510
rect 21088 29446 21140 29452
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21192 29306 21220 29446
rect 21180 29300 21232 29306
rect 21180 29242 21232 29248
rect 21284 28626 21312 29650
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21180 28008 21232 28014
rect 21180 27950 21232 27956
rect 21272 28008 21324 28014
rect 21272 27950 21324 27956
rect 21192 27674 21220 27950
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 21284 27130 21312 27950
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21468 26858 21496 33254
rect 21557 33212 21865 33232
rect 21557 33210 21563 33212
rect 21619 33210 21643 33212
rect 21699 33210 21723 33212
rect 21779 33210 21803 33212
rect 21859 33210 21865 33212
rect 21619 33158 21621 33210
rect 21801 33158 21803 33210
rect 21557 33156 21563 33158
rect 21619 33156 21643 33158
rect 21699 33156 21723 33158
rect 21779 33156 21803 33158
rect 21859 33156 21865 33158
rect 21557 33136 21865 33156
rect 21928 32774 21956 33254
rect 22204 32978 22232 35430
rect 22388 35154 22416 35430
rect 22468 35284 22520 35290
rect 22468 35226 22520 35232
rect 22376 35148 22428 35154
rect 22376 35090 22428 35096
rect 22480 35086 22508 35226
rect 22468 35080 22520 35086
rect 22468 35022 22520 35028
rect 22376 35012 22428 35018
rect 22376 34954 22428 34960
rect 22388 34066 22416 34954
rect 22376 34060 22428 34066
rect 22376 34002 22428 34008
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22296 33114 22324 33934
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 22192 32972 22244 32978
rect 22192 32914 22244 32920
rect 21916 32768 21968 32774
rect 21916 32710 21968 32716
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 22112 32570 22140 32710
rect 22204 32570 22232 32914
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22192 32564 22244 32570
rect 22192 32506 22244 32512
rect 21916 32360 21968 32366
rect 21968 32308 22232 32314
rect 21916 32302 22232 32308
rect 21928 32286 22232 32302
rect 22008 32224 22060 32230
rect 22008 32166 22060 32172
rect 21557 32124 21865 32144
rect 21557 32122 21563 32124
rect 21619 32122 21643 32124
rect 21699 32122 21723 32124
rect 21779 32122 21803 32124
rect 21859 32122 21865 32124
rect 21619 32070 21621 32122
rect 21801 32070 21803 32122
rect 21557 32068 21563 32070
rect 21619 32068 21643 32070
rect 21699 32068 21723 32070
rect 21779 32068 21803 32070
rect 21859 32068 21865 32070
rect 21557 32048 21865 32068
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 21928 31754 21956 31962
rect 22020 31890 22048 32166
rect 22008 31884 22060 31890
rect 22060 31844 22140 31872
rect 22008 31826 22060 31832
rect 21916 31748 21968 31754
rect 21916 31690 21968 31696
rect 22008 31748 22060 31754
rect 22008 31690 22060 31696
rect 21640 31476 21692 31482
rect 21640 31418 21692 31424
rect 21652 31210 21680 31418
rect 21640 31204 21692 31210
rect 21640 31146 21692 31152
rect 21557 31036 21865 31056
rect 21557 31034 21563 31036
rect 21619 31034 21643 31036
rect 21699 31034 21723 31036
rect 21779 31034 21803 31036
rect 21859 31034 21865 31036
rect 21619 30982 21621 31034
rect 21801 30982 21803 31034
rect 21557 30980 21563 30982
rect 21619 30980 21643 30982
rect 21699 30980 21723 30982
rect 21779 30980 21803 30982
rect 21859 30980 21865 30982
rect 21557 30960 21865 30980
rect 21824 30796 21876 30802
rect 21824 30738 21876 30744
rect 21836 30190 21864 30738
rect 21928 30666 21956 31690
rect 22020 31278 22048 31690
rect 22008 31272 22060 31278
rect 22008 31214 22060 31220
rect 21916 30660 21968 30666
rect 21916 30602 21968 30608
rect 21824 30184 21876 30190
rect 21824 30126 21876 30132
rect 21557 29948 21865 29968
rect 21557 29946 21563 29948
rect 21619 29946 21643 29948
rect 21699 29946 21723 29948
rect 21779 29946 21803 29948
rect 21859 29946 21865 29948
rect 21619 29894 21621 29946
rect 21801 29894 21803 29946
rect 21557 29892 21563 29894
rect 21619 29892 21643 29894
rect 21699 29892 21723 29894
rect 21779 29892 21803 29894
rect 21859 29892 21865 29894
rect 21557 29872 21865 29892
rect 22020 29102 22048 31214
rect 22112 30734 22140 31844
rect 22204 30734 22232 32286
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22296 31278 22324 32166
rect 22284 31272 22336 31278
rect 22284 31214 22336 31220
rect 22284 31136 22336 31142
rect 22284 31078 22336 31084
rect 22296 30802 22324 31078
rect 22284 30796 22336 30802
rect 22284 30738 22336 30744
rect 22100 30728 22152 30734
rect 22100 30670 22152 30676
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 22112 29646 22140 30670
rect 22204 30258 22232 30670
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22204 29714 22232 30194
rect 22192 29708 22244 29714
rect 22192 29650 22244 29656
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 22284 29640 22336 29646
rect 22388 29628 22416 33798
rect 22480 32978 22508 35022
rect 22572 33114 22600 36586
rect 22756 36038 22784 37062
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22664 34066 22692 34342
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 22560 33108 22612 33114
rect 22560 33050 22612 33056
rect 22468 32972 22520 32978
rect 22468 32914 22520 32920
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22572 30938 22600 31826
rect 22664 31142 22692 34002
rect 22756 33454 22784 35974
rect 22836 35556 22888 35562
rect 22836 35498 22888 35504
rect 22848 33862 22876 35498
rect 22836 33856 22888 33862
rect 22836 33798 22888 33804
rect 22744 33448 22796 33454
rect 22744 33390 22796 33396
rect 22744 33108 22796 33114
rect 22744 33050 22796 33056
rect 22756 31754 22784 33050
rect 22756 31726 22876 31754
rect 22744 31272 22796 31278
rect 22744 31214 22796 31220
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22468 30184 22520 30190
rect 22468 30126 22520 30132
rect 22480 29714 22508 30126
rect 22756 29782 22784 31214
rect 22744 29776 22796 29782
rect 22664 29736 22744 29764
rect 22468 29708 22520 29714
rect 22468 29650 22520 29656
rect 22336 29600 22416 29628
rect 22284 29582 22336 29588
rect 22100 29300 22152 29306
rect 22100 29242 22152 29248
rect 22008 29096 22060 29102
rect 22008 29038 22060 29044
rect 21557 28860 21865 28880
rect 21557 28858 21563 28860
rect 21619 28858 21643 28860
rect 21699 28858 21723 28860
rect 21779 28858 21803 28860
rect 21859 28858 21865 28860
rect 21619 28806 21621 28858
rect 21801 28806 21803 28858
rect 21557 28804 21563 28806
rect 21619 28804 21643 28806
rect 21699 28804 21723 28806
rect 21779 28804 21803 28806
rect 21859 28804 21865 28806
rect 21557 28784 21865 28804
rect 22112 28694 22140 29242
rect 22192 29096 22244 29102
rect 22192 29038 22244 29044
rect 22204 28694 22232 29038
rect 22100 28688 22152 28694
rect 22100 28630 22152 28636
rect 22192 28688 22244 28694
rect 22192 28630 22244 28636
rect 22008 28008 22060 28014
rect 22008 27950 22060 27956
rect 21557 27772 21865 27792
rect 21557 27770 21563 27772
rect 21619 27770 21643 27772
rect 21699 27770 21723 27772
rect 21779 27770 21803 27772
rect 21859 27770 21865 27772
rect 21619 27718 21621 27770
rect 21801 27718 21803 27770
rect 21557 27716 21563 27718
rect 21619 27716 21643 27718
rect 21699 27716 21723 27718
rect 21779 27716 21803 27718
rect 21859 27716 21865 27718
rect 21557 27696 21865 27716
rect 22020 26994 22048 27950
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 20904 26852 20956 26858
rect 20904 26794 20956 26800
rect 21456 26852 21508 26858
rect 21456 26794 21508 26800
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 20720 26512 20772 26518
rect 20720 26454 20772 26460
rect 20444 26444 20496 26450
rect 20444 26386 20496 26392
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 20076 25764 20128 25770
rect 20076 25706 20128 25712
rect 20088 24818 20116 25706
rect 20180 25702 20208 26318
rect 20260 25832 20312 25838
rect 20260 25774 20312 25780
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19628 23662 19656 23802
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19524 22772 19576 22778
rect 19628 22760 19656 23598
rect 19996 23322 20024 24142
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 19708 22772 19760 22778
rect 19628 22732 19708 22760
rect 19524 22714 19576 22720
rect 19708 22714 19760 22720
rect 19444 22630 19564 22658
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19260 22234 19380 22250
rect 19248 22228 19380 22234
rect 19300 22222 19380 22228
rect 19248 22170 19300 22176
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 19352 21418 19380 22102
rect 19444 21690 19472 22374
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19156 20800 19208 20806
rect 19156 20742 19208 20748
rect 19168 19718 19196 20742
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19260 18970 19288 19382
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19352 18630 19380 18838
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 19168 16946 19196 18090
rect 19260 18068 19288 18362
rect 19340 18216 19392 18222
rect 19444 18204 19472 18770
rect 19392 18176 19472 18204
rect 19340 18158 19392 18164
rect 19260 18040 19380 18068
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19076 16918 19196 16946
rect 19076 16658 19104 16918
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 19168 16250 19196 16458
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19260 15858 19288 17274
rect 19352 16114 19380 18040
rect 19536 17882 19564 22630
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19628 19922 19656 21966
rect 19720 21486 19748 22714
rect 19800 22500 19852 22506
rect 19800 22442 19852 22448
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19812 20806 19840 22442
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19904 21894 19932 22034
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19996 21622 20024 23258
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 20088 20942 20116 23530
rect 20168 21412 20220 21418
rect 20168 21354 20220 21360
rect 20180 20942 20208 21354
rect 20272 21350 20300 25774
rect 20456 24818 20484 26386
rect 20548 25702 20576 26386
rect 20732 26314 20944 26330
rect 20720 26308 20944 26314
rect 20772 26302 20944 26308
rect 20720 26250 20772 26256
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 20456 23254 20484 23666
rect 20444 23248 20496 23254
rect 20444 23190 20496 23196
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19720 19122 19748 20402
rect 20180 20398 20208 20878
rect 20272 20602 20300 21286
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 19628 19094 19748 19122
rect 19628 18766 19656 19094
rect 19800 18964 19852 18970
rect 19720 18924 19800 18952
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19628 18154 19656 18702
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19076 15830 19288 15858
rect 19076 15586 19104 15830
rect 18972 15564 19024 15570
rect 19076 15558 19196 15586
rect 19536 15570 19564 17002
rect 18972 15506 19024 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 18984 14958 19012 15370
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 19076 14804 19104 15438
rect 18984 14776 19104 14804
rect 18984 14090 19012 14776
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 19076 14278 19104 14554
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18984 14062 19104 14090
rect 18892 12406 19012 12434
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 18156 7002 18184 7958
rect 18248 7546 18276 8502
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18144 6860 18196 6866
rect 18064 6820 18144 6848
rect 18144 6802 18196 6808
rect 17972 5766 18092 5794
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17972 5166 18000 5578
rect 18064 5574 18092 5766
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 18064 5098 18092 5170
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17972 4282 18000 4490
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17776 2576 17828 2582
rect 17972 2564 18000 4218
rect 18064 4146 18092 5034
rect 18156 4282 18184 5102
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18248 4214 18276 5306
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18340 4146 18368 8434
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18524 7818 18552 8230
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 7478 18460 7686
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18524 6798 18552 7278
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18616 6202 18644 11766
rect 18708 10810 18736 12038
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18708 10130 18736 10406
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18432 6174 18644 6202
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18248 3194 18276 4014
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18340 2990 18368 3470
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 17828 2536 18000 2564
rect 17776 2518 17828 2524
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 17316 1760 17368 1766
rect 17316 1702 17368 1708
rect 17316 1488 17368 1494
rect 17316 1430 17368 1436
rect 17184 1244 17264 1272
rect 17132 1226 17184 1232
rect 17236 882 17264 1244
rect 17224 876 17276 882
rect 17224 818 17276 824
rect 17328 814 17356 1430
rect 17420 1426 17448 2450
rect 17972 2446 18000 2536
rect 18064 2514 18092 2858
rect 18432 2774 18460 6174
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18616 5302 18644 5646
rect 18708 5370 18736 7346
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18604 5296 18656 5302
rect 18604 5238 18656 5244
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18616 4758 18644 5102
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18512 3460 18564 3466
rect 18512 3402 18564 3408
rect 18524 2990 18552 3402
rect 18708 2990 18736 3674
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18432 2746 18552 2774
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18064 2378 18092 2450
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18432 1766 18460 2450
rect 18420 1760 18472 1766
rect 18420 1702 18472 1708
rect 17408 1420 17460 1426
rect 17408 1362 17460 1368
rect 17500 1420 17552 1426
rect 17500 1362 17552 1368
rect 17512 1018 17540 1362
rect 18524 1018 18552 2746
rect 18708 2514 18736 2926
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18616 1902 18644 2246
rect 18800 2106 18828 8570
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18892 5030 18920 7822
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18892 4690 18920 4966
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18880 2372 18932 2378
rect 18880 2314 18932 2320
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18604 1896 18656 1902
rect 18604 1838 18656 1844
rect 18892 1562 18920 2314
rect 18880 1556 18932 1562
rect 18880 1498 18932 1504
rect 18984 1018 19012 12406
rect 19076 11354 19104 14062
rect 19168 12782 19196 15558
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19260 15094 19288 15506
rect 19628 15162 19656 17070
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19260 14618 19288 15030
rect 19352 14958 19380 15030
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19352 13258 19380 14894
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 14346 19564 14418
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19536 13938 19564 14282
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19536 13394 19564 13874
rect 19628 13530 19656 14826
rect 19720 14074 19748 18924
rect 19800 18906 19852 18912
rect 20180 18834 20208 20334
rect 20364 19446 20392 21830
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20272 18714 20300 19246
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 19996 18686 20300 18714
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19812 18222 19840 18566
rect 19904 18358 19932 18566
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19812 17610 19840 18158
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19904 16658 19932 18022
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19812 14362 19840 15438
rect 19904 15144 19932 16050
rect 19996 15366 20024 18686
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19984 15156 20036 15162
rect 19904 15116 19984 15144
rect 19984 15098 20036 15104
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19904 14482 19932 14758
rect 19996 14618 20024 14758
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19812 14334 19932 14362
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19720 13394 19748 14010
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19708 13388 19760 13394
rect 19708 13330 19760 13336
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 12306 19196 12718
rect 19352 12322 19380 13194
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19432 12436 19484 12442
rect 19536 12424 19564 12786
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19484 12396 19564 12424
rect 19432 12378 19484 12384
rect 19156 12300 19208 12306
rect 19352 12294 19564 12322
rect 19156 12242 19208 12248
rect 19168 11694 19196 12242
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19352 11762 19380 12174
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19444 11694 19472 12174
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19168 10198 19196 11086
rect 19340 10600 19392 10606
rect 19444 10588 19472 11630
rect 19392 10560 19472 10588
rect 19340 10542 19392 10548
rect 19444 10266 19472 10560
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19168 8838 19196 10134
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 8498 19196 8774
rect 19352 8650 19380 9590
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19260 8622 19380 8650
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19168 7886 19196 8434
rect 19260 8294 19288 8622
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19076 5914 19104 6122
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19076 4758 19104 5850
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19076 3534 19104 4558
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19076 1494 19104 2926
rect 19064 1488 19116 1494
rect 19064 1430 19116 1436
rect 19168 1358 19196 7822
rect 19352 6866 19380 8502
rect 19444 8004 19472 9318
rect 19536 8634 19564 12294
rect 19628 11898 19656 12718
rect 19708 12708 19760 12714
rect 19708 12650 19760 12656
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19628 10674 19656 11834
rect 19720 11830 19748 12650
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19812 11558 19840 12242
rect 19904 12220 19932 14334
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19996 12986 20024 13738
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20088 12374 20116 17818
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 20180 16046 20208 17750
rect 20364 17746 20392 18770
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20272 16794 20300 17546
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20272 15586 20300 16730
rect 20180 15558 20300 15586
rect 20180 15162 20208 15558
rect 20260 15428 20312 15434
rect 20260 15370 20312 15376
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 20180 13462 20208 14826
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 19984 12232 20036 12238
rect 19904 12192 19984 12220
rect 19984 12174 20036 12180
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19812 10810 19840 11494
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19800 10532 19852 10538
rect 19800 10474 19852 10480
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19524 8016 19576 8022
rect 19444 7976 19524 8004
rect 19524 7958 19576 7964
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19260 4826 19288 6190
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19260 4214 19288 4762
rect 19248 4208 19300 4214
rect 19248 4150 19300 4156
rect 19260 3738 19288 4150
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 2514 19288 3538
rect 19352 3194 19380 3946
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19260 2106 19288 2450
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19156 1352 19208 1358
rect 19156 1294 19208 1300
rect 19444 1018 19472 7278
rect 19720 6866 19748 7890
rect 19812 7750 19840 10474
rect 19904 10130 19932 12038
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 11286 20024 11494
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 20088 10674 20116 12310
rect 20180 12170 20208 13398
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19904 7546 19932 9454
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 19628 4826 19656 5714
rect 19812 5166 19840 6190
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19812 4622 19840 5102
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19720 3602 19748 4014
rect 19812 3602 19840 4558
rect 19904 4486 19932 6258
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19720 2854 19748 3538
rect 19812 3058 19840 3538
rect 19904 3534 19932 4422
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19812 2582 19840 2994
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 19524 2508 19576 2514
rect 19576 2468 19656 2496
rect 19524 2450 19576 2456
rect 19628 2378 19656 2468
rect 19616 2372 19668 2378
rect 19616 2314 19668 2320
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 19812 1494 19840 2246
rect 19800 1488 19852 1494
rect 19800 1430 19852 1436
rect 17500 1012 17552 1018
rect 17500 954 17552 960
rect 18512 1012 18564 1018
rect 18512 954 18564 960
rect 18972 1012 19024 1018
rect 18972 954 19024 960
rect 19432 1012 19484 1018
rect 19432 954 19484 960
rect 20088 950 20116 8842
rect 20180 7274 20208 12106
rect 20272 9382 20300 15370
rect 20364 15094 20392 17682
rect 20456 17134 20484 18362
rect 20548 18358 20576 25638
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20640 23662 20668 24210
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20640 23186 20668 23598
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20536 18080 20588 18086
rect 20732 18034 20760 25366
rect 20824 24750 20852 26182
rect 20916 25294 20944 26302
rect 21100 26246 21128 26726
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21008 25362 21036 26182
rect 21468 26042 21496 26794
rect 21557 26684 21865 26704
rect 21557 26682 21563 26684
rect 21619 26682 21643 26684
rect 21699 26682 21723 26684
rect 21779 26682 21803 26684
rect 21859 26682 21865 26684
rect 21619 26630 21621 26682
rect 21801 26630 21803 26682
rect 21557 26628 21563 26630
rect 21619 26628 21643 26630
rect 21699 26628 21723 26630
rect 21779 26628 21803 26630
rect 21859 26628 21865 26630
rect 21557 26608 21865 26628
rect 22008 26308 22060 26314
rect 22008 26250 22060 26256
rect 21456 26036 21508 26042
rect 21284 25996 21456 26024
rect 21284 25498 21312 25996
rect 21456 25978 21508 25984
rect 21916 25764 21968 25770
rect 21916 25706 21968 25712
rect 21557 25596 21865 25616
rect 21557 25594 21563 25596
rect 21619 25594 21643 25596
rect 21699 25594 21723 25596
rect 21779 25594 21803 25596
rect 21859 25594 21865 25596
rect 21619 25542 21621 25594
rect 21801 25542 21803 25594
rect 21557 25540 21563 25542
rect 21619 25540 21643 25542
rect 21699 25540 21723 25542
rect 21779 25540 21803 25542
rect 21859 25540 21865 25542
rect 21557 25520 21865 25540
rect 21272 25492 21324 25498
rect 21272 25434 21324 25440
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20904 24880 20956 24886
rect 20904 24822 20956 24828
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20812 24336 20864 24342
rect 20812 24278 20864 24284
rect 20824 23662 20852 24278
rect 20916 24274 20944 24822
rect 21088 24676 21140 24682
rect 21088 24618 21140 24624
rect 21100 24274 21128 24618
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20916 23322 20944 24210
rect 21284 23882 21312 25434
rect 21364 24676 21416 24682
rect 21364 24618 21416 24624
rect 21376 24410 21404 24618
rect 21928 24614 21956 25706
rect 22020 25702 22048 26250
rect 22112 25974 22140 27474
rect 22100 25968 22152 25974
rect 22100 25910 22152 25916
rect 22204 25906 22232 28630
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22296 26450 22324 28358
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22296 25838 22324 26386
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21557 24508 21865 24528
rect 21557 24506 21563 24508
rect 21619 24506 21643 24508
rect 21699 24506 21723 24508
rect 21779 24506 21803 24508
rect 21859 24506 21865 24508
rect 21619 24454 21621 24506
rect 21801 24454 21803 24506
rect 21557 24452 21563 24454
rect 21619 24452 21643 24454
rect 21699 24452 21723 24454
rect 21779 24452 21803 24454
rect 21859 24452 21865 24454
rect 21557 24432 21865 24452
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21284 23854 21496 23882
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20916 21434 20944 22918
rect 21008 22234 21036 23666
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21284 22506 21312 23122
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20824 21406 20944 21434
rect 20824 21350 20852 21406
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 20262 20852 21286
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20916 20398 20944 20946
rect 21100 20398 21128 21490
rect 21376 21078 21404 22714
rect 21468 21690 21496 23854
rect 21560 23798 21588 24006
rect 21548 23792 21600 23798
rect 21548 23734 21600 23740
rect 21557 23420 21865 23440
rect 21557 23418 21563 23420
rect 21619 23418 21643 23420
rect 21699 23418 21723 23420
rect 21779 23418 21803 23420
rect 21859 23418 21865 23420
rect 21619 23366 21621 23418
rect 21801 23366 21803 23418
rect 21557 23364 21563 23366
rect 21619 23364 21643 23366
rect 21699 23364 21723 23366
rect 21779 23364 21803 23366
rect 21859 23364 21865 23366
rect 21557 23344 21865 23364
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21836 23050 21864 23122
rect 21824 23044 21876 23050
rect 21824 22986 21876 22992
rect 21557 22332 21865 22352
rect 21557 22330 21563 22332
rect 21619 22330 21643 22332
rect 21699 22330 21723 22332
rect 21779 22330 21803 22332
rect 21859 22330 21865 22332
rect 21619 22278 21621 22330
rect 21801 22278 21803 22330
rect 21557 22276 21563 22278
rect 21619 22276 21643 22278
rect 21699 22276 21723 22278
rect 21779 22276 21803 22278
rect 21859 22276 21865 22278
rect 21557 22256 21865 22276
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21557 21244 21865 21264
rect 21557 21242 21563 21244
rect 21619 21242 21643 21244
rect 21699 21242 21723 21244
rect 21779 21242 21803 21244
rect 21859 21242 21865 21244
rect 21619 21190 21621 21242
rect 21801 21190 21803 21242
rect 21557 21188 21563 21190
rect 21619 21188 21643 21190
rect 21699 21188 21723 21190
rect 21779 21188 21803 21190
rect 21859 21188 21865 21190
rect 21557 21168 21865 21188
rect 21928 21146 21956 24550
rect 22112 23662 22140 25162
rect 22296 24954 22324 25298
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22008 23180 22060 23186
rect 22008 23122 22060 23128
rect 22020 23050 22048 23122
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22112 22778 22140 23598
rect 22296 23526 22324 24074
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22388 22930 22416 29600
rect 22480 28422 22508 29650
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22572 28626 22600 29446
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 22468 28416 22520 28422
rect 22468 28358 22520 28364
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22572 26586 22600 26862
rect 22560 26580 22612 26586
rect 22560 26522 22612 26528
rect 22664 26518 22692 29736
rect 22744 29718 22796 29724
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22756 27470 22784 28358
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22744 26920 22796 26926
rect 22744 26862 22796 26868
rect 22652 26512 22704 26518
rect 22572 26460 22652 26466
rect 22572 26454 22704 26460
rect 22572 26438 22692 26454
rect 22572 26042 22600 26438
rect 22652 26308 22704 26314
rect 22652 26250 22704 26256
rect 22560 26036 22612 26042
rect 22560 25978 22612 25984
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 22480 24698 22508 24890
rect 22480 24670 22600 24698
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22480 23594 22508 24550
rect 22572 24274 22600 24670
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22468 23588 22520 23594
rect 22468 23530 22520 23536
rect 22560 23588 22612 23594
rect 22560 23530 22612 23536
rect 22572 23322 22600 23530
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22388 22902 22508 22930
rect 22100 22772 22152 22778
rect 22100 22714 22152 22720
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22112 22234 22140 22714
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22112 22098 22140 22170
rect 22100 22092 22152 22098
rect 22100 22034 22152 22040
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21364 20528 21416 20534
rect 21364 20470 21416 20476
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20916 20040 20944 20334
rect 20824 20012 20944 20040
rect 20824 18766 20852 20012
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20916 18970 20944 19858
rect 21100 19496 21128 20334
rect 21180 20324 21232 20330
rect 21180 20266 21232 20272
rect 21192 20058 21220 20266
rect 21376 20262 21404 20470
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21180 19508 21232 19514
rect 21100 19468 21180 19496
rect 21180 19450 21232 19456
rect 21284 19310 21312 20198
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20824 18290 20852 18702
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20536 18022 20588 18028
rect 20548 17678 20576 18022
rect 20640 18006 20760 18034
rect 20640 17882 20668 18006
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20824 17218 20852 17614
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20732 17190 20852 17218
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20456 12186 20484 17070
rect 20548 16658 20576 17138
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 13734 20576 15302
rect 20640 15162 20668 15506
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20732 13394 20760 17190
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20824 16726 20852 17070
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20824 16250 20852 16662
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20824 15026 20852 16186
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20824 14550 20852 14962
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20916 14074 20944 18702
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 20996 17536 21048 17542
rect 21100 17524 21128 18022
rect 21376 17678 21404 19654
rect 21468 18902 21496 20538
rect 22112 20466 22140 21490
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21557 20156 21865 20176
rect 21557 20154 21563 20156
rect 21619 20154 21643 20156
rect 21699 20154 21723 20156
rect 21779 20154 21803 20156
rect 21859 20154 21865 20156
rect 21619 20102 21621 20154
rect 21801 20102 21803 20154
rect 21557 20100 21563 20102
rect 21619 20100 21643 20102
rect 21699 20100 21723 20102
rect 21779 20100 21803 20102
rect 21859 20100 21865 20102
rect 21557 20080 21865 20100
rect 21557 19068 21865 19088
rect 21557 19066 21563 19068
rect 21619 19066 21643 19068
rect 21699 19066 21723 19068
rect 21779 19066 21803 19068
rect 21859 19066 21865 19068
rect 21619 19014 21621 19066
rect 21801 19014 21803 19066
rect 21557 19012 21563 19014
rect 21619 19012 21643 19014
rect 21699 19012 21723 19014
rect 21779 19012 21803 19014
rect 21859 19012 21865 19014
rect 21557 18992 21865 19012
rect 21928 18970 21956 20334
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 22020 19514 22048 20266
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21456 18896 21508 18902
rect 21456 18838 21508 18844
rect 22020 18834 22048 19450
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 21557 17980 21865 18000
rect 21557 17978 21563 17980
rect 21619 17978 21643 17980
rect 21699 17978 21723 17980
rect 21779 17978 21803 17980
rect 21859 17978 21865 17980
rect 21619 17926 21621 17978
rect 21801 17926 21803 17978
rect 21557 17924 21563 17926
rect 21619 17924 21643 17926
rect 21699 17924 21723 17926
rect 21779 17924 21803 17926
rect 21859 17924 21865 17926
rect 21557 17904 21865 17924
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21048 17496 21128 17524
rect 20996 17478 21048 17484
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20732 13190 20760 13330
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20824 12782 20852 12854
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12434 20760 12582
rect 20732 12406 20944 12434
rect 20812 12232 20864 12238
rect 20456 12158 20760 12186
rect 20812 12174 20864 12180
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 10810 20484 12038
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20640 11762 20668 11834
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20640 11354 20668 11698
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20364 10266 20392 10474
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20272 6390 20300 8910
rect 20456 8838 20484 9454
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7410 20392 7822
rect 20548 7818 20576 8978
rect 20732 8294 20760 12158
rect 20824 10198 20852 12174
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20180 4690 20208 6054
rect 20456 5710 20484 7278
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20456 4758 20484 5646
rect 20732 5302 20760 6598
rect 20720 5296 20772 5302
rect 20720 5238 20772 5244
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 20732 4690 20760 4966
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20272 1902 20300 2450
rect 20260 1896 20312 1902
rect 20260 1838 20312 1844
rect 20272 1358 20300 1838
rect 20732 1834 20760 3470
rect 20720 1828 20772 1834
rect 20720 1770 20772 1776
rect 20260 1352 20312 1358
rect 20260 1294 20312 1300
rect 20824 1018 20852 7210
rect 20916 6322 20944 12406
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21008 8634 21036 10746
rect 21100 10742 21128 17496
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 15570 21220 17478
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 13530 21220 14214
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21284 12918 21312 14010
rect 21376 13462 21404 17614
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21468 16250 21496 17002
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21557 16892 21865 16912
rect 21557 16890 21563 16892
rect 21619 16890 21643 16892
rect 21699 16890 21723 16892
rect 21779 16890 21803 16892
rect 21859 16890 21865 16892
rect 21619 16838 21621 16890
rect 21801 16838 21803 16890
rect 21557 16836 21563 16838
rect 21619 16836 21643 16838
rect 21699 16836 21723 16838
rect 21779 16836 21803 16838
rect 21859 16836 21865 16838
rect 21557 16816 21865 16836
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21557 15804 21865 15824
rect 21557 15802 21563 15804
rect 21619 15802 21643 15804
rect 21699 15802 21723 15804
rect 21779 15802 21803 15804
rect 21859 15802 21865 15804
rect 21619 15750 21621 15802
rect 21801 15750 21803 15802
rect 21557 15748 21563 15750
rect 21619 15748 21643 15750
rect 21699 15748 21723 15750
rect 21779 15748 21803 15750
rect 21859 15748 21865 15750
rect 21557 15728 21865 15748
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21468 14074 21496 14826
rect 21928 14770 21956 16934
rect 22020 16658 22048 18090
rect 22112 17542 22140 19926
rect 22204 18086 22232 21626
rect 22296 19922 22324 21966
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22296 19310 22324 19858
rect 22388 19310 22416 22714
rect 22480 21690 22508 22902
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22480 20602 22508 20878
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22296 17746 22324 19246
rect 22480 18970 22508 19858
rect 22572 19174 22600 20946
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22664 18222 22692 26250
rect 22756 26042 22784 26862
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 22756 24818 22784 25842
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22756 23186 22784 24006
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22848 22094 22876 31726
rect 22940 28082 22968 37130
rect 23032 36718 23060 37198
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 23388 37120 23440 37126
rect 23388 37062 23440 37068
rect 23112 36780 23164 36786
rect 23112 36722 23164 36728
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 23032 36038 23060 36654
rect 23020 36032 23072 36038
rect 23020 35974 23072 35980
rect 23020 33924 23072 33930
rect 23020 33866 23072 33872
rect 23032 32230 23060 33866
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 23124 31754 23152 36722
rect 23216 36650 23244 37062
rect 23296 36916 23348 36922
rect 23296 36858 23348 36864
rect 23204 36644 23256 36650
rect 23204 36586 23256 36592
rect 23308 36242 23336 36858
rect 23296 36236 23348 36242
rect 23296 36178 23348 36184
rect 23204 35760 23256 35766
rect 23204 35702 23256 35708
rect 23216 33522 23244 35702
rect 23400 33998 23428 37062
rect 23676 36922 23704 37742
rect 23756 37732 23808 37738
rect 23756 37674 23808 37680
rect 23664 36916 23716 36922
rect 23664 36858 23716 36864
rect 23768 36786 23796 37674
rect 23860 37398 23888 38150
rect 23848 37392 23900 37398
rect 23848 37334 23900 37340
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23848 36712 23900 36718
rect 23848 36654 23900 36660
rect 23572 36304 23624 36310
rect 23572 36246 23624 36252
rect 23584 35290 23612 36246
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35630 23704 35974
rect 23860 35698 23888 36654
rect 23952 36242 23980 38814
rect 23940 36236 23992 36242
rect 23940 36178 23992 36184
rect 23848 35692 23900 35698
rect 23848 35634 23900 35640
rect 23664 35624 23716 35630
rect 23664 35566 23716 35572
rect 23848 35556 23900 35562
rect 23848 35498 23900 35504
rect 23572 35284 23624 35290
rect 23572 35226 23624 35232
rect 23664 34128 23716 34134
rect 23664 34070 23716 34076
rect 23388 33992 23440 33998
rect 23388 33934 23440 33940
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 23204 33516 23256 33522
rect 23256 33476 23336 33504
rect 23204 33458 23256 33464
rect 23204 33380 23256 33386
rect 23204 33322 23256 33328
rect 23216 32026 23244 33322
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23308 31754 23336 33476
rect 23400 33386 23428 33798
rect 23388 33380 23440 33386
rect 23388 33322 23440 33328
rect 23676 33114 23704 34070
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23664 33108 23716 33114
rect 23664 33050 23716 33056
rect 23572 32972 23624 32978
rect 23572 32914 23624 32920
rect 23584 32570 23612 32914
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 23388 32360 23440 32366
rect 23388 32302 23440 32308
rect 23032 31726 23152 31754
rect 23216 31726 23336 31754
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 22940 22778 22968 27406
rect 23032 27062 23060 31726
rect 23112 30592 23164 30598
rect 23112 30534 23164 30540
rect 23124 30394 23152 30534
rect 23112 30388 23164 30394
rect 23112 30330 23164 30336
rect 23216 30326 23244 31726
rect 23400 31414 23428 32302
rect 23388 31408 23440 31414
rect 23388 31350 23440 31356
rect 23388 31204 23440 31210
rect 23388 31146 23440 31152
rect 23400 30734 23428 31146
rect 23492 30802 23520 32370
rect 23768 32348 23796 33254
rect 23584 32320 23796 32348
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 23296 30660 23348 30666
rect 23296 30602 23348 30608
rect 23308 30546 23336 30602
rect 23308 30518 23428 30546
rect 23204 30320 23256 30326
rect 23204 30262 23256 30268
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 23204 30048 23256 30054
rect 23204 29990 23256 29996
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 23124 27606 23152 29514
rect 23216 29102 23244 29990
rect 23308 29306 23336 30126
rect 23296 29300 23348 29306
rect 23296 29242 23348 29248
rect 23204 29096 23256 29102
rect 23204 29038 23256 29044
rect 23204 28960 23256 28966
rect 23204 28902 23256 28908
rect 23216 28694 23244 28902
rect 23204 28688 23256 28694
rect 23204 28630 23256 28636
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 23020 27056 23072 27062
rect 23020 26998 23072 27004
rect 23204 26920 23256 26926
rect 23204 26862 23256 26868
rect 23216 26518 23244 26862
rect 23204 26512 23256 26518
rect 23204 26454 23256 26460
rect 23112 26444 23164 26450
rect 23112 26386 23164 26392
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 24206 23060 26182
rect 23124 24750 23152 26386
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 23216 24886 23244 26318
rect 23308 25838 23336 29242
rect 23400 29186 23428 30518
rect 23400 29158 23520 29186
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23400 28966 23428 29038
rect 23388 28960 23440 28966
rect 23388 28902 23440 28908
rect 23492 28506 23520 29158
rect 23400 28478 23520 28506
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23204 24880 23256 24886
rect 23204 24822 23256 24828
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 23032 22250 23060 24142
rect 23124 23730 23152 24142
rect 23216 24070 23244 24210
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 23112 23588 23164 23594
rect 23216 23576 23244 24006
rect 23308 23866 23336 24890
rect 23400 24614 23428 28478
rect 23584 27520 23612 32320
rect 23756 32224 23808 32230
rect 23756 32166 23808 32172
rect 23768 30734 23796 32166
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23676 27946 23704 29990
rect 23756 28620 23808 28626
rect 23756 28562 23808 28568
rect 23664 27940 23716 27946
rect 23664 27882 23716 27888
rect 23492 27492 23612 27520
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23492 24426 23520 27492
rect 23572 27396 23624 27402
rect 23572 27338 23624 27344
rect 23584 26450 23612 27338
rect 23676 27062 23704 27882
rect 23768 27538 23796 28562
rect 23860 28082 23888 35498
rect 23952 34950 23980 36178
rect 23940 34944 23992 34950
rect 23940 34886 23992 34892
rect 23952 34678 23980 34886
rect 23940 34672 23992 34678
rect 23940 34614 23992 34620
rect 23940 32836 23992 32842
rect 23940 32778 23992 32784
rect 23952 32366 23980 32778
rect 23940 32360 23992 32366
rect 23940 32302 23992 32308
rect 23940 31680 23992 31686
rect 23940 31622 23992 31628
rect 23952 31414 23980 31622
rect 23940 31408 23992 31414
rect 23940 31350 23992 31356
rect 23940 30320 23992 30326
rect 23940 30262 23992 30268
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23664 27056 23716 27062
rect 23664 26998 23716 27004
rect 23572 26444 23624 26450
rect 23572 26386 23624 26392
rect 23584 24954 23612 26386
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23400 24398 23520 24426
rect 23400 24342 23428 24398
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23164 23548 23244 23576
rect 23112 23530 23164 23536
rect 23124 23050 23152 23530
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23112 23044 23164 23050
rect 23112 22986 23164 22992
rect 23124 22778 23152 22986
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23032 22222 23152 22250
rect 23308 22234 23336 23054
rect 23020 22160 23072 22166
rect 23020 22102 23072 22108
rect 22756 22066 22876 22094
rect 22756 19310 22784 22066
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22940 19174 22968 20810
rect 22928 19168 22980 19174
rect 22928 19110 22980 19116
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 16658 22232 16934
rect 22480 16794 22508 17274
rect 22572 16794 22600 17682
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22112 15706 22140 15982
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 21928 14742 22048 14770
rect 21557 14716 21865 14736
rect 21557 14714 21563 14716
rect 21619 14714 21643 14716
rect 21699 14714 21723 14716
rect 21779 14714 21803 14716
rect 21859 14714 21865 14716
rect 21619 14662 21621 14714
rect 21801 14662 21803 14714
rect 21557 14660 21563 14662
rect 21619 14660 21643 14662
rect 21699 14660 21723 14662
rect 21779 14660 21803 14662
rect 21859 14660 21865 14662
rect 21557 14640 21865 14660
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21652 14006 21680 14214
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 21824 13864 21876 13870
rect 21928 13818 21956 14010
rect 21876 13812 21956 13818
rect 21824 13806 21956 13812
rect 21456 13796 21508 13802
rect 21836 13790 21956 13806
rect 21456 13738 21508 13744
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21468 13190 21496 13738
rect 21557 13628 21865 13648
rect 21557 13626 21563 13628
rect 21619 13626 21643 13628
rect 21699 13626 21723 13628
rect 21779 13626 21803 13628
rect 21859 13626 21865 13628
rect 21619 13574 21621 13626
rect 21801 13574 21803 13626
rect 21557 13572 21563 13574
rect 21619 13572 21643 13574
rect 21699 13572 21723 13574
rect 21779 13572 21803 13574
rect 21859 13572 21865 13574
rect 21557 13552 21865 13572
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 21560 13190 21588 13398
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21272 12912 21324 12918
rect 21272 12854 21324 12860
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 21192 9602 21220 12582
rect 21284 11830 21312 12854
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21376 11642 21404 12174
rect 21284 11614 21404 11642
rect 21284 11218 21312 11614
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21091 9574 21220 9602
rect 21091 9194 21119 9574
rect 21091 9166 21312 9194
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21100 6730 21128 8230
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20916 1018 20944 6122
rect 21100 5778 21128 6190
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21008 5234 21036 5510
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21100 4486 21128 5714
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 21100 3466 21128 4422
rect 21192 4078 21220 9046
rect 21284 8906 21312 9166
rect 21376 9160 21404 10678
rect 21468 10130 21496 13126
rect 21836 12628 21864 13398
rect 21928 12782 21956 13790
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 21916 12640 21968 12646
rect 21836 12600 21916 12628
rect 21916 12582 21968 12588
rect 21557 12540 21865 12560
rect 21557 12538 21563 12540
rect 21619 12538 21643 12540
rect 21699 12538 21723 12540
rect 21779 12538 21803 12540
rect 21859 12538 21865 12540
rect 21619 12486 21621 12538
rect 21801 12486 21803 12538
rect 21557 12484 21563 12486
rect 21619 12484 21643 12486
rect 21699 12484 21723 12486
rect 21779 12484 21803 12486
rect 21859 12484 21865 12486
rect 21557 12464 21865 12484
rect 21916 12436 21968 12442
rect 21836 12396 21916 12424
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21560 11898 21588 12174
rect 21836 12170 21864 12396
rect 21916 12378 21968 12384
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 21557 11452 21865 11472
rect 21557 11450 21563 11452
rect 21619 11450 21643 11452
rect 21699 11450 21723 11452
rect 21779 11450 21803 11452
rect 21859 11450 21865 11452
rect 21619 11398 21621 11450
rect 21801 11398 21803 11450
rect 21557 11396 21563 11398
rect 21619 11396 21643 11398
rect 21699 11396 21723 11398
rect 21779 11396 21803 11398
rect 21859 11396 21865 11398
rect 21557 11376 21865 11396
rect 21928 10810 21956 11494
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 22020 10674 22048 14742
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22112 13394 22140 13942
rect 22296 13530 22324 15574
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22388 13394 22416 15574
rect 22480 15502 22508 15846
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22480 15366 22508 15438
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22664 14906 22692 18158
rect 22572 14878 22692 14906
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22480 14618 22508 14758
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22572 13802 22600 14878
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 13870 22692 14758
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22112 11898 22140 12242
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22204 11762 22232 12650
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22112 10554 22140 11154
rect 22020 10526 22140 10554
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 21557 10364 21865 10384
rect 21557 10362 21563 10364
rect 21619 10362 21643 10364
rect 21699 10362 21723 10364
rect 21779 10362 21803 10364
rect 21859 10362 21865 10364
rect 21619 10310 21621 10362
rect 21801 10310 21803 10362
rect 21557 10308 21563 10310
rect 21619 10308 21643 10310
rect 21699 10308 21723 10310
rect 21779 10308 21803 10310
rect 21859 10308 21865 10310
rect 21557 10288 21865 10308
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21744 9364 21772 10066
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21836 9586 21864 9862
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21928 9500 21956 10202
rect 22020 9586 22048 10526
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22112 9722 22140 9930
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22204 9654 22232 10542
rect 22296 10266 22324 13126
rect 22388 12714 22416 13330
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22480 12782 22508 13262
rect 22756 12986 22784 18770
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22848 16658 22876 18022
rect 23032 17882 23060 22102
rect 23124 21162 23152 22222
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 23124 21134 23244 21162
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 23124 20602 23152 21014
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 23124 16998 23152 18566
rect 23216 17762 23244 21134
rect 23308 21010 23336 22170
rect 23676 21894 23704 26998
rect 23768 26858 23796 27474
rect 23756 26852 23808 26858
rect 23756 26794 23808 26800
rect 23848 26444 23900 26450
rect 23848 26386 23900 26392
rect 23860 24410 23888 26386
rect 23848 24404 23900 24410
rect 23848 24346 23900 24352
rect 23952 22094 23980 30262
rect 24044 26518 24072 38950
rect 24032 26512 24084 26518
rect 24032 26454 24084 26460
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 24044 25702 24072 26318
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 24044 22794 24072 25638
rect 24136 25430 24164 44474
rect 24228 44470 24256 44814
rect 24320 44810 24348 45766
rect 24412 44946 24440 45766
rect 24400 44940 24452 44946
rect 24400 44882 24452 44888
rect 24492 44940 24544 44946
rect 24492 44882 24544 44888
rect 24308 44804 24360 44810
rect 24308 44746 24360 44752
rect 24216 44464 24268 44470
rect 24216 44406 24268 44412
rect 24216 44260 24268 44266
rect 24216 44202 24268 44208
rect 24228 43994 24256 44202
rect 24216 43988 24268 43994
rect 24216 43930 24268 43936
rect 24412 43858 24440 44882
rect 24504 44470 24532 44882
rect 24492 44464 24544 44470
rect 24492 44406 24544 44412
rect 24596 44334 24624 46464
rect 25136 46368 25188 46374
rect 25136 46310 25188 46316
rect 25688 46368 25740 46374
rect 25688 46310 25740 46316
rect 25148 46102 25176 46310
rect 25136 46096 25188 46102
rect 25136 46038 25188 46044
rect 25700 44946 25728 46310
rect 30668 46034 30696 46854
rect 30656 46028 30708 46034
rect 30656 45970 30708 45976
rect 31576 46028 31628 46034
rect 31576 45970 31628 45976
rect 26148 45960 26200 45966
rect 26148 45902 26200 45908
rect 26160 45626 26188 45902
rect 26240 45824 26292 45830
rect 26240 45766 26292 45772
rect 26252 45626 26280 45766
rect 26709 45724 27017 45744
rect 26709 45722 26715 45724
rect 26771 45722 26795 45724
rect 26851 45722 26875 45724
rect 26931 45722 26955 45724
rect 27011 45722 27017 45724
rect 26771 45670 26773 45722
rect 26953 45670 26955 45722
rect 26709 45668 26715 45670
rect 26771 45668 26795 45670
rect 26851 45668 26875 45670
rect 26931 45668 26955 45670
rect 27011 45668 27017 45670
rect 26709 45648 27017 45668
rect 26148 45620 26200 45626
rect 26148 45562 26200 45568
rect 26240 45620 26292 45626
rect 26240 45562 26292 45568
rect 26160 45490 26188 45562
rect 26148 45484 26200 45490
rect 26148 45426 26200 45432
rect 26056 45280 26108 45286
rect 26056 45222 26108 45228
rect 25688 44940 25740 44946
rect 25688 44882 25740 44888
rect 24768 44804 24820 44810
rect 24768 44746 24820 44752
rect 24584 44328 24636 44334
rect 24584 44270 24636 44276
rect 24400 43852 24452 43858
rect 24400 43794 24452 43800
rect 24676 43444 24728 43450
rect 24676 43386 24728 43392
rect 24400 43240 24452 43246
rect 24400 43182 24452 43188
rect 24216 42764 24268 42770
rect 24216 42706 24268 42712
rect 24228 42022 24256 42706
rect 24308 42560 24360 42566
rect 24308 42502 24360 42508
rect 24320 42090 24348 42502
rect 24412 42158 24440 43182
rect 24400 42152 24452 42158
rect 24400 42094 24452 42100
rect 24308 42084 24360 42090
rect 24308 42026 24360 42032
rect 24216 42016 24268 42022
rect 24216 41958 24268 41964
rect 24308 41268 24360 41274
rect 24308 41210 24360 41216
rect 24216 40996 24268 41002
rect 24216 40938 24268 40944
rect 24228 40662 24256 40938
rect 24216 40656 24268 40662
rect 24216 40598 24268 40604
rect 24228 39982 24256 40598
rect 24216 39976 24268 39982
rect 24216 39918 24268 39924
rect 24228 38554 24256 39918
rect 24320 39642 24348 41210
rect 24584 41200 24636 41206
rect 24584 41142 24636 41148
rect 24596 39982 24624 41142
rect 24584 39976 24636 39982
rect 24584 39918 24636 39924
rect 24308 39636 24360 39642
rect 24308 39578 24360 39584
rect 24400 39364 24452 39370
rect 24400 39306 24452 39312
rect 24308 38752 24360 38758
rect 24308 38694 24360 38700
rect 24216 38548 24268 38554
rect 24216 38490 24268 38496
rect 24320 34762 24348 38694
rect 24412 38214 24440 39306
rect 24584 39024 24636 39030
rect 24584 38966 24636 38972
rect 24492 38548 24544 38554
rect 24492 38490 24544 38496
rect 24400 38208 24452 38214
rect 24400 38150 24452 38156
rect 24400 37868 24452 37874
rect 24400 37810 24452 37816
rect 24412 37346 24440 37810
rect 24504 37806 24532 38490
rect 24492 37800 24544 37806
rect 24492 37742 24544 37748
rect 24504 37466 24532 37742
rect 24492 37460 24544 37466
rect 24492 37402 24544 37408
rect 24412 37330 24532 37346
rect 24412 37324 24544 37330
rect 24412 37318 24492 37324
rect 24492 37266 24544 37272
rect 24492 36100 24544 36106
rect 24228 34734 24348 34762
rect 24412 36060 24492 36088
rect 24228 30666 24256 34734
rect 24308 34672 24360 34678
rect 24308 34614 24360 34620
rect 24216 30660 24268 30666
rect 24216 30602 24268 30608
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24124 25424 24176 25430
rect 24124 25366 24176 25372
rect 24124 24676 24176 24682
rect 24228 24664 24256 30262
rect 24320 28762 24348 34614
rect 24308 28756 24360 28762
rect 24308 28698 24360 28704
rect 24320 27606 24348 28698
rect 24412 28150 24440 36060
rect 24492 36042 24544 36048
rect 24596 34134 24624 38966
rect 24584 34128 24636 34134
rect 24584 34070 24636 34076
rect 24492 33448 24544 33454
rect 24492 33390 24544 33396
rect 24504 33130 24532 33390
rect 24596 33318 24624 34070
rect 24584 33312 24636 33318
rect 24584 33254 24636 33260
rect 24504 33114 24624 33130
rect 24504 33108 24636 33114
rect 24504 33102 24584 33108
rect 24584 33050 24636 33056
rect 24492 31952 24544 31958
rect 24492 31894 24544 31900
rect 24504 31686 24532 31894
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 24596 31226 24624 33050
rect 24688 31754 24716 43386
rect 24780 40186 24808 44746
rect 24860 44736 24912 44742
rect 24860 44678 24912 44684
rect 24872 43926 24900 44678
rect 25320 44192 25372 44198
rect 25320 44134 25372 44140
rect 25872 44192 25924 44198
rect 25872 44134 25924 44140
rect 24860 43920 24912 43926
rect 24860 43862 24912 43868
rect 25228 43648 25280 43654
rect 25228 43590 25280 43596
rect 25044 42764 25096 42770
rect 25044 42706 25096 42712
rect 24952 42696 25004 42702
rect 24952 42638 25004 42644
rect 24860 41676 24912 41682
rect 24860 41618 24912 41624
rect 24872 40526 24900 41618
rect 24964 41562 24992 42638
rect 25056 42158 25084 42706
rect 25044 42152 25096 42158
rect 25044 42094 25096 42100
rect 25056 41682 25084 42094
rect 25044 41676 25096 41682
rect 25044 41618 25096 41624
rect 24964 41534 25176 41562
rect 24952 41472 25004 41478
rect 24952 41414 25004 41420
rect 25044 41472 25096 41478
rect 25044 41414 25096 41420
rect 24964 40526 24992 41414
rect 24860 40520 24912 40526
rect 24860 40462 24912 40468
rect 24952 40520 25004 40526
rect 24952 40462 25004 40468
rect 24768 40180 24820 40186
rect 24768 40122 24820 40128
rect 24872 39982 24900 40462
rect 24860 39976 24912 39982
rect 24860 39918 24912 39924
rect 24768 38956 24820 38962
rect 24768 38898 24820 38904
rect 24780 38214 24808 38898
rect 24872 38282 24900 39918
rect 24952 39568 25004 39574
rect 24952 39510 25004 39516
rect 24964 38654 24992 39510
rect 25056 38758 25084 41414
rect 25148 41138 25176 41534
rect 25136 41132 25188 41138
rect 25136 41074 25188 41080
rect 25044 38752 25096 38758
rect 25044 38694 25096 38700
rect 24964 38626 25084 38654
rect 24860 38276 24912 38282
rect 24860 38218 24912 38224
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 24872 37398 24900 38218
rect 24860 37392 24912 37398
rect 24860 37334 24912 37340
rect 24860 36848 24912 36854
rect 24860 36790 24912 36796
rect 24872 35290 24900 36790
rect 24952 36576 25004 36582
rect 24952 36518 25004 36524
rect 24964 35766 24992 36518
rect 24952 35760 25004 35766
rect 24952 35702 25004 35708
rect 24860 35284 24912 35290
rect 24860 35226 24912 35232
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 24860 34536 24912 34542
rect 24860 34478 24912 34484
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24780 33114 24808 33934
rect 24872 33454 24900 34478
rect 24860 33448 24912 33454
rect 24860 33390 24912 33396
rect 24768 33108 24820 33114
rect 24768 33050 24820 33056
rect 24872 32978 24900 33390
rect 24964 33046 24992 34886
rect 25056 33318 25084 38626
rect 25240 38536 25268 43590
rect 25332 41478 25360 44134
rect 25884 43858 25912 44134
rect 25688 43852 25740 43858
rect 25688 43794 25740 43800
rect 25872 43852 25924 43858
rect 25872 43794 25924 43800
rect 25700 42702 25728 43794
rect 25688 42696 25740 42702
rect 25688 42638 25740 42644
rect 25884 41818 25912 43794
rect 25872 41812 25924 41818
rect 25872 41754 25924 41760
rect 25412 41744 25464 41750
rect 25412 41686 25464 41692
rect 25320 41472 25372 41478
rect 25320 41414 25372 41420
rect 25320 40520 25372 40526
rect 25320 40462 25372 40468
rect 25332 39846 25360 40462
rect 25320 39840 25372 39846
rect 25320 39782 25372 39788
rect 25332 39506 25360 39782
rect 25320 39500 25372 39506
rect 25320 39442 25372 39448
rect 25332 39098 25360 39442
rect 25320 39092 25372 39098
rect 25320 39034 25372 39040
rect 25148 38508 25268 38536
rect 25148 38282 25176 38508
rect 25332 38486 25360 39034
rect 25424 39030 25452 41686
rect 25780 41676 25832 41682
rect 25780 41618 25832 41624
rect 25792 41274 25820 41618
rect 25780 41268 25832 41274
rect 25780 41210 25832 41216
rect 26068 40662 26096 45222
rect 26252 44198 26280 45562
rect 27620 45484 27672 45490
rect 27620 45426 27672 45432
rect 27528 45416 27580 45422
rect 27528 45358 27580 45364
rect 26424 44940 26476 44946
rect 26424 44882 26476 44888
rect 26332 44736 26384 44742
rect 26332 44678 26384 44684
rect 26240 44192 26292 44198
rect 26240 44134 26292 44140
rect 26344 44010 26372 44678
rect 26252 43982 26372 44010
rect 26436 43994 26464 44882
rect 26709 44636 27017 44656
rect 26709 44634 26715 44636
rect 26771 44634 26795 44636
rect 26851 44634 26875 44636
rect 26931 44634 26955 44636
rect 27011 44634 27017 44636
rect 26771 44582 26773 44634
rect 26953 44582 26955 44634
rect 26709 44580 26715 44582
rect 26771 44580 26795 44582
rect 26851 44580 26875 44582
rect 26931 44580 26955 44582
rect 27011 44580 27017 44582
rect 26709 44560 27017 44580
rect 27540 44470 27568 45358
rect 27632 44742 27660 45426
rect 27620 44736 27672 44742
rect 27620 44678 27672 44684
rect 30932 44736 30984 44742
rect 30932 44678 30984 44684
rect 27068 44464 27120 44470
rect 27068 44406 27120 44412
rect 27528 44464 27580 44470
rect 27528 44406 27580 44412
rect 26608 44260 26660 44266
rect 26608 44202 26660 44208
rect 26424 43988 26476 43994
rect 26252 43858 26280 43982
rect 26424 43930 26476 43936
rect 26240 43852 26292 43858
rect 26240 43794 26292 43800
rect 26148 43716 26200 43722
rect 26148 43658 26200 43664
rect 26160 43382 26188 43658
rect 26148 43376 26200 43382
rect 26148 43318 26200 43324
rect 26252 43178 26280 43794
rect 26332 43784 26384 43790
rect 26332 43726 26384 43732
rect 26344 43314 26372 43726
rect 26332 43308 26384 43314
rect 26332 43250 26384 43256
rect 26240 43172 26292 43178
rect 26240 43114 26292 43120
rect 26148 43104 26200 43110
rect 26148 43046 26200 43052
rect 26160 42752 26188 43046
rect 26240 42764 26292 42770
rect 26160 42724 26240 42752
rect 26240 42706 26292 42712
rect 26344 42650 26372 43250
rect 26424 43240 26476 43246
rect 26424 43182 26476 43188
rect 26436 42702 26464 43182
rect 26160 42622 26372 42650
rect 26424 42696 26476 42702
rect 26424 42638 26476 42644
rect 26160 41614 26188 42622
rect 26332 42560 26384 42566
rect 26332 42502 26384 42508
rect 26344 42362 26372 42502
rect 26332 42356 26384 42362
rect 26332 42298 26384 42304
rect 26436 42242 26464 42638
rect 26516 42560 26568 42566
rect 26516 42502 26568 42508
rect 26344 42214 26464 42242
rect 26240 42152 26292 42158
rect 26344 42140 26372 42214
rect 26292 42112 26372 42140
rect 26240 42094 26292 42100
rect 26148 41608 26200 41614
rect 26148 41550 26200 41556
rect 26160 41138 26188 41550
rect 26240 41540 26292 41546
rect 26240 41482 26292 41488
rect 26148 41132 26200 41138
rect 26148 41074 26200 41080
rect 26056 40656 26108 40662
rect 26056 40598 26108 40604
rect 25504 40588 25556 40594
rect 25504 40530 25556 40536
rect 25516 40474 25544 40530
rect 26056 40520 26108 40526
rect 25516 40446 25728 40474
rect 26160 40508 26188 41074
rect 26252 41070 26280 41482
rect 26344 41206 26372 42112
rect 26424 42130 26476 42136
rect 26424 42072 26476 42078
rect 26436 41478 26464 42072
rect 26424 41472 26476 41478
rect 26424 41414 26476 41420
rect 26332 41200 26384 41206
rect 26332 41142 26384 41148
rect 26240 41064 26292 41070
rect 26240 41006 26292 41012
rect 26332 41064 26384 41070
rect 26332 41006 26384 41012
rect 26108 40480 26188 40508
rect 26056 40462 26108 40468
rect 25412 39024 25464 39030
rect 25412 38966 25464 38972
rect 25320 38480 25372 38486
rect 25320 38422 25372 38428
rect 25228 38412 25280 38418
rect 25228 38354 25280 38360
rect 25136 38276 25188 38282
rect 25136 38218 25188 38224
rect 25240 38010 25268 38354
rect 25320 38276 25372 38282
rect 25320 38218 25372 38224
rect 25228 38004 25280 38010
rect 25228 37946 25280 37952
rect 25136 37936 25188 37942
rect 25136 37878 25188 37884
rect 25148 36038 25176 37878
rect 25332 36922 25360 38218
rect 25412 38208 25464 38214
rect 25412 38150 25464 38156
rect 25424 37806 25452 38150
rect 25412 37800 25464 37806
rect 25412 37742 25464 37748
rect 25320 36916 25372 36922
rect 25320 36858 25372 36864
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25148 35630 25176 35974
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25044 33312 25096 33318
rect 25044 33254 25096 33260
rect 24952 33040 25004 33046
rect 24952 32982 25004 32988
rect 25044 33040 25096 33046
rect 25044 32982 25096 32988
rect 24860 32972 24912 32978
rect 24780 32932 24860 32960
rect 24780 32366 24808 32932
rect 24860 32914 24912 32920
rect 24952 32904 25004 32910
rect 24952 32846 25004 32852
rect 24768 32360 24820 32366
rect 24768 32302 24820 32308
rect 24860 32292 24912 32298
rect 24964 32280 24992 32846
rect 25056 32502 25084 32982
rect 25044 32496 25096 32502
rect 25044 32438 25096 32444
rect 25148 32348 25176 35566
rect 25332 35562 25360 36858
rect 25504 36032 25556 36038
rect 25504 35974 25556 35980
rect 25320 35556 25372 35562
rect 25320 35498 25372 35504
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 25240 34678 25268 35430
rect 25412 35284 25464 35290
rect 25412 35226 25464 35232
rect 25228 34672 25280 34678
rect 25228 34614 25280 34620
rect 25240 33930 25268 34614
rect 25424 34542 25452 35226
rect 25320 34536 25372 34542
rect 25320 34478 25372 34484
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25332 34406 25360 34478
rect 25320 34400 25372 34406
rect 25320 34342 25372 34348
rect 25228 33924 25280 33930
rect 25228 33866 25280 33872
rect 25240 33522 25268 33866
rect 25228 33516 25280 33522
rect 25228 33458 25280 33464
rect 25228 33380 25280 33386
rect 25332 33368 25360 34342
rect 25424 34134 25452 34478
rect 25412 34128 25464 34134
rect 25412 34070 25464 34076
rect 25424 33862 25452 34070
rect 25412 33856 25464 33862
rect 25412 33798 25464 33804
rect 25280 33340 25360 33368
rect 25228 33322 25280 33328
rect 25412 33312 25464 33318
rect 25412 33254 25464 33260
rect 25424 32994 25452 33254
rect 25516 33114 25544 35974
rect 25596 35148 25648 35154
rect 25596 35090 25648 35096
rect 25608 34678 25636 35090
rect 25596 34672 25648 34678
rect 25596 34614 25648 34620
rect 25596 34196 25648 34202
rect 25596 34138 25648 34144
rect 25608 33590 25636 34138
rect 25596 33584 25648 33590
rect 25596 33526 25648 33532
rect 25596 33448 25648 33454
rect 25596 33390 25648 33396
rect 25504 33108 25556 33114
rect 25504 33050 25556 33056
rect 25332 32966 25452 32994
rect 25608 32978 25636 33390
rect 25596 32972 25648 32978
rect 24912 32252 24992 32280
rect 25056 32320 25176 32348
rect 25228 32360 25280 32366
rect 24860 32234 24912 32240
rect 25056 32212 25084 32320
rect 25228 32302 25280 32308
rect 24964 32184 25084 32212
rect 24964 32008 24992 32184
rect 24964 31980 25176 32008
rect 24688 31726 24808 31754
rect 24596 31198 24716 31226
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24492 30796 24544 30802
rect 24492 30738 24544 30744
rect 24504 28506 24532 30738
rect 24596 29034 24624 31078
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24504 28478 24624 28506
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24504 28014 24532 28358
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 24400 27668 24452 27674
rect 24400 27610 24452 27616
rect 24308 27600 24360 27606
rect 24308 27542 24360 27548
rect 24320 27402 24348 27542
rect 24308 27396 24360 27402
rect 24308 27338 24360 27344
rect 24412 27062 24440 27610
rect 24400 27056 24452 27062
rect 24400 26998 24452 27004
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24492 26784 24544 26790
rect 24492 26726 24544 26732
rect 24412 26518 24440 26726
rect 24400 26512 24452 26518
rect 24400 26454 24452 26460
rect 24308 26308 24360 26314
rect 24308 26250 24360 26256
rect 24176 24636 24256 24664
rect 24124 24618 24176 24624
rect 24136 24410 24164 24618
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24320 24342 24348 26250
rect 24504 25498 24532 26726
rect 24596 26314 24624 28478
rect 24688 28218 24716 31198
rect 24780 30326 24808 31726
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24952 31476 25004 31482
rect 24952 31418 25004 31424
rect 24872 30870 24900 31418
rect 24964 31346 24992 31418
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24860 30864 24912 30870
rect 24860 30806 24912 30812
rect 24768 30320 24820 30326
rect 24768 30262 24820 30268
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 24872 29034 24900 29650
rect 24860 29028 24912 29034
rect 24860 28970 24912 28976
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24688 26450 24716 28154
rect 24780 27606 24808 28630
rect 24872 28082 24900 28970
rect 24964 28694 24992 31282
rect 25044 31204 25096 31210
rect 25044 31146 25096 31152
rect 25056 28966 25084 31146
rect 25044 28960 25096 28966
rect 25044 28902 25096 28908
rect 24952 28688 25004 28694
rect 24952 28630 25004 28636
rect 25056 28626 25084 28902
rect 25044 28620 25096 28626
rect 25044 28562 25096 28568
rect 24952 28416 25004 28422
rect 24952 28358 25004 28364
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24964 27656 24992 28358
rect 24872 27628 24992 27656
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24780 27130 24808 27542
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 24584 26308 24636 26314
rect 24584 26250 24636 26256
rect 24676 25832 24728 25838
rect 24676 25774 24728 25780
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24400 25356 24452 25362
rect 24400 25298 24452 25304
rect 24412 24954 24440 25298
rect 24400 24948 24452 24954
rect 24400 24890 24452 24896
rect 24492 24948 24544 24954
rect 24492 24890 24544 24896
rect 24308 24336 24360 24342
rect 24308 24278 24360 24284
rect 24216 24200 24268 24206
rect 24216 24142 24268 24148
rect 24044 22766 24164 22794
rect 23952 22066 24072 22094
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23572 21412 23624 21418
rect 23572 21354 23624 21360
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 23388 20460 23440 20466
rect 23584 20448 23612 21354
rect 23676 21078 23704 21422
rect 23860 21146 23888 21966
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 23952 21690 23980 21830
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 23440 20420 23612 20448
rect 23388 20402 23440 20408
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23308 19310 23336 19654
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23492 18834 23520 19314
rect 23584 18970 23612 20420
rect 23860 20398 23888 21082
rect 24044 21010 24072 22066
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24136 20890 24164 22766
rect 24044 20862 24164 20890
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23848 20392 23900 20398
rect 23848 20334 23900 20340
rect 23676 20058 23704 20334
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23860 19378 23888 20334
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23664 18692 23716 18698
rect 23664 18634 23716 18640
rect 23676 18426 23704 18634
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23400 17882 23428 18158
rect 23768 18154 23796 19246
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23216 17734 23428 17762
rect 23400 17490 23428 17734
rect 23308 17462 23428 17490
rect 23204 17060 23256 17066
rect 23204 17002 23256 17008
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23124 16658 23152 16934
rect 22836 16652 22888 16658
rect 23112 16652 23164 16658
rect 22836 16594 22888 16600
rect 23032 16612 23112 16640
rect 22848 16454 22876 16594
rect 22928 16516 22980 16522
rect 22928 16458 22980 16464
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22940 15162 22968 16458
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22848 13870 22876 14962
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 13870 22968 14214
rect 23032 14074 23060 16612
rect 23112 16594 23164 16600
rect 23216 16590 23244 17002
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23124 14958 23152 15506
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23308 14278 23336 17462
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23492 16250 23520 17070
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23492 14550 23520 15914
rect 23584 15706 23612 16594
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23676 15502 23704 18022
rect 23768 16794 23796 18090
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23860 16658 23888 17138
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23676 15094 23704 15438
rect 23768 15162 23796 15914
rect 23952 15570 23980 17478
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23952 15366 23980 15506
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23664 15088 23716 15094
rect 24044 15042 24072 20862
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 23664 15030 23716 15036
rect 23768 15014 24072 15042
rect 23768 14958 23796 15014
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23400 14074 23428 14418
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22480 10606 22508 11630
rect 22572 10606 22600 12854
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22388 10130 22416 10406
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22296 9674 22324 10066
rect 22192 9648 22244 9654
rect 22296 9646 22416 9674
rect 22192 9590 22244 9596
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 21928 9472 21972 9500
rect 21944 9466 21972 9472
rect 21944 9438 22094 9466
rect 21744 9336 21956 9364
rect 21557 9276 21865 9296
rect 21557 9274 21563 9276
rect 21619 9274 21643 9276
rect 21699 9274 21723 9276
rect 21779 9274 21803 9276
rect 21859 9274 21865 9276
rect 21619 9222 21621 9274
rect 21801 9222 21803 9274
rect 21557 9220 21563 9222
rect 21619 9220 21643 9222
rect 21699 9220 21723 9222
rect 21779 9220 21803 9222
rect 21859 9220 21865 9222
rect 21557 9200 21865 9220
rect 21376 9132 21588 9160
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 21456 8560 21508 8566
rect 21456 8502 21508 8508
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21284 8022 21312 8230
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21284 6458 21312 7754
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 21376 3040 21404 8298
rect 21468 5710 21496 8502
rect 21560 8276 21588 9132
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21652 8634 21680 8774
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21836 8430 21864 8774
rect 21928 8566 21956 9336
rect 22066 9330 22094 9438
rect 22020 9302 22094 9330
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21560 8248 21956 8276
rect 21557 8188 21865 8208
rect 21557 8186 21563 8188
rect 21619 8186 21643 8188
rect 21699 8186 21723 8188
rect 21779 8186 21803 8188
rect 21859 8186 21865 8188
rect 21619 8134 21621 8186
rect 21801 8134 21803 8186
rect 21557 8132 21563 8134
rect 21619 8132 21643 8134
rect 21699 8132 21723 8134
rect 21779 8132 21803 8134
rect 21859 8132 21865 8134
rect 21557 8112 21865 8132
rect 21557 7100 21865 7120
rect 21557 7098 21563 7100
rect 21619 7098 21643 7100
rect 21699 7098 21723 7100
rect 21779 7098 21803 7100
rect 21859 7098 21865 7100
rect 21619 7046 21621 7098
rect 21801 7046 21803 7098
rect 21557 7044 21563 7046
rect 21619 7044 21643 7046
rect 21699 7044 21723 7046
rect 21779 7044 21803 7046
rect 21859 7044 21865 7046
rect 21557 7024 21865 7044
rect 21928 6458 21956 8248
rect 22020 7818 22048 9302
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22112 8362 22140 9114
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 22112 7546 22140 7890
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 22020 7002 22048 7210
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22112 6866 22140 7482
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 21557 6012 21865 6032
rect 21557 6010 21563 6012
rect 21619 6010 21643 6012
rect 21699 6010 21723 6012
rect 21779 6010 21803 6012
rect 21859 6010 21865 6012
rect 21619 5958 21621 6010
rect 21801 5958 21803 6010
rect 21557 5956 21563 5958
rect 21619 5956 21643 5958
rect 21699 5956 21723 5958
rect 21779 5956 21803 5958
rect 21859 5956 21865 5958
rect 21557 5936 21865 5956
rect 21928 5914 21956 6258
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21824 5092 21876 5098
rect 21876 5052 21956 5080
rect 21824 5034 21876 5040
rect 21557 4924 21865 4944
rect 21557 4922 21563 4924
rect 21619 4922 21643 4924
rect 21699 4922 21723 4924
rect 21779 4922 21803 4924
rect 21859 4922 21865 4924
rect 21619 4870 21621 4922
rect 21801 4870 21803 4922
rect 21557 4868 21563 4870
rect 21619 4868 21643 4870
rect 21699 4868 21723 4870
rect 21779 4868 21803 4870
rect 21859 4868 21865 4870
rect 21557 4848 21865 4868
rect 21928 4826 21956 5052
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 22020 4196 22048 6190
rect 22204 4758 22232 9590
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22296 7886 22324 8910
rect 22388 8838 22416 9646
rect 22572 9518 22600 10542
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22664 9178 22692 12718
rect 22756 12306 22784 12786
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22848 11694 22876 13806
rect 22940 13190 22968 13806
rect 23124 13530 23152 13806
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23492 13444 23520 14486
rect 23768 13530 23796 14894
rect 24044 14618 24072 14894
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23664 13456 23716 13462
rect 23492 13416 23664 13444
rect 23664 13398 23716 13404
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 22928 12708 22980 12714
rect 22928 12650 22980 12656
rect 22940 12238 22968 12650
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 22940 11626 22968 12174
rect 22928 11620 22980 11626
rect 22928 11562 22980 11568
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22756 10538 22784 11086
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 22744 10532 22796 10538
rect 22744 10474 22796 10480
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22296 6866 22324 7822
rect 22388 7342 22416 8366
rect 22480 7954 22508 8842
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22296 6322 22324 6802
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21928 4168 22048 4196
rect 21557 3836 21865 3856
rect 21557 3834 21563 3836
rect 21619 3834 21643 3836
rect 21699 3834 21723 3836
rect 21779 3834 21803 3836
rect 21859 3834 21865 3836
rect 21619 3782 21621 3834
rect 21801 3782 21803 3834
rect 21557 3780 21563 3782
rect 21619 3780 21643 3782
rect 21699 3780 21723 3782
rect 21779 3780 21803 3782
rect 21859 3780 21865 3782
rect 21557 3760 21865 3780
rect 21928 3534 21956 4168
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 21376 3012 21496 3040
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21376 2446 21404 2858
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 21468 1562 21496 3012
rect 21928 2922 21956 3470
rect 22204 3126 22232 4558
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 21916 2916 21968 2922
rect 21916 2858 21968 2864
rect 22112 2802 22140 2926
rect 22020 2774 22140 2802
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 21557 2748 21865 2768
rect 21557 2746 21563 2748
rect 21619 2746 21643 2748
rect 21699 2746 21723 2748
rect 21779 2746 21803 2748
rect 21859 2746 21865 2748
rect 21619 2694 21621 2746
rect 21801 2694 21803 2746
rect 21557 2692 21563 2694
rect 21619 2692 21643 2694
rect 21699 2692 21723 2694
rect 21779 2692 21803 2694
rect 21859 2692 21865 2694
rect 21557 2672 21865 2692
rect 22020 2650 22048 2774
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22204 2582 22232 2790
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 21557 1660 21865 1680
rect 21557 1658 21563 1660
rect 21619 1658 21643 1660
rect 21699 1658 21723 1660
rect 21779 1658 21803 1660
rect 21859 1658 21865 1660
rect 21619 1606 21621 1658
rect 21801 1606 21803 1658
rect 21557 1604 21563 1606
rect 21619 1604 21643 1606
rect 21699 1604 21723 1606
rect 21779 1604 21803 1606
rect 21859 1604 21865 1606
rect 21557 1584 21865 1604
rect 21456 1556 21508 1562
rect 21456 1498 21508 1504
rect 22296 1018 22324 5646
rect 22388 5234 22416 7278
rect 22480 6730 22508 7890
rect 22572 7800 22600 8978
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22664 8090 22692 8298
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22652 7812 22704 7818
rect 22572 7772 22652 7800
rect 22652 7754 22704 7760
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22572 6338 22600 7414
rect 22664 6866 22692 7754
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22480 6310 22600 6338
rect 22480 6186 22508 6310
rect 22560 6248 22612 6254
rect 22664 6236 22692 6802
rect 22612 6208 22692 6236
rect 22560 6190 22612 6196
rect 22468 6180 22520 6186
rect 22468 6122 22520 6128
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22388 4282 22416 5170
rect 22572 4690 22600 6190
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22388 2990 22416 4218
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22652 1828 22704 1834
rect 22652 1770 22704 1776
rect 22664 1358 22692 1770
rect 22652 1352 22704 1358
rect 22652 1294 22704 1300
rect 22756 1018 22784 10474
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22848 7886 22876 8978
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22940 7002 22968 7686
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22848 5234 22876 6258
rect 22940 6254 22968 6666
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 22940 5234 22968 6190
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22848 4622 22876 5170
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22848 2922 22876 3538
rect 22836 2916 22888 2922
rect 22836 2858 22888 2864
rect 22848 2106 22876 2858
rect 22836 2100 22888 2106
rect 22836 2042 22888 2048
rect 22848 1426 22876 2042
rect 22836 1420 22888 1426
rect 22836 1362 22888 1368
rect 20812 1012 20864 1018
rect 20812 954 20864 960
rect 20904 1012 20956 1018
rect 20904 954 20956 960
rect 22284 1012 22336 1018
rect 22284 954 22336 960
rect 22744 1012 22796 1018
rect 22744 954 22796 960
rect 23032 950 23060 9998
rect 23124 7546 23152 10542
rect 23216 10266 23244 11154
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 2106 23152 6394
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 23216 950 23244 8774
rect 23308 6984 23336 12378
rect 23676 12306 23704 12922
rect 24136 12434 24164 20742
rect 24228 17882 24256 24142
rect 24504 23866 24532 24890
rect 24596 24750 24624 25638
rect 24584 24744 24636 24750
rect 24584 24686 24636 24692
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24492 23860 24544 23866
rect 24492 23802 24544 23808
rect 24596 23662 24624 24006
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24492 23248 24544 23254
rect 24492 23190 24544 23196
rect 24400 23180 24452 23186
rect 24400 23122 24452 23128
rect 24412 21690 24440 23122
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24504 21570 24532 23190
rect 24412 21554 24532 21570
rect 24400 21548 24532 21554
rect 24452 21542 24532 21548
rect 24400 21490 24452 21496
rect 24308 21004 24360 21010
rect 24308 20946 24360 20952
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24228 17338 24256 17682
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24320 16674 24348 20946
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24412 19310 24440 19654
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24228 16646 24348 16674
rect 24228 12986 24256 16646
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 24320 16046 24348 16526
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24320 15570 24348 15982
rect 24308 15564 24360 15570
rect 24308 15506 24360 15512
rect 24320 15162 24348 15506
rect 24308 15156 24360 15162
rect 24308 15098 24360 15104
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24044 12406 24164 12434
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23492 10606 23520 11222
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23400 10130 23428 10406
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23492 9178 23520 10542
rect 24044 10538 24072 12406
rect 24412 12186 24440 19246
rect 24504 16522 24532 21542
rect 24688 21162 24716 25774
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24780 25430 24808 25706
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24872 24596 24900 27628
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 24964 25362 24992 26318
rect 25056 25838 25084 28562
rect 25148 27130 25176 31980
rect 25240 31890 25268 32302
rect 25228 31884 25280 31890
rect 25228 31826 25280 31832
rect 25228 31748 25280 31754
rect 25228 31690 25280 31696
rect 25240 27606 25268 31690
rect 25332 30598 25360 32966
rect 25596 32914 25648 32920
rect 25608 32824 25636 32914
rect 25424 32796 25636 32824
rect 25424 32230 25452 32796
rect 25504 32360 25556 32366
rect 25504 32302 25556 32308
rect 25412 32224 25464 32230
rect 25412 32166 25464 32172
rect 25516 31958 25544 32302
rect 25700 32178 25728 40446
rect 25780 40384 25832 40390
rect 25780 40326 25832 40332
rect 25792 39982 25820 40326
rect 25780 39976 25832 39982
rect 25780 39918 25832 39924
rect 26160 39574 26188 40480
rect 26252 40050 26280 41006
rect 26344 40526 26372 41006
rect 26332 40520 26384 40526
rect 26332 40462 26384 40468
rect 26240 40044 26292 40050
rect 26240 39986 26292 39992
rect 26344 39846 26372 40462
rect 26528 39982 26556 42502
rect 26620 42362 26648 44202
rect 26709 43548 27017 43568
rect 26709 43546 26715 43548
rect 26771 43546 26795 43548
rect 26851 43546 26875 43548
rect 26931 43546 26955 43548
rect 27011 43546 27017 43548
rect 26771 43494 26773 43546
rect 26953 43494 26955 43546
rect 26709 43492 26715 43494
rect 26771 43492 26795 43494
rect 26851 43492 26875 43494
rect 26931 43492 26955 43494
rect 27011 43492 27017 43494
rect 26709 43472 27017 43492
rect 26884 43240 26936 43246
rect 26936 43200 27016 43228
rect 26884 43182 26936 43188
rect 26988 42702 27016 43200
rect 26976 42696 27028 42702
rect 26976 42638 27028 42644
rect 26709 42460 27017 42480
rect 26709 42458 26715 42460
rect 26771 42458 26795 42460
rect 26851 42458 26875 42460
rect 26931 42458 26955 42460
rect 27011 42458 27017 42460
rect 26771 42406 26773 42458
rect 26953 42406 26955 42458
rect 26709 42404 26715 42406
rect 26771 42404 26795 42406
rect 26851 42404 26875 42406
rect 26931 42404 26955 42406
rect 27011 42404 27017 42406
rect 26709 42384 27017 42404
rect 26608 42356 26660 42362
rect 26608 42298 26660 42304
rect 26700 42152 26752 42158
rect 26700 42094 26752 42100
rect 26792 42152 26844 42158
rect 26792 42094 26844 42100
rect 26712 41614 26740 42094
rect 26804 41818 26832 42094
rect 26884 42084 26936 42090
rect 26884 42026 26936 42032
rect 26792 41812 26844 41818
rect 26792 41754 26844 41760
rect 26804 41682 26832 41754
rect 26792 41676 26844 41682
rect 26792 41618 26844 41624
rect 26700 41608 26752 41614
rect 26700 41550 26752 41556
rect 26896 41546 26924 42026
rect 26884 41540 26936 41546
rect 26884 41482 26936 41488
rect 26608 41472 26660 41478
rect 26608 41414 26660 41420
rect 26620 41002 26648 41414
rect 26709 41372 27017 41392
rect 26709 41370 26715 41372
rect 26771 41370 26795 41372
rect 26851 41370 26875 41372
rect 26931 41370 26955 41372
rect 27011 41370 27017 41372
rect 26771 41318 26773 41370
rect 26953 41318 26955 41370
rect 26709 41316 26715 41318
rect 26771 41316 26795 41318
rect 26851 41316 26875 41318
rect 26931 41316 26955 41318
rect 27011 41316 27017 41318
rect 26709 41296 27017 41316
rect 27080 41070 27108 44406
rect 27632 44334 27660 44678
rect 29368 44464 29420 44470
rect 29368 44406 29420 44412
rect 27620 44328 27672 44334
rect 27620 44270 27672 44276
rect 27344 44260 27396 44266
rect 27344 44202 27396 44208
rect 27160 43852 27212 43858
rect 27160 43794 27212 43800
rect 27172 43450 27200 43794
rect 27160 43444 27212 43450
rect 27160 43386 27212 43392
rect 27160 43104 27212 43110
rect 27160 43046 27212 43052
rect 27172 42158 27200 43046
rect 27160 42152 27212 42158
rect 27356 42106 27384 44202
rect 27632 43654 27660 44270
rect 29380 43994 29408 44406
rect 30656 44192 30708 44198
rect 30656 44134 30708 44140
rect 29368 43988 29420 43994
rect 29368 43930 29420 43936
rect 27620 43648 27672 43654
rect 27620 43590 27672 43596
rect 28724 43648 28776 43654
rect 28724 43590 28776 43596
rect 27632 43246 27660 43590
rect 27620 43240 27672 43246
rect 27620 43182 27672 43188
rect 28632 43240 28684 43246
rect 28632 43182 28684 43188
rect 27632 42838 27660 43182
rect 27712 43172 27764 43178
rect 27712 43114 27764 43120
rect 28264 43172 28316 43178
rect 28264 43114 28316 43120
rect 27620 42832 27672 42838
rect 27620 42774 27672 42780
rect 27724 42770 27752 43114
rect 28276 42906 28304 43114
rect 28264 42900 28316 42906
rect 28264 42842 28316 42848
rect 27712 42764 27764 42770
rect 27712 42706 27764 42712
rect 27804 42696 27856 42702
rect 27804 42638 27856 42644
rect 27896 42696 27948 42702
rect 27896 42638 27948 42644
rect 27436 42560 27488 42566
rect 27436 42502 27488 42508
rect 27160 42094 27212 42100
rect 27264 42078 27384 42106
rect 27160 41472 27212 41478
rect 27160 41414 27212 41420
rect 27068 41064 27120 41070
rect 27068 41006 27120 41012
rect 26608 40996 26660 41002
rect 26608 40938 26660 40944
rect 26516 39976 26568 39982
rect 26516 39918 26568 39924
rect 26332 39840 26384 39846
rect 26332 39782 26384 39788
rect 26148 39568 26200 39574
rect 26148 39510 26200 39516
rect 25780 39092 25832 39098
rect 25780 39034 25832 39040
rect 25792 38826 25820 39034
rect 26240 38888 26292 38894
rect 26240 38830 26292 38836
rect 25780 38820 25832 38826
rect 25780 38762 25832 38768
rect 25792 37738 25820 38762
rect 26252 38486 26280 38830
rect 26240 38480 26292 38486
rect 26240 38422 26292 38428
rect 26240 38276 26292 38282
rect 26240 38218 26292 38224
rect 26252 37806 26280 38218
rect 26240 37800 26292 37806
rect 26240 37742 26292 37748
rect 25780 37732 25832 37738
rect 25780 37674 25832 37680
rect 26252 37398 26280 37742
rect 26240 37392 26292 37398
rect 26240 37334 26292 37340
rect 26056 36576 26108 36582
rect 26056 36518 26108 36524
rect 26068 36378 26096 36518
rect 26056 36372 26108 36378
rect 26056 36314 26108 36320
rect 26056 36236 26108 36242
rect 26056 36178 26108 36184
rect 26068 34950 26096 36178
rect 26252 35086 26280 37334
rect 26344 36378 26372 39782
rect 26424 39500 26476 39506
rect 26424 39442 26476 39448
rect 26436 38758 26464 39442
rect 26528 39098 26556 39918
rect 26516 39092 26568 39098
rect 26516 39034 26568 39040
rect 26620 38894 26648 40938
rect 26709 40284 27017 40304
rect 26709 40282 26715 40284
rect 26771 40282 26795 40284
rect 26851 40282 26875 40284
rect 26931 40282 26955 40284
rect 27011 40282 27017 40284
rect 26771 40230 26773 40282
rect 26953 40230 26955 40282
rect 26709 40228 26715 40230
rect 26771 40228 26795 40230
rect 26851 40228 26875 40230
rect 26931 40228 26955 40230
rect 27011 40228 27017 40230
rect 26709 40208 27017 40228
rect 27172 39506 27200 41414
rect 27264 40730 27292 42078
rect 27344 42016 27396 42022
rect 27344 41958 27396 41964
rect 27252 40724 27304 40730
rect 27252 40666 27304 40672
rect 27356 40662 27384 41958
rect 27344 40656 27396 40662
rect 27344 40598 27396 40604
rect 27448 40594 27476 42502
rect 27528 42016 27580 42022
rect 27528 41958 27580 41964
rect 27252 40588 27304 40594
rect 27252 40530 27304 40536
rect 27436 40588 27488 40594
rect 27436 40530 27488 40536
rect 27264 39574 27292 40530
rect 27344 40384 27396 40390
rect 27344 40326 27396 40332
rect 27252 39568 27304 39574
rect 27252 39510 27304 39516
rect 27160 39500 27212 39506
rect 27160 39442 27212 39448
rect 26709 39196 27017 39216
rect 26709 39194 26715 39196
rect 26771 39194 26795 39196
rect 26851 39194 26875 39196
rect 26931 39194 26955 39196
rect 27011 39194 27017 39196
rect 26771 39142 26773 39194
rect 26953 39142 26955 39194
rect 26709 39140 26715 39142
rect 26771 39140 26795 39142
rect 26851 39140 26875 39142
rect 26931 39140 26955 39142
rect 27011 39140 27017 39142
rect 26709 39120 27017 39140
rect 26608 38888 26660 38894
rect 26608 38830 26660 38836
rect 26424 38752 26476 38758
rect 26476 38712 26556 38740
rect 26424 38694 26476 38700
rect 26424 37732 26476 37738
rect 26424 37674 26476 37680
rect 26436 37466 26464 37674
rect 26424 37460 26476 37466
rect 26424 37402 26476 37408
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 26332 36372 26384 36378
rect 26332 36314 26384 36320
rect 26436 36174 26464 37062
rect 26528 36310 26556 38712
rect 26608 38412 26660 38418
rect 26608 38354 26660 38360
rect 26620 38010 26648 38354
rect 26709 38108 27017 38128
rect 26709 38106 26715 38108
rect 26771 38106 26795 38108
rect 26851 38106 26875 38108
rect 26931 38106 26955 38108
rect 27011 38106 27017 38108
rect 26771 38054 26773 38106
rect 26953 38054 26955 38106
rect 26709 38052 26715 38054
rect 26771 38052 26795 38054
rect 26851 38052 26875 38054
rect 26931 38052 26955 38054
rect 27011 38052 27017 38054
rect 26709 38032 27017 38052
rect 26608 38004 26660 38010
rect 26608 37946 26660 37952
rect 27264 37942 27292 39510
rect 27356 38554 27384 40326
rect 27436 39840 27488 39846
rect 27436 39782 27488 39788
rect 27448 39386 27476 39782
rect 27540 39506 27568 41958
rect 27816 41546 27844 42638
rect 27908 42294 27936 42638
rect 27896 42288 27948 42294
rect 27896 42230 27948 42236
rect 28264 42016 28316 42022
rect 28264 41958 28316 41964
rect 27804 41540 27856 41546
rect 27804 41482 27856 41488
rect 27896 41472 27948 41478
rect 27896 41414 27948 41420
rect 27620 40452 27672 40458
rect 27620 40394 27672 40400
rect 27528 39500 27580 39506
rect 27528 39442 27580 39448
rect 27448 39358 27568 39386
rect 27436 39296 27488 39302
rect 27436 39238 27488 39244
rect 27344 38548 27396 38554
rect 27344 38490 27396 38496
rect 27356 38010 27384 38490
rect 27344 38004 27396 38010
rect 27344 37946 27396 37952
rect 27252 37936 27304 37942
rect 27252 37878 27304 37884
rect 27356 37398 27384 37946
rect 27252 37392 27304 37398
rect 27252 37334 27304 37340
rect 27344 37392 27396 37398
rect 27344 37334 27396 37340
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 26709 37020 27017 37040
rect 26709 37018 26715 37020
rect 26771 37018 26795 37020
rect 26851 37018 26875 37020
rect 26931 37018 26955 37020
rect 27011 37018 27017 37020
rect 26771 36966 26773 37018
rect 26953 36966 26955 37018
rect 26709 36964 26715 36966
rect 26771 36964 26795 36966
rect 26851 36964 26875 36966
rect 26931 36964 26955 36966
rect 27011 36964 27017 36966
rect 26709 36944 27017 36964
rect 27080 36904 27108 37198
rect 26804 36876 27108 36904
rect 26804 36718 26832 36876
rect 26608 36712 26660 36718
rect 26608 36654 26660 36660
rect 26792 36712 26844 36718
rect 26792 36654 26844 36660
rect 27068 36712 27120 36718
rect 27068 36654 27120 36660
rect 27160 36712 27212 36718
rect 27160 36654 27212 36660
rect 26516 36304 26568 36310
rect 26516 36246 26568 36252
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26056 34944 26108 34950
rect 26056 34886 26108 34892
rect 26068 34542 26096 34886
rect 26056 34536 26108 34542
rect 26056 34478 26108 34484
rect 26148 34468 26200 34474
rect 26148 34410 26200 34416
rect 26056 34128 26108 34134
rect 26056 34070 26108 34076
rect 25872 33924 25924 33930
rect 25872 33866 25924 33872
rect 25780 33380 25832 33386
rect 25780 33322 25832 33328
rect 25792 32978 25820 33322
rect 25884 33114 25912 33866
rect 25872 33108 25924 33114
rect 25872 33050 25924 33056
rect 25780 32972 25832 32978
rect 25780 32914 25832 32920
rect 25792 32230 25820 32914
rect 25884 32910 25912 33050
rect 26068 33046 26096 34070
rect 26160 33862 26188 34410
rect 26148 33856 26200 33862
rect 26148 33798 26200 33804
rect 26160 33130 26188 33798
rect 26252 33454 26280 35022
rect 26528 34542 26556 36246
rect 26620 35562 26648 36654
rect 26804 36106 26832 36654
rect 26792 36100 26844 36106
rect 26792 36042 26844 36048
rect 26709 35932 27017 35952
rect 26709 35930 26715 35932
rect 26771 35930 26795 35932
rect 26851 35930 26875 35932
rect 26931 35930 26955 35932
rect 27011 35930 27017 35932
rect 26771 35878 26773 35930
rect 26953 35878 26955 35930
rect 26709 35876 26715 35878
rect 26771 35876 26795 35878
rect 26851 35876 26875 35878
rect 26931 35876 26955 35878
rect 27011 35876 27017 35878
rect 26709 35856 27017 35876
rect 26608 35556 26660 35562
rect 26608 35498 26660 35504
rect 26620 34746 26648 35498
rect 27080 35290 27108 36654
rect 27172 36378 27200 36654
rect 27160 36372 27212 36378
rect 27160 36314 27212 36320
rect 27160 35828 27212 35834
rect 27160 35770 27212 35776
rect 27172 35494 27200 35770
rect 27264 35630 27292 37334
rect 27356 36310 27384 37334
rect 27344 36304 27396 36310
rect 27344 36246 27396 36252
rect 27448 36242 27476 39238
rect 27540 38894 27568 39358
rect 27632 38894 27660 40394
rect 27712 39500 27764 39506
rect 27712 39442 27764 39448
rect 27724 39098 27752 39442
rect 27804 39364 27856 39370
rect 27804 39306 27856 39312
rect 27712 39092 27764 39098
rect 27712 39034 27764 39040
rect 27816 38962 27844 39306
rect 27804 38956 27856 38962
rect 27804 38898 27856 38904
rect 27528 38888 27580 38894
rect 27528 38830 27580 38836
rect 27620 38888 27672 38894
rect 27620 38830 27672 38836
rect 27540 38486 27568 38830
rect 27528 38480 27580 38486
rect 27528 38422 27580 38428
rect 27712 38344 27764 38350
rect 27712 38286 27764 38292
rect 27528 38004 27580 38010
rect 27528 37946 27580 37952
rect 27540 37194 27568 37946
rect 27620 37800 27672 37806
rect 27620 37742 27672 37748
rect 27632 37466 27660 37742
rect 27620 37460 27672 37466
rect 27620 37402 27672 37408
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 27528 37188 27580 37194
rect 27528 37130 27580 37136
rect 27528 36576 27580 36582
rect 27528 36518 27580 36524
rect 27436 36236 27488 36242
rect 27436 36178 27488 36184
rect 27344 36168 27396 36174
rect 27344 36110 27396 36116
rect 27356 35834 27384 36110
rect 27344 35828 27396 35834
rect 27344 35770 27396 35776
rect 27540 35714 27568 36518
rect 27632 36242 27660 37266
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 27632 35766 27660 36178
rect 27724 35766 27752 38286
rect 27816 38214 27844 38898
rect 27908 38894 27936 41414
rect 28172 40520 28224 40526
rect 28172 40462 28224 40468
rect 28184 40050 28212 40462
rect 28172 40044 28224 40050
rect 28172 39986 28224 39992
rect 28184 39642 28212 39986
rect 28172 39636 28224 39642
rect 28172 39578 28224 39584
rect 27988 39432 28040 39438
rect 27988 39374 28040 39380
rect 28000 38894 28028 39374
rect 28172 39364 28224 39370
rect 28172 39306 28224 39312
rect 27896 38888 27948 38894
rect 27896 38830 27948 38836
rect 27988 38888 28040 38894
rect 27988 38830 28040 38836
rect 27896 38344 27948 38350
rect 27896 38286 27948 38292
rect 27804 38208 27856 38214
rect 27804 38150 27856 38156
rect 27816 36650 27844 38150
rect 27908 37874 27936 38286
rect 27896 37868 27948 37874
rect 27896 37810 27948 37816
rect 27896 37664 27948 37670
rect 27896 37606 27948 37612
rect 27908 36718 27936 37606
rect 28000 36786 28028 38830
rect 28184 38418 28212 39306
rect 28276 38894 28304 41958
rect 28644 41614 28672 43182
rect 28736 42770 28764 43590
rect 29184 43104 29236 43110
rect 29184 43046 29236 43052
rect 29552 43104 29604 43110
rect 29552 43046 29604 43052
rect 28724 42764 28776 42770
rect 28724 42706 28776 42712
rect 29196 42702 29224 43046
rect 29368 42764 29420 42770
rect 29368 42706 29420 42712
rect 29184 42696 29236 42702
rect 29184 42638 29236 42644
rect 28908 42220 28960 42226
rect 28908 42162 28960 42168
rect 28632 41608 28684 41614
rect 28632 41550 28684 41556
rect 28644 41138 28672 41550
rect 28632 41132 28684 41138
rect 28632 41074 28684 41080
rect 28644 40594 28672 41074
rect 28632 40588 28684 40594
rect 28632 40530 28684 40536
rect 28920 40526 28948 42162
rect 29092 42152 29144 42158
rect 29092 42094 29144 42100
rect 29000 41744 29052 41750
rect 29000 41686 29052 41692
rect 28540 40520 28592 40526
rect 28540 40462 28592 40468
rect 28908 40520 28960 40526
rect 28908 40462 28960 40468
rect 28448 39976 28500 39982
rect 28448 39918 28500 39924
rect 28552 39930 28580 40462
rect 28356 39636 28408 39642
rect 28356 39578 28408 39584
rect 28264 38888 28316 38894
rect 28264 38830 28316 38836
rect 28368 38654 28396 39578
rect 28460 39030 28488 39918
rect 28552 39914 28672 39930
rect 28552 39908 28684 39914
rect 28552 39902 28632 39908
rect 28552 39506 28580 39902
rect 28632 39850 28684 39856
rect 29012 39642 29040 41686
rect 29000 39636 29052 39642
rect 29000 39578 29052 39584
rect 29104 39506 29132 42094
rect 29196 42022 29224 42638
rect 29380 42362 29408 42706
rect 29368 42356 29420 42362
rect 29368 42298 29420 42304
rect 29276 42152 29328 42158
rect 29276 42094 29328 42100
rect 29184 42016 29236 42022
rect 29184 41958 29236 41964
rect 29196 39574 29224 41958
rect 29288 39982 29316 42094
rect 29460 40044 29512 40050
rect 29460 39986 29512 39992
rect 29276 39976 29328 39982
rect 29276 39918 29328 39924
rect 29184 39568 29236 39574
rect 29184 39510 29236 39516
rect 28540 39500 28592 39506
rect 28540 39442 28592 39448
rect 29092 39500 29144 39506
rect 29092 39442 29144 39448
rect 28448 39024 28500 39030
rect 28448 38966 28500 38972
rect 28448 38752 28500 38758
rect 28448 38694 28500 38700
rect 28276 38626 28396 38654
rect 28276 38486 28304 38626
rect 28264 38480 28316 38486
rect 28264 38422 28316 38428
rect 28172 38412 28224 38418
rect 28460 38400 28488 38694
rect 28552 38486 28580 39442
rect 28632 39432 28684 39438
rect 28632 39374 28684 39380
rect 28540 38480 28592 38486
rect 28540 38422 28592 38428
rect 28460 38372 28497 38400
rect 28172 38354 28224 38360
rect 28080 38208 28132 38214
rect 28080 38150 28132 38156
rect 28092 37738 28120 38150
rect 28184 37806 28212 38354
rect 28469 38264 28497 38372
rect 28644 38350 28672 39374
rect 29288 39370 29316 39918
rect 29472 39642 29500 39986
rect 29460 39636 29512 39642
rect 29460 39578 29512 39584
rect 29276 39364 29328 39370
rect 29276 39306 29328 39312
rect 29092 39296 29144 39302
rect 29092 39238 29144 39244
rect 28724 38412 28776 38418
rect 28724 38354 28776 38360
rect 28632 38344 28684 38350
rect 28632 38286 28684 38292
rect 28460 38236 28497 38264
rect 28172 37800 28224 37806
rect 28172 37742 28224 37748
rect 28080 37732 28132 37738
rect 28080 37674 28132 37680
rect 28184 37448 28212 37742
rect 28092 37420 28212 37448
rect 28092 37330 28120 37420
rect 28080 37324 28132 37330
rect 28080 37266 28132 37272
rect 28172 37324 28224 37330
rect 28172 37266 28224 37272
rect 27988 36780 28040 36786
rect 27988 36722 28040 36728
rect 27896 36712 27948 36718
rect 27896 36654 27948 36660
rect 27804 36644 27856 36650
rect 27804 36586 27856 36592
rect 27448 35686 27568 35714
rect 27620 35760 27672 35766
rect 27620 35702 27672 35708
rect 27712 35760 27764 35766
rect 27712 35702 27764 35708
rect 27252 35624 27304 35630
rect 27252 35566 27304 35572
rect 27160 35488 27212 35494
rect 27160 35430 27212 35436
rect 27068 35284 27120 35290
rect 27068 35226 27120 35232
rect 27264 34950 27292 35566
rect 27448 35154 27476 35686
rect 27816 35630 27844 36586
rect 27896 35760 27948 35766
rect 27896 35702 27948 35708
rect 27712 35624 27764 35630
rect 27712 35566 27764 35572
rect 27804 35624 27856 35630
rect 27804 35566 27856 35572
rect 27528 35556 27580 35562
rect 27528 35498 27580 35504
rect 27436 35148 27488 35154
rect 27436 35090 27488 35096
rect 27252 34944 27304 34950
rect 27252 34886 27304 34892
rect 26709 34844 27017 34864
rect 26709 34842 26715 34844
rect 26771 34842 26795 34844
rect 26851 34842 26875 34844
rect 26931 34842 26955 34844
rect 27011 34842 27017 34844
rect 26771 34790 26773 34842
rect 26953 34790 26955 34842
rect 26709 34788 26715 34790
rect 26771 34788 26795 34790
rect 26851 34788 26875 34790
rect 26931 34788 26955 34790
rect 27011 34788 27017 34790
rect 26709 34768 27017 34788
rect 26608 34740 26660 34746
rect 26608 34682 26660 34688
rect 26608 34604 26660 34610
rect 26608 34546 26660 34552
rect 26516 34536 26568 34542
rect 26516 34478 26568 34484
rect 26516 34060 26568 34066
rect 26516 34002 26568 34008
rect 26240 33448 26292 33454
rect 26240 33390 26292 33396
rect 26160 33102 26280 33130
rect 26056 33040 26108 33046
rect 26056 32982 26108 32988
rect 26148 32972 26200 32978
rect 26148 32914 26200 32920
rect 25872 32904 25924 32910
rect 25872 32846 25924 32852
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26068 32230 26096 32846
rect 26160 32366 26188 32914
rect 26148 32360 26200 32366
rect 26148 32302 26200 32308
rect 25608 32150 25728 32178
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 25964 32224 26016 32230
rect 25964 32166 26016 32172
rect 26056 32224 26108 32230
rect 26056 32166 26108 32172
rect 25504 31952 25556 31958
rect 25504 31894 25556 31900
rect 25412 31884 25464 31890
rect 25412 31826 25464 31832
rect 25424 31278 25452 31826
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 25516 31278 25544 31758
rect 25608 31754 25636 32150
rect 25976 31890 26004 32166
rect 25780 31884 25832 31890
rect 25780 31826 25832 31832
rect 25964 31884 26016 31890
rect 25964 31826 26016 31832
rect 25596 31748 25648 31754
rect 25596 31690 25648 31696
rect 25792 31668 25820 31826
rect 26068 31668 26096 32166
rect 26252 32026 26280 33102
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 26240 32020 26292 32026
rect 26240 31962 26292 31968
rect 26344 31822 26372 33050
rect 26528 31822 26556 34002
rect 26620 33114 26648 34546
rect 27540 34202 27568 35498
rect 27724 34202 27752 35566
rect 27908 35154 27936 35702
rect 28000 35698 28028 36722
rect 28080 36712 28132 36718
rect 28080 36654 28132 36660
rect 28092 35834 28120 36654
rect 28080 35828 28132 35834
rect 28080 35770 28132 35776
rect 27988 35692 28040 35698
rect 27988 35634 28040 35640
rect 27896 35148 27948 35154
rect 27896 35090 27948 35096
rect 28080 34400 28132 34406
rect 28080 34342 28132 34348
rect 27528 34196 27580 34202
rect 27528 34138 27580 34144
rect 27712 34196 27764 34202
rect 27712 34138 27764 34144
rect 27988 34060 28040 34066
rect 27988 34002 28040 34008
rect 26709 33756 27017 33776
rect 26709 33754 26715 33756
rect 26771 33754 26795 33756
rect 26851 33754 26875 33756
rect 26931 33754 26955 33756
rect 27011 33754 27017 33756
rect 26771 33702 26773 33754
rect 26953 33702 26955 33754
rect 26709 33700 26715 33702
rect 26771 33700 26795 33702
rect 26851 33700 26875 33702
rect 26931 33700 26955 33702
rect 27011 33700 27017 33702
rect 26709 33680 27017 33700
rect 28000 33454 28028 34002
rect 28092 33522 28120 34342
rect 28080 33516 28132 33522
rect 28080 33458 28132 33464
rect 27988 33448 28040 33454
rect 27988 33390 28040 33396
rect 26608 33108 26660 33114
rect 26608 33050 26660 33056
rect 27620 32768 27672 32774
rect 27620 32710 27672 32716
rect 26709 32668 27017 32688
rect 26709 32666 26715 32668
rect 26771 32666 26795 32668
rect 26851 32666 26875 32668
rect 26931 32666 26955 32668
rect 27011 32666 27017 32668
rect 26771 32614 26773 32666
rect 26953 32614 26955 32666
rect 26709 32612 26715 32614
rect 26771 32612 26795 32614
rect 26851 32612 26875 32614
rect 26931 32612 26955 32614
rect 27011 32612 27017 32614
rect 26709 32592 27017 32612
rect 26608 32564 26660 32570
rect 26608 32506 26660 32512
rect 26620 32026 26648 32506
rect 27528 32292 27580 32298
rect 27528 32234 27580 32240
rect 27540 32026 27568 32234
rect 26608 32020 26660 32026
rect 26608 31962 26660 31968
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 26332 31816 26384 31822
rect 25792 31640 26096 31668
rect 26252 31776 26332 31804
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25412 31272 25464 31278
rect 25412 31214 25464 31220
rect 25504 31272 25556 31278
rect 25504 31214 25556 31220
rect 25424 30802 25452 31214
rect 25608 31210 25636 31282
rect 26148 31272 26200 31278
rect 26148 31214 26200 31220
rect 25596 31204 25648 31210
rect 25596 31146 25648 31152
rect 25504 31136 25556 31142
rect 25504 31078 25556 31084
rect 25412 30796 25464 30802
rect 25412 30738 25464 30744
rect 25320 30592 25372 30598
rect 25320 30534 25372 30540
rect 25332 30190 25360 30534
rect 25320 30184 25372 30190
rect 25320 30126 25372 30132
rect 25320 29028 25372 29034
rect 25320 28970 25372 28976
rect 25228 27600 25280 27606
rect 25228 27542 25280 27548
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25148 26994 25176 27066
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25136 26444 25188 26450
rect 25136 26386 25188 26392
rect 25044 25832 25096 25838
rect 25044 25774 25096 25780
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 25044 25356 25096 25362
rect 25044 25298 25096 25304
rect 24952 24676 25004 24682
rect 24952 24618 25004 24624
rect 24780 24568 24900 24596
rect 24780 24206 24808 24568
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24872 22778 24900 24210
rect 24964 24070 24992 24618
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 25056 23662 25084 25298
rect 25148 24818 25176 26386
rect 25240 25158 25268 26862
rect 25332 25362 25360 28970
rect 25412 27600 25464 27606
rect 25412 27542 25464 27548
rect 25424 25362 25452 27542
rect 25320 25356 25372 25362
rect 25320 25298 25372 25304
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25424 25242 25452 25298
rect 25332 25214 25452 25242
rect 25228 25152 25280 25158
rect 25228 25094 25280 25100
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24964 22234 24992 23258
rect 25148 23202 25176 24142
rect 25240 23322 25268 25094
rect 25332 24274 25360 25214
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 25424 24206 25452 25094
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25320 23588 25372 23594
rect 25320 23530 25372 23536
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25148 23174 25268 23202
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 24952 22228 25004 22234
rect 24952 22170 25004 22176
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24596 21134 24716 21162
rect 24596 20806 24624 21134
rect 24780 21010 24808 21966
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24872 21486 24900 21898
rect 24964 21622 24992 22170
rect 25056 22098 25084 22714
rect 25136 22500 25188 22506
rect 25136 22442 25188 22448
rect 25148 22234 25176 22442
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 24952 21616 25004 21622
rect 24952 21558 25004 21564
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24596 20534 24624 20742
rect 24584 20528 24636 20534
rect 24584 20470 24636 20476
rect 24780 20398 24808 20946
rect 24964 20806 24992 21422
rect 25148 21146 25176 21422
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 24768 20392 24820 20398
rect 24768 20334 24820 20340
rect 25148 20330 25176 20742
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24596 18766 24624 18906
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 24688 16250 24716 16594
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24688 15434 24716 16186
rect 24964 15706 24992 20198
rect 25240 18170 25268 23174
rect 25332 21690 25360 23530
rect 25516 22094 25544 31078
rect 26160 30802 26188 31214
rect 26252 31210 26280 31776
rect 26332 31758 26384 31764
rect 26516 31816 26568 31822
rect 26516 31758 26568 31764
rect 26332 31680 26384 31686
rect 26332 31622 26384 31628
rect 26344 31346 26372 31622
rect 26620 31362 26648 31962
rect 26709 31580 27017 31600
rect 26709 31578 26715 31580
rect 26771 31578 26795 31580
rect 26851 31578 26875 31580
rect 26931 31578 26955 31580
rect 27011 31578 27017 31580
rect 26771 31526 26773 31578
rect 26953 31526 26955 31578
rect 26709 31524 26715 31526
rect 26771 31524 26795 31526
rect 26851 31524 26875 31526
rect 26931 31524 26955 31526
rect 27011 31524 27017 31526
rect 26709 31504 27017 31524
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 26528 31334 26648 31362
rect 27540 31346 27568 31962
rect 27632 31482 27660 32710
rect 28000 32570 28028 33390
rect 28184 32978 28212 37266
rect 28460 36854 28488 38236
rect 28736 37670 28764 38354
rect 28908 38208 28960 38214
rect 28908 38150 28960 38156
rect 28920 37806 28948 38150
rect 29000 37936 29052 37942
rect 29000 37878 29052 37884
rect 28908 37800 28960 37806
rect 28908 37742 28960 37748
rect 28724 37664 28776 37670
rect 28724 37606 28776 37612
rect 28448 36848 28500 36854
rect 28448 36790 28500 36796
rect 28264 36032 28316 36038
rect 28264 35974 28316 35980
rect 28276 35630 28304 35974
rect 29012 35766 29040 37878
rect 29104 36310 29132 39238
rect 29368 38344 29420 38350
rect 29368 38286 29420 38292
rect 29380 37874 29408 38286
rect 29184 37868 29236 37874
rect 29184 37810 29236 37816
rect 29368 37868 29420 37874
rect 29368 37810 29420 37816
rect 29196 37670 29224 37810
rect 29184 37664 29236 37670
rect 29184 37606 29236 37612
rect 29196 36650 29224 37606
rect 29184 36644 29236 36650
rect 29184 36586 29236 36592
rect 29092 36304 29144 36310
rect 29092 36246 29144 36252
rect 29000 35760 29052 35766
rect 29000 35702 29052 35708
rect 28816 35692 28868 35698
rect 28816 35634 28868 35640
rect 28264 35624 28316 35630
rect 28264 35566 28316 35572
rect 28540 35284 28592 35290
rect 28540 35226 28592 35232
rect 28356 34060 28408 34066
rect 28356 34002 28408 34008
rect 28368 33454 28396 34002
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 28368 33046 28396 33390
rect 28448 33312 28500 33318
rect 28448 33254 28500 33260
rect 28356 33040 28408 33046
rect 28356 32982 28408 32988
rect 28172 32972 28224 32978
rect 28172 32914 28224 32920
rect 27988 32564 28040 32570
rect 27988 32506 28040 32512
rect 27988 32292 28040 32298
rect 27988 32234 28040 32240
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27344 31340 27396 31346
rect 26240 31204 26292 31210
rect 26240 31146 26292 31152
rect 25688 30796 25740 30802
rect 25688 30738 25740 30744
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25608 30326 25636 30670
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 25608 30122 25636 30262
rect 25700 30190 25728 30738
rect 25688 30184 25740 30190
rect 25688 30126 25740 30132
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 25596 30116 25648 30122
rect 25596 30058 25648 30064
rect 25608 29850 25636 30058
rect 25596 29844 25648 29850
rect 25596 29786 25648 29792
rect 25700 28626 25728 30126
rect 26056 29708 26108 29714
rect 26160 29696 26188 30126
rect 26108 29668 26188 29696
rect 26056 29650 26108 29656
rect 26056 29504 26108 29510
rect 26056 29446 26108 29452
rect 25688 28620 25740 28626
rect 25688 28562 25740 28568
rect 25872 28620 25924 28626
rect 25872 28562 25924 28568
rect 25884 28490 25912 28562
rect 25872 28484 25924 28490
rect 25872 28426 25924 28432
rect 25688 27872 25740 27878
rect 25688 27814 25740 27820
rect 25780 27872 25832 27878
rect 25884 27860 25912 28426
rect 25832 27832 25912 27860
rect 25780 27814 25832 27820
rect 25700 27470 25728 27814
rect 25688 27464 25740 27470
rect 25608 27424 25688 27452
rect 25608 24834 25636 27424
rect 25688 27406 25740 27412
rect 25688 26852 25740 26858
rect 25688 26794 25740 26800
rect 25700 25906 25728 26794
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 25608 24806 25728 24834
rect 25700 24426 25728 24806
rect 25424 22066 25544 22094
rect 25608 24398 25728 24426
rect 25320 21684 25372 21690
rect 25320 21626 25372 21632
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25056 18142 25268 18170
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24584 15088 24636 15094
rect 24584 15030 24636 15036
rect 24596 14482 24624 15030
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24688 14618 24716 14962
rect 24780 14890 24808 15438
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24872 15162 24900 15302
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24964 15094 24992 15642
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24768 14884 24820 14890
rect 24768 14826 24820 14832
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24780 14414 24808 14826
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24872 14618 24900 14758
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24780 14006 24808 14350
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24872 14006 24900 14214
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24964 13870 24992 14418
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24780 13190 24808 13670
rect 24964 13530 24992 13806
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24504 12442 24532 12718
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24136 12158 24440 12186
rect 24136 11354 24164 12158
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24412 11898 24440 12038
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24320 11354 24348 11494
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24032 10532 24084 10538
rect 24032 10474 24084 10480
rect 24044 10130 24072 10474
rect 24032 10124 24084 10130
rect 24032 10066 24084 10072
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23584 9042 23612 9658
rect 24032 9512 24084 9518
rect 24032 9454 24084 9460
rect 23848 9104 23900 9110
rect 23848 9046 23900 9052
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23400 8566 23428 8910
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23492 8022 23520 8774
rect 23584 8634 23612 8842
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23308 6956 23612 6984
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23492 6186 23520 6802
rect 23584 6746 23612 6956
rect 23768 6934 23796 7142
rect 23756 6928 23808 6934
rect 23756 6870 23808 6876
rect 23860 6798 23888 9046
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23952 8430 23980 8774
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23940 7744 23992 7750
rect 23940 7686 23992 7692
rect 23848 6792 23900 6798
rect 23584 6718 23796 6746
rect 23848 6734 23900 6740
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23676 6390 23704 6598
rect 23664 6384 23716 6390
rect 23664 6326 23716 6332
rect 23768 6322 23796 6718
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23860 6254 23888 6734
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23308 5846 23336 6054
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 23492 5166 23520 6122
rect 23860 5914 23888 6190
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23952 5778 23980 7686
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23492 4826 23520 5102
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23676 4078 23704 5034
rect 23952 4758 23980 5714
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23584 2990 23612 3674
rect 23676 3074 23704 4014
rect 23676 3046 23796 3074
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23400 1358 23428 2926
rect 23676 2650 23704 3046
rect 23768 2990 23796 3046
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23388 1352 23440 1358
rect 23388 1294 23440 1300
rect 20076 944 20128 950
rect 19352 870 19472 898
rect 20076 886 20128 892
rect 23020 944 23072 950
rect 23020 886 23072 892
rect 23204 944 23256 950
rect 23204 886 23256 892
rect 15936 808 15988 814
rect 15936 750 15988 756
rect 16764 808 16816 814
rect 16764 750 16816 756
rect 16948 808 17000 814
rect 16948 750 17000 756
rect 17316 808 17368 814
rect 19352 800 19380 870
rect 19444 814 19472 870
rect 19432 808 19484 814
rect 17316 750 17368 756
rect 14648 672 14700 678
rect 14648 614 14700 620
rect 19338 0 19394 800
rect 19432 750 19484 756
rect 20168 672 20220 678
rect 20168 614 20220 620
rect 20180 406 20208 614
rect 21557 572 21865 592
rect 21557 570 21563 572
rect 21619 570 21643 572
rect 21699 570 21723 572
rect 21779 570 21803 572
rect 21859 570 21865 572
rect 21619 518 21621 570
rect 21801 518 21803 570
rect 21557 516 21563 518
rect 21619 516 21643 518
rect 21699 516 21723 518
rect 21779 516 21803 518
rect 21859 516 21865 518
rect 21557 496 21865 516
rect 23032 474 23060 886
rect 24044 814 24072 9454
rect 24136 7750 24164 11290
rect 24504 10810 24532 11834
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24504 9722 24532 10746
rect 24596 10606 24624 12310
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 11218 24808 12174
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24964 11014 24992 11630
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 10198 24624 10542
rect 24584 10192 24636 10198
rect 24584 10134 24636 10140
rect 24492 9716 24544 9722
rect 24492 9658 24544 9664
rect 24504 8090 24532 9658
rect 24596 9518 24624 10134
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24780 8634 24808 9046
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24412 5846 24440 6598
rect 24504 5914 24532 7346
rect 24688 6662 24716 7890
rect 24780 7546 24808 8298
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24872 7342 24900 9386
rect 24964 8566 24992 10950
rect 25056 10010 25084 18142
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 17542 25268 18022
rect 25332 17814 25360 18566
rect 25320 17808 25372 17814
rect 25320 17750 25372 17756
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25240 17134 25268 17478
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25240 16114 25268 17070
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25136 14544 25188 14550
rect 25136 14486 25188 14492
rect 25148 14414 25176 14486
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 25136 14408 25188 14414
rect 25136 14350 25188 14356
rect 25148 13938 25176 14350
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25136 13932 25188 13938
rect 25136 13874 25188 13880
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 25148 13394 25176 13670
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25148 11014 25176 12786
rect 25240 12374 25268 14214
rect 25332 12442 25360 14418
rect 25424 12714 25452 22066
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25516 20602 25544 21286
rect 25608 20942 25636 24398
rect 25688 24336 25740 24342
rect 25688 24278 25740 24284
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25608 19310 25636 20878
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 25516 12850 25544 19110
rect 25700 16130 25728 24278
rect 25792 23186 25820 27814
rect 25872 26240 25924 26246
rect 25872 26182 25924 26188
rect 25884 25838 25912 26182
rect 26068 25838 26096 29446
rect 26160 29170 26188 29668
rect 26240 29708 26292 29714
rect 26240 29650 26292 29656
rect 26252 29306 26280 29650
rect 26240 29300 26292 29306
rect 26240 29242 26292 29248
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 26160 28558 26188 28698
rect 26252 28626 26280 29242
rect 26528 29186 26556 31334
rect 27344 31282 27396 31288
rect 27528 31340 27580 31346
rect 27528 31282 27580 31288
rect 26608 31272 26660 31278
rect 26608 31214 26660 31220
rect 27252 31272 27304 31278
rect 27252 31214 27304 31220
rect 26620 29714 26648 31214
rect 27068 31136 27120 31142
rect 27068 31078 27120 31084
rect 26709 30492 27017 30512
rect 26709 30490 26715 30492
rect 26771 30490 26795 30492
rect 26851 30490 26875 30492
rect 26931 30490 26955 30492
rect 27011 30490 27017 30492
rect 26771 30438 26773 30490
rect 26953 30438 26955 30490
rect 26709 30436 26715 30438
rect 26771 30436 26795 30438
rect 26851 30436 26875 30438
rect 26931 30436 26955 30438
rect 27011 30436 27017 30438
rect 26709 30416 27017 30436
rect 27080 30138 27108 31078
rect 27264 30802 27292 31214
rect 27252 30796 27304 30802
rect 27252 30738 27304 30744
rect 27356 30734 27384 31282
rect 27436 31204 27488 31210
rect 27436 31146 27488 31152
rect 27344 30728 27396 30734
rect 27344 30670 27396 30676
rect 27356 30274 27384 30670
rect 27448 30666 27476 31146
rect 27620 31136 27672 31142
rect 27620 31078 27672 31084
rect 27632 30938 27660 31078
rect 27620 30932 27672 30938
rect 27620 30874 27672 30880
rect 27620 30796 27672 30802
rect 27620 30738 27672 30744
rect 27436 30660 27488 30666
rect 27436 30602 27488 30608
rect 27356 30246 27568 30274
rect 26988 30122 27108 30138
rect 27344 30184 27396 30190
rect 27344 30126 27396 30132
rect 26976 30116 27108 30122
rect 27028 30110 27108 30116
rect 27160 30116 27212 30122
rect 26976 30058 27028 30064
rect 27160 30058 27212 30064
rect 27172 29782 27200 30058
rect 27160 29776 27212 29782
rect 27160 29718 27212 29724
rect 26608 29708 26660 29714
rect 26608 29650 26660 29656
rect 26709 29404 27017 29424
rect 26709 29402 26715 29404
rect 26771 29402 26795 29404
rect 26851 29402 26875 29404
rect 26931 29402 26955 29404
rect 27011 29402 27017 29404
rect 26771 29350 26773 29402
rect 26953 29350 26955 29402
rect 26709 29348 26715 29350
rect 26771 29348 26795 29350
rect 26851 29348 26875 29350
rect 26931 29348 26955 29350
rect 27011 29348 27017 29350
rect 26709 29328 27017 29348
rect 26528 29158 26648 29186
rect 26516 29028 26568 29034
rect 26516 28970 26568 28976
rect 26528 28762 26556 28970
rect 26516 28756 26568 28762
rect 26516 28698 26568 28704
rect 26240 28620 26292 28626
rect 26240 28562 26292 28568
rect 26148 28552 26200 28558
rect 26148 28494 26200 28500
rect 26160 27606 26188 28494
rect 26620 27878 26648 29158
rect 26709 28316 27017 28336
rect 26709 28314 26715 28316
rect 26771 28314 26795 28316
rect 26851 28314 26875 28316
rect 26931 28314 26955 28316
rect 27011 28314 27017 28316
rect 26771 28262 26773 28314
rect 26953 28262 26955 28314
rect 26709 28260 26715 28262
rect 26771 28260 26795 28262
rect 26851 28260 26875 28262
rect 26931 28260 26955 28262
rect 27011 28260 27017 28262
rect 26709 28240 27017 28260
rect 26424 27872 26476 27878
rect 26424 27814 26476 27820
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 26332 26784 26384 26790
rect 26332 26726 26384 26732
rect 26240 26512 26292 26518
rect 26240 26454 26292 26460
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 25872 25832 25924 25838
rect 25872 25774 25924 25780
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 25964 25696 26016 25702
rect 26160 25684 26188 26386
rect 25964 25638 26016 25644
rect 26068 25656 26188 25684
rect 25976 25498 26004 25638
rect 25964 25492 26016 25498
rect 25964 25434 26016 25440
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25780 21616 25832 21622
rect 25780 21558 25832 21564
rect 25792 21010 25820 21558
rect 25884 21146 25912 25230
rect 25964 25220 26016 25226
rect 26068 25208 26096 25656
rect 26148 25356 26200 25362
rect 26148 25298 26200 25304
rect 26016 25180 26096 25208
rect 25964 25162 26016 25168
rect 25976 24274 26004 25162
rect 25964 24268 26016 24274
rect 25964 24210 26016 24216
rect 26056 23588 26108 23594
rect 26056 23530 26108 23536
rect 26068 22982 26096 23530
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 26068 22250 26096 22918
rect 25976 22222 26096 22250
rect 25976 22166 26004 22222
rect 25964 22160 26016 22166
rect 25964 22102 26016 22108
rect 25872 21140 25924 21146
rect 25872 21082 25924 21088
rect 25976 21078 26004 22102
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 26068 21418 26096 21898
rect 26160 21486 26188 25298
rect 26252 24682 26280 26454
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26344 24342 26372 26726
rect 26436 25974 26464 27814
rect 27252 27396 27304 27402
rect 27252 27338 27304 27344
rect 26709 27228 27017 27248
rect 26709 27226 26715 27228
rect 26771 27226 26795 27228
rect 26851 27226 26875 27228
rect 26931 27226 26955 27228
rect 27011 27226 27017 27228
rect 26771 27174 26773 27226
rect 26953 27174 26955 27226
rect 26709 27172 26715 27174
rect 26771 27172 26795 27174
rect 26851 27172 26875 27174
rect 26931 27172 26955 27174
rect 27011 27172 27017 27174
rect 26709 27152 27017 27172
rect 26608 26920 26660 26926
rect 26608 26862 26660 26868
rect 26976 26920 27028 26926
rect 26976 26862 27028 26868
rect 26516 26240 26568 26246
rect 26516 26182 26568 26188
rect 26424 25968 26476 25974
rect 26424 25910 26476 25916
rect 26528 25906 26556 26182
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26516 25764 26568 25770
rect 26516 25706 26568 25712
rect 26424 25696 26476 25702
rect 26424 25638 26476 25644
rect 26436 24886 26464 25638
rect 26424 24880 26476 24886
rect 26424 24822 26476 24828
rect 26424 24744 26476 24750
rect 26424 24686 26476 24692
rect 26436 24410 26464 24686
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26332 24336 26384 24342
rect 26332 24278 26384 24284
rect 26344 24070 26372 24278
rect 26332 24064 26384 24070
rect 26332 24006 26384 24012
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25780 21004 25832 21010
rect 25780 20946 25832 20952
rect 26160 20058 26188 21422
rect 26252 20398 26280 22510
rect 26344 22166 26372 23462
rect 26528 23322 26556 25706
rect 26620 24954 26648 26862
rect 26988 26228 27016 26862
rect 27264 26382 27292 27338
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 27160 26308 27212 26314
rect 27160 26250 27212 26256
rect 26988 26200 27108 26228
rect 26709 26140 27017 26160
rect 26709 26138 26715 26140
rect 26771 26138 26795 26140
rect 26851 26138 26875 26140
rect 26931 26138 26955 26140
rect 27011 26138 27017 26140
rect 26771 26086 26773 26138
rect 26953 26086 26955 26138
rect 26709 26084 26715 26086
rect 26771 26084 26795 26086
rect 26851 26084 26875 26086
rect 26931 26084 26955 26086
rect 27011 26084 27017 26086
rect 26709 26064 27017 26084
rect 26700 25968 26752 25974
rect 26700 25910 26752 25916
rect 26712 25226 26740 25910
rect 26700 25220 26752 25226
rect 26700 25162 26752 25168
rect 26709 25052 27017 25072
rect 26709 25050 26715 25052
rect 26771 25050 26795 25052
rect 26851 25050 26875 25052
rect 26931 25050 26955 25052
rect 27011 25050 27017 25052
rect 26771 24998 26773 25050
rect 26953 24998 26955 25050
rect 26709 24996 26715 24998
rect 26771 24996 26795 24998
rect 26851 24996 26875 24998
rect 26931 24996 26955 24998
rect 27011 24996 27017 24998
rect 26709 24976 27017 24996
rect 26608 24948 26660 24954
rect 26608 24890 26660 24896
rect 27080 24750 27108 26200
rect 26608 24744 26660 24750
rect 26608 24686 26660 24692
rect 27068 24744 27120 24750
rect 27068 24686 27120 24692
rect 26516 23316 26568 23322
rect 26516 23258 26568 23264
rect 26620 22778 26648 24686
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 26712 24274 26740 24550
rect 27080 24410 27108 24686
rect 27172 24682 27200 26250
rect 27356 25974 27384 30126
rect 27540 28490 27568 30246
rect 27632 29510 27660 30738
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 27724 30394 27752 30670
rect 27804 30592 27856 30598
rect 27804 30534 27856 30540
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27816 29782 27844 30534
rect 27804 29776 27856 29782
rect 27804 29718 27856 29724
rect 28000 29714 28028 32234
rect 28080 31272 28132 31278
rect 28080 31214 28132 31220
rect 28092 30326 28120 31214
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 28184 29850 28212 32914
rect 28460 32366 28488 33254
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28276 30870 28304 31282
rect 28264 30864 28316 30870
rect 28264 30806 28316 30812
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28172 29844 28224 29850
rect 28172 29786 28224 29792
rect 27988 29708 28040 29714
rect 27988 29650 28040 29656
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27632 28626 27660 29446
rect 28184 29170 28212 29786
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 27528 28484 27580 28490
rect 27528 28426 27580 28432
rect 27540 28082 27568 28426
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27632 28014 27660 28562
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27620 27872 27672 27878
rect 27620 27814 27672 27820
rect 28264 27872 28316 27878
rect 28264 27814 28316 27820
rect 27528 27668 27580 27674
rect 27528 27610 27580 27616
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27448 25974 27476 26862
rect 27540 26858 27568 27610
rect 27632 27334 27660 27814
rect 27988 27464 28040 27470
rect 27988 27406 28040 27412
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27632 27130 27660 27270
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27528 26852 27580 26858
rect 27528 26794 27580 26800
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27908 26450 27936 26726
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 27896 26444 27948 26450
rect 27896 26386 27948 26392
rect 27528 26376 27580 26382
rect 27528 26318 27580 26324
rect 27540 26042 27568 26318
rect 27724 26042 27752 26386
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27712 26036 27764 26042
rect 27712 25978 27764 25984
rect 27344 25968 27396 25974
rect 27344 25910 27396 25916
rect 27436 25968 27488 25974
rect 27436 25910 27488 25916
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27264 25362 27292 25842
rect 27252 25356 27304 25362
rect 27252 25298 27304 25304
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27068 24404 27120 24410
rect 27068 24346 27120 24352
rect 27172 24342 27200 24618
rect 27160 24336 27212 24342
rect 27160 24278 27212 24284
rect 26700 24268 26752 24274
rect 26700 24210 26752 24216
rect 26709 23964 27017 23984
rect 26709 23962 26715 23964
rect 26771 23962 26795 23964
rect 26851 23962 26875 23964
rect 26931 23962 26955 23964
rect 27011 23962 27017 23964
rect 26771 23910 26773 23962
rect 26953 23910 26955 23962
rect 26709 23908 26715 23910
rect 26771 23908 26795 23910
rect 26851 23908 26875 23910
rect 26931 23908 26955 23910
rect 27011 23908 27017 23910
rect 26709 23888 27017 23908
rect 27264 23866 27292 25298
rect 27448 25158 27476 25910
rect 27436 25152 27488 25158
rect 27436 25094 27488 25100
rect 27344 24676 27396 24682
rect 27344 24618 27396 24624
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27068 23792 27120 23798
rect 27068 23734 27120 23740
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26712 23050 26740 23462
rect 26700 23044 26752 23050
rect 26700 22986 26752 22992
rect 26709 22876 27017 22896
rect 26709 22874 26715 22876
rect 26771 22874 26795 22876
rect 26851 22874 26875 22876
rect 26931 22874 26955 22876
rect 27011 22874 27017 22876
rect 26771 22822 26773 22874
rect 26953 22822 26955 22874
rect 26709 22820 26715 22822
rect 26771 22820 26795 22822
rect 26851 22820 26875 22822
rect 26931 22820 26955 22822
rect 27011 22820 27017 22822
rect 26709 22800 27017 22820
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26424 22704 26476 22710
rect 27080 22658 27108 23734
rect 27160 23588 27212 23594
rect 27160 23530 27212 23536
rect 27172 23118 27200 23530
rect 27264 23118 27292 23802
rect 27356 23798 27384 24618
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 26424 22646 26476 22652
rect 26436 22234 26464 22646
rect 26896 22630 27108 22658
rect 26896 22574 26924 22630
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 27068 22568 27120 22574
rect 27068 22510 27120 22516
rect 26424 22228 26476 22234
rect 26424 22170 26476 22176
rect 26332 22160 26384 22166
rect 26332 22102 26384 22108
rect 27080 21894 27108 22510
rect 27172 22234 27200 23054
rect 27448 23050 27476 25094
rect 27540 24818 27568 25978
rect 28000 25294 28028 27406
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28080 26376 28132 26382
rect 28080 26318 28132 26324
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27436 23044 27488 23050
rect 27436 22986 27488 22992
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27264 22574 27292 22918
rect 27540 22710 27568 24754
rect 27632 24750 27660 25094
rect 28092 24818 28120 26318
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 27620 24744 27672 24750
rect 27620 24686 27672 24692
rect 27804 24744 27856 24750
rect 28184 24698 28212 27270
rect 28276 25838 28304 27814
rect 28460 27062 28488 30194
rect 28552 28422 28580 35226
rect 28828 34066 28856 35634
rect 29012 34678 29040 35702
rect 29000 34672 29052 34678
rect 29000 34614 29052 34620
rect 29012 34082 29040 34614
rect 28816 34060 28868 34066
rect 29012 34054 29132 34082
rect 29196 34066 29224 36586
rect 29564 35222 29592 43046
rect 30668 42770 30696 44134
rect 30944 43450 30972 44678
rect 31116 44328 31168 44334
rect 31116 44270 31168 44276
rect 31024 43648 31076 43654
rect 31024 43590 31076 43596
rect 30932 43444 30984 43450
rect 30932 43386 30984 43392
rect 30656 42764 30708 42770
rect 30656 42706 30708 42712
rect 30380 42560 30432 42566
rect 30380 42502 30432 42508
rect 29920 42220 29972 42226
rect 29920 42162 29972 42168
rect 29932 39982 29960 42162
rect 30012 42084 30064 42090
rect 30012 42026 30064 42032
rect 30024 41818 30052 42026
rect 30288 42016 30340 42022
rect 30288 41958 30340 41964
rect 30012 41812 30064 41818
rect 30012 41754 30064 41760
rect 30300 41070 30328 41958
rect 30288 41064 30340 41070
rect 30288 41006 30340 41012
rect 30288 40588 30340 40594
rect 30288 40530 30340 40536
rect 30300 40186 30328 40530
rect 30392 40186 30420 42502
rect 30472 42152 30524 42158
rect 30472 42094 30524 42100
rect 30484 41682 30512 42094
rect 30944 41818 30972 43386
rect 31036 43330 31064 43590
rect 31128 43450 31156 44270
rect 31116 43444 31168 43450
rect 31116 43386 31168 43392
rect 31036 43302 31156 43330
rect 31128 43246 31156 43302
rect 31116 43240 31168 43246
rect 31116 43182 31168 43188
rect 31128 42158 31156 43182
rect 31208 42764 31260 42770
rect 31208 42706 31260 42712
rect 31116 42152 31168 42158
rect 31116 42094 31168 42100
rect 30932 41812 30984 41818
rect 30932 41754 30984 41760
rect 30472 41676 30524 41682
rect 30472 41618 30524 41624
rect 30484 41562 30512 41618
rect 30484 41534 30604 41562
rect 30472 41472 30524 41478
rect 30472 41414 30524 41420
rect 30288 40180 30340 40186
rect 30288 40122 30340 40128
rect 30380 40180 30432 40186
rect 30380 40122 30432 40128
rect 30484 40066 30512 41414
rect 30576 40934 30604 41534
rect 30564 40928 30616 40934
rect 30564 40870 30616 40876
rect 30564 40384 30616 40390
rect 30564 40326 30616 40332
rect 30208 40038 30512 40066
rect 29920 39976 29972 39982
rect 29920 39918 29972 39924
rect 29644 39840 29696 39846
rect 29644 39782 29696 39788
rect 29656 39574 29684 39782
rect 29644 39568 29696 39574
rect 29644 39510 29696 39516
rect 29932 39438 29960 39918
rect 29920 39432 29972 39438
rect 29920 39374 29972 39380
rect 29932 39098 29960 39374
rect 29920 39092 29972 39098
rect 29920 39034 29972 39040
rect 30104 36236 30156 36242
rect 30104 36178 30156 36184
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 29736 36032 29788 36038
rect 29736 35974 29788 35980
rect 29644 35624 29696 35630
rect 29644 35566 29696 35572
rect 29552 35216 29604 35222
rect 29552 35158 29604 35164
rect 29276 35080 29328 35086
rect 29656 35034 29684 35566
rect 29748 35290 29776 35974
rect 29828 35624 29880 35630
rect 29828 35566 29880 35572
rect 29736 35284 29788 35290
rect 29736 35226 29788 35232
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 29276 35022 29328 35028
rect 29288 34066 29316 35022
rect 29564 35006 29684 35034
rect 29564 34950 29592 35006
rect 29552 34944 29604 34950
rect 29552 34886 29604 34892
rect 29564 34066 29592 34886
rect 29644 34740 29696 34746
rect 29644 34682 29696 34688
rect 28816 34002 28868 34008
rect 28828 33454 28856 34002
rect 29104 33998 29132 34054
rect 29184 34060 29236 34066
rect 29184 34002 29236 34008
rect 29276 34060 29328 34066
rect 29276 34002 29328 34008
rect 29552 34060 29604 34066
rect 29552 34002 29604 34008
rect 29092 33992 29144 33998
rect 29092 33934 29144 33940
rect 29104 33590 29132 33934
rect 29092 33584 29144 33590
rect 29092 33526 29144 33532
rect 29288 33522 29316 34002
rect 29276 33516 29328 33522
rect 29276 33458 29328 33464
rect 29656 33454 29684 34682
rect 29748 34202 29776 35090
rect 29840 35086 29868 35566
rect 29828 35080 29880 35086
rect 29828 35022 29880 35028
rect 29932 34202 29960 36110
rect 30116 35630 30144 36178
rect 30104 35624 30156 35630
rect 30104 35566 30156 35572
rect 30116 34762 30144 35566
rect 30024 34746 30144 34762
rect 30012 34740 30144 34746
rect 30064 34734 30144 34740
rect 30012 34682 30064 34688
rect 29736 34196 29788 34202
rect 29736 34138 29788 34144
rect 29920 34196 29972 34202
rect 29920 34138 29972 34144
rect 30012 34060 30064 34066
rect 30012 34002 30064 34008
rect 29736 33584 29788 33590
rect 29736 33526 29788 33532
rect 28632 33448 28684 33454
rect 28632 33390 28684 33396
rect 28816 33448 28868 33454
rect 28816 33390 28868 33396
rect 29644 33448 29696 33454
rect 29644 33390 29696 33396
rect 28644 33046 28672 33390
rect 28632 33040 28684 33046
rect 28632 32982 28684 32988
rect 28644 32910 28672 32982
rect 29748 32978 29776 33526
rect 29828 33516 29880 33522
rect 29828 33458 29880 33464
rect 28816 32972 28868 32978
rect 28816 32914 28868 32920
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 28632 32904 28684 32910
rect 28632 32846 28684 32852
rect 28828 32026 28856 32914
rect 29840 32910 29868 33458
rect 30024 33454 30052 34002
rect 30012 33448 30064 33454
rect 29932 33408 30012 33436
rect 29932 32978 29960 33408
rect 30012 33390 30064 33396
rect 29920 32972 29972 32978
rect 29920 32914 29972 32920
rect 29828 32904 29880 32910
rect 29828 32846 29880 32852
rect 29000 32836 29052 32842
rect 29000 32778 29052 32784
rect 28816 32020 28868 32026
rect 28816 31962 28868 31968
rect 28816 29504 28868 29510
rect 28816 29446 28868 29452
rect 28632 29096 28684 29102
rect 28632 29038 28684 29044
rect 28644 28626 28672 29038
rect 28632 28620 28684 28626
rect 28632 28562 28684 28568
rect 28540 28416 28592 28422
rect 28540 28358 28592 28364
rect 28644 28014 28672 28562
rect 28724 28552 28776 28558
rect 28828 28506 28856 29446
rect 29012 29170 29040 32778
rect 29368 32768 29420 32774
rect 29368 32710 29420 32716
rect 29828 32768 29880 32774
rect 29828 32710 29880 32716
rect 29092 32292 29144 32298
rect 29092 32234 29144 32240
rect 29104 30938 29132 32234
rect 29380 31958 29408 32710
rect 29368 31952 29420 31958
rect 29368 31894 29420 31900
rect 29644 31884 29696 31890
rect 29840 31872 29868 32710
rect 29932 32570 29960 32914
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 29696 31844 29868 31872
rect 29644 31826 29696 31832
rect 29092 30932 29144 30938
rect 29092 30874 29144 30880
rect 29184 29844 29236 29850
rect 29184 29786 29236 29792
rect 29000 29164 29052 29170
rect 29000 29106 29052 29112
rect 29092 28960 29144 28966
rect 29092 28902 29144 28908
rect 29104 28626 29132 28902
rect 29092 28620 29144 28626
rect 29092 28562 29144 28568
rect 28776 28500 28856 28506
rect 28724 28494 28856 28500
rect 28908 28552 28960 28558
rect 28908 28494 28960 28500
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 28736 28478 28856 28494
rect 28632 28008 28684 28014
rect 28632 27950 28684 27956
rect 28828 27878 28856 28478
rect 28816 27872 28868 27878
rect 28816 27814 28868 27820
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28736 27334 28764 27406
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28448 27056 28500 27062
rect 28448 26998 28500 27004
rect 28736 26586 28764 27270
rect 28724 26580 28776 26586
rect 28724 26522 28776 26528
rect 28828 25906 28856 27814
rect 28920 27538 28948 28494
rect 29012 28218 29040 28494
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 29012 27606 29040 28154
rect 29104 28082 29132 28562
rect 29092 28076 29144 28082
rect 29092 28018 29144 28024
rect 29000 27600 29052 27606
rect 29000 27542 29052 27548
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 29104 26926 29132 28018
rect 29092 26920 29144 26926
rect 29092 26862 29144 26868
rect 28908 26784 28960 26790
rect 28908 26726 28960 26732
rect 28920 26450 28948 26726
rect 28908 26444 28960 26450
rect 28908 26386 28960 26392
rect 28816 25900 28868 25906
rect 28816 25842 28868 25848
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28816 25356 28868 25362
rect 28816 25298 28868 25304
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 27804 24686 27856 24692
rect 27816 24410 27844 24686
rect 28092 24670 28212 24698
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27528 22704 27580 22710
rect 27528 22646 27580 22652
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 26709 21788 27017 21808
rect 26709 21786 26715 21788
rect 26771 21786 26795 21788
rect 26851 21786 26875 21788
rect 26931 21786 26955 21788
rect 27011 21786 27017 21788
rect 26771 21734 26773 21786
rect 26953 21734 26955 21786
rect 26709 21732 26715 21734
rect 26771 21732 26795 21734
rect 26851 21732 26875 21734
rect 26931 21732 26955 21734
rect 27011 21732 27017 21734
rect 26709 21712 27017 21732
rect 27540 21690 27568 22034
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27540 21486 27568 21626
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26608 21344 26660 21350
rect 26608 21286 26660 21292
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26252 19854 26280 20334
rect 26344 19990 26372 21286
rect 26620 20330 26648 21286
rect 27160 20800 27212 20806
rect 27160 20742 27212 20748
rect 26709 20700 27017 20720
rect 26709 20698 26715 20700
rect 26771 20698 26795 20700
rect 26851 20698 26875 20700
rect 26931 20698 26955 20700
rect 27011 20698 27017 20700
rect 26771 20646 26773 20698
rect 26953 20646 26955 20698
rect 26709 20644 26715 20646
rect 26771 20644 26795 20646
rect 26851 20644 26875 20646
rect 26931 20644 26955 20646
rect 27011 20644 27017 20646
rect 26709 20624 27017 20644
rect 26608 20324 26660 20330
rect 26608 20266 26660 20272
rect 26332 19984 26384 19990
rect 26332 19926 26384 19932
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26252 18086 26280 19790
rect 26709 19612 27017 19632
rect 26709 19610 26715 19612
rect 26771 19610 26795 19612
rect 26851 19610 26875 19612
rect 26931 19610 26955 19612
rect 27011 19610 27017 19612
rect 26771 19558 26773 19610
rect 26953 19558 26955 19610
rect 26709 19556 26715 19558
rect 26771 19556 26795 19558
rect 26851 19556 26875 19558
rect 26931 19556 26955 19558
rect 27011 19556 27017 19558
rect 26709 19536 27017 19556
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26344 18698 26372 19110
rect 27172 18902 27200 20742
rect 27540 19922 27568 21422
rect 28092 21350 28120 24670
rect 28552 23662 28580 25230
rect 28828 24410 28856 25298
rect 29000 24744 29052 24750
rect 29000 24686 29052 24692
rect 29012 24614 29040 24686
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28816 24404 28868 24410
rect 28816 24346 28868 24352
rect 28816 24268 28868 24274
rect 28816 24210 28868 24216
rect 28828 23662 28856 24210
rect 29012 23730 29040 24550
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 28172 23656 28224 23662
rect 28172 23598 28224 23604
rect 28540 23656 28592 23662
rect 28540 23598 28592 23604
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28184 22574 28212 23598
rect 28448 23520 28500 23526
rect 28448 23462 28500 23468
rect 28460 22642 28488 23462
rect 28552 22642 28580 23598
rect 28828 23526 28856 23598
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28632 23180 28684 23186
rect 28632 23122 28684 23128
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28540 22636 28592 22642
rect 28540 22578 28592 22584
rect 28172 22568 28224 22574
rect 28172 22510 28224 22516
rect 28184 22098 28212 22510
rect 28264 22500 28316 22506
rect 28264 22442 28316 22448
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 28172 21956 28224 21962
rect 28172 21898 28224 21904
rect 28184 21486 28212 21898
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 28000 20398 28028 21286
rect 28092 20942 28120 21286
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 28092 20210 28120 20878
rect 28000 20182 28120 20210
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27160 18896 27212 18902
rect 27160 18838 27212 18844
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26332 18692 26384 18698
rect 26332 18634 26384 18640
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26344 17898 26372 18634
rect 26252 17870 26372 17898
rect 25872 17808 25924 17814
rect 25872 17750 25924 17756
rect 25884 16658 25912 17750
rect 26148 17128 26200 17134
rect 26148 17070 26200 17076
rect 26160 16794 26188 17070
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 25700 16102 25912 16130
rect 25780 15972 25832 15978
rect 25780 15914 25832 15920
rect 25792 15162 25820 15914
rect 25780 15156 25832 15162
rect 25780 15098 25832 15104
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25608 14278 25636 14418
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25608 13870 25636 14214
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25700 13734 25728 14010
rect 25884 13954 25912 16102
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 25964 14816 26016 14822
rect 25964 14758 26016 14764
rect 25976 14482 26004 14758
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25884 13926 26004 13954
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25700 12782 25728 13670
rect 25884 13274 25912 13806
rect 25976 13462 26004 13926
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 26068 13274 26096 15982
rect 26160 14958 26188 16594
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 26160 14550 26188 14894
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 26160 14414 26188 14486
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 25884 13246 26096 13274
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25412 12708 25464 12714
rect 25412 12650 25464 12656
rect 25872 12708 25924 12714
rect 25872 12650 25924 12656
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25228 12368 25280 12374
rect 25228 12310 25280 12316
rect 25332 11762 25360 12378
rect 25424 11898 25452 12378
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25424 11218 25452 11834
rect 25700 11694 25728 12582
rect 25884 12442 25912 12650
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25976 11830 26004 13126
rect 26068 12714 26096 13246
rect 26056 12708 26108 12714
rect 26056 12650 26108 12656
rect 26068 12306 26096 12650
rect 26056 12300 26108 12306
rect 26056 12242 26108 12248
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25412 11212 25464 11218
rect 25412 11154 25464 11160
rect 25700 11082 25728 11630
rect 25792 11218 25820 11698
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 25884 11354 25912 11630
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25976 11218 26004 11766
rect 25780 11212 25832 11218
rect 25780 11154 25832 11160
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25320 10056 25372 10062
rect 25056 9982 25176 10010
rect 25320 9998 25372 10004
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25056 8974 25084 9862
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25148 8838 25176 9982
rect 25332 9518 25360 9998
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 25516 8022 25544 10610
rect 25964 10532 26016 10538
rect 25964 10474 26016 10480
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25700 9110 25728 10406
rect 25976 10130 26004 10474
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 25964 10124 26016 10130
rect 25964 10066 26016 10072
rect 25976 9518 26004 10066
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 26160 9160 26188 10406
rect 26252 9450 26280 17870
rect 26436 17542 26464 18702
rect 27172 18630 27200 18838
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 26709 18524 27017 18544
rect 26709 18522 26715 18524
rect 26771 18522 26795 18524
rect 26851 18522 26875 18524
rect 26931 18522 26955 18524
rect 27011 18522 27017 18524
rect 26771 18470 26773 18522
rect 26953 18470 26955 18522
rect 26709 18468 26715 18470
rect 26771 18468 26795 18470
rect 26851 18468 26875 18470
rect 26931 18468 26955 18470
rect 27011 18468 27017 18470
rect 26709 18448 27017 18468
rect 27068 18420 27120 18426
rect 27068 18362 27120 18368
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26344 14482 26372 14894
rect 26332 14476 26384 14482
rect 26332 14418 26384 14424
rect 26436 14362 26464 17478
rect 26528 17134 26556 17682
rect 26709 17436 27017 17456
rect 26709 17434 26715 17436
rect 26771 17434 26795 17436
rect 26851 17434 26875 17436
rect 26931 17434 26955 17436
rect 27011 17434 27017 17436
rect 26771 17382 26773 17434
rect 26953 17382 26955 17434
rect 26709 17380 26715 17382
rect 26771 17380 26795 17382
rect 26851 17380 26875 17382
rect 26931 17380 26955 17382
rect 27011 17380 27017 17382
rect 26709 17360 27017 17380
rect 26516 17128 26568 17134
rect 26516 17070 26568 17076
rect 26528 15570 26556 17070
rect 26976 16992 27028 16998
rect 26976 16934 27028 16940
rect 26988 16794 27016 16934
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 26709 16348 27017 16368
rect 26709 16346 26715 16348
rect 26771 16346 26795 16348
rect 26851 16346 26875 16348
rect 26931 16346 26955 16348
rect 27011 16346 27017 16348
rect 26771 16294 26773 16346
rect 26953 16294 26955 16346
rect 26709 16292 26715 16294
rect 26771 16292 26795 16294
rect 26851 16292 26875 16294
rect 26931 16292 26955 16294
rect 27011 16292 27017 16294
rect 26709 16272 27017 16292
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26528 14958 26556 15506
rect 26620 15502 26648 15846
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26620 15026 26648 15438
rect 26709 15260 27017 15280
rect 26709 15258 26715 15260
rect 26771 15258 26795 15260
rect 26851 15258 26875 15260
rect 26931 15258 26955 15260
rect 27011 15258 27017 15260
rect 26771 15206 26773 15258
rect 26953 15206 26955 15258
rect 26709 15204 26715 15206
rect 26771 15204 26795 15206
rect 26851 15204 26875 15206
rect 26931 15204 26955 15206
rect 27011 15204 27017 15206
rect 26709 15184 27017 15204
rect 27080 15162 27108 18362
rect 27172 17202 27200 18566
rect 27264 18086 27292 19246
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27264 17814 27292 18022
rect 27252 17808 27304 17814
rect 27252 17750 27304 17756
rect 27252 17672 27304 17678
rect 27356 17660 27384 19314
rect 27712 19304 27764 19310
rect 27540 19252 27712 19258
rect 27540 19246 27764 19252
rect 27540 19242 27752 19246
rect 27528 19236 27752 19242
rect 27580 19230 27752 19236
rect 27528 19178 27580 19184
rect 27804 19168 27856 19174
rect 27804 19110 27856 19116
rect 27816 18970 27844 19110
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 28000 18834 28028 20182
rect 28080 19916 28132 19922
rect 28080 19858 28132 19864
rect 28092 18902 28120 19858
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 28080 18896 28132 18902
rect 28080 18838 28132 18844
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 27804 18148 27856 18154
rect 27804 18090 27856 18096
rect 27816 17882 27844 18090
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 27620 17808 27672 17814
rect 27620 17750 27672 17756
rect 27304 17632 27384 17660
rect 27252 17614 27304 17620
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27264 16590 27292 17614
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 27264 15502 27292 16526
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26344 14334 26464 14362
rect 26528 14346 26556 14894
rect 26516 14340 26568 14346
rect 26240 9444 26292 9450
rect 26240 9386 26292 9392
rect 26160 9132 26280 9160
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25872 9036 25924 9042
rect 25872 8978 25924 8984
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25504 8016 25556 8022
rect 25504 7958 25556 7964
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 24872 6934 24900 7278
rect 24860 6928 24912 6934
rect 24860 6870 24912 6876
rect 24872 6798 24900 6870
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24400 5840 24452 5846
rect 24400 5782 24452 5788
rect 24596 5302 24624 6190
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24780 5778 24808 6122
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24308 5024 24360 5030
rect 24308 4966 24360 4972
rect 24320 4690 24348 4966
rect 24308 4684 24360 4690
rect 24308 4626 24360 4632
rect 24504 3534 24532 5170
rect 24596 4078 24624 5238
rect 24688 4146 24716 5714
rect 24964 5370 24992 6802
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24860 5160 24912 5166
rect 24912 5120 24992 5148
rect 24860 5102 24912 5108
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24780 4162 24808 4626
rect 24676 4140 24728 4146
rect 24780 4134 24900 4162
rect 24676 4082 24728 4088
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24596 3738 24624 4014
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 24688 3602 24716 3674
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24320 3194 24348 3334
rect 24308 3188 24360 3194
rect 24308 3130 24360 3136
rect 24596 2650 24624 3538
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 24596 1426 24624 2586
rect 24688 2106 24716 3538
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24780 3058 24808 3470
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24780 2310 24808 2994
rect 24872 2650 24900 4134
rect 24964 3516 24992 5120
rect 25056 4690 25084 7686
rect 25516 7478 25544 7958
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25148 6866 25176 7142
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25516 6798 25544 7414
rect 25608 6866 25636 7890
rect 25700 7342 25728 8774
rect 25884 8566 25912 8978
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 25976 8090 26004 8366
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 25976 7342 26004 8026
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 25964 7336 26016 7342
rect 25964 7278 26016 7284
rect 25780 7268 25832 7274
rect 25780 7210 25832 7216
rect 25792 6866 25820 7210
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25780 6860 25832 6866
rect 25780 6802 25832 6808
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25424 5914 25452 6666
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 26068 5778 26096 8910
rect 26160 6186 26188 8978
rect 26252 6236 26280 9132
rect 26344 8362 26372 14334
rect 26516 14282 26568 14288
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 26436 13870 26464 14214
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26620 13326 26648 14962
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 26709 14172 27017 14192
rect 26709 14170 26715 14172
rect 26771 14170 26795 14172
rect 26851 14170 26875 14172
rect 26931 14170 26955 14172
rect 27011 14170 27017 14172
rect 26771 14118 26773 14170
rect 26953 14118 26955 14170
rect 26709 14116 26715 14118
rect 26771 14116 26795 14118
rect 26851 14116 26875 14118
rect 26931 14116 26955 14118
rect 27011 14116 27017 14118
rect 26709 14096 27017 14116
rect 27080 13394 27108 14214
rect 27172 14074 27200 14418
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27264 13802 27292 15438
rect 27252 13796 27304 13802
rect 27252 13738 27304 13744
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 27080 13274 27108 13330
rect 26620 12374 26648 13262
rect 27080 13246 27200 13274
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 26709 13084 27017 13104
rect 26709 13082 26715 13084
rect 26771 13082 26795 13084
rect 26851 13082 26875 13084
rect 26931 13082 26955 13084
rect 27011 13082 27017 13084
rect 26771 13030 26773 13082
rect 26953 13030 26955 13082
rect 26709 13028 26715 13030
rect 26771 13028 26795 13030
rect 26851 13028 26875 13030
rect 26931 13028 26955 13030
rect 27011 13028 27017 13030
rect 26709 13008 27017 13028
rect 27080 12782 27108 13126
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 26608 12368 26660 12374
rect 26608 12310 26660 12316
rect 27172 12102 27200 13246
rect 27356 12866 27384 16390
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27448 15570 27476 16186
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27540 14074 27568 15846
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27436 13728 27488 13734
rect 27436 13670 27488 13676
rect 27264 12850 27384 12866
rect 27252 12844 27384 12850
rect 27304 12838 27384 12844
rect 27252 12786 27304 12792
rect 27344 12776 27396 12782
rect 27344 12718 27396 12724
rect 27356 12442 27384 12718
rect 27344 12436 27396 12442
rect 27344 12378 27396 12384
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 26709 11996 27017 12016
rect 26709 11994 26715 11996
rect 26771 11994 26795 11996
rect 26851 11994 26875 11996
rect 26931 11994 26955 11996
rect 27011 11994 27017 11996
rect 26771 11942 26773 11994
rect 26953 11942 26955 11994
rect 26709 11940 26715 11942
rect 26771 11940 26795 11942
rect 26851 11940 26875 11942
rect 26931 11940 26955 11942
rect 27011 11940 27017 11942
rect 26709 11920 27017 11940
rect 27448 11914 27476 13670
rect 27632 12832 27660 17750
rect 27712 15972 27764 15978
rect 27712 15914 27764 15920
rect 27724 15706 27752 15914
rect 27712 15700 27764 15706
rect 27712 15642 27764 15648
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27632 12804 27752 12832
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27264 11886 27476 11914
rect 26516 11688 26568 11694
rect 26516 11630 26568 11636
rect 27160 11688 27212 11694
rect 27160 11630 27212 11636
rect 26528 10674 26556 11630
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 27068 11552 27120 11558
rect 27068 11494 27120 11500
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26620 10606 26648 11494
rect 26709 10908 27017 10928
rect 26709 10906 26715 10908
rect 26771 10906 26795 10908
rect 26851 10906 26875 10908
rect 26931 10906 26955 10908
rect 27011 10906 27017 10908
rect 26771 10854 26773 10906
rect 26953 10854 26955 10906
rect 26709 10852 26715 10854
rect 26771 10852 26795 10854
rect 26851 10852 26875 10854
rect 26931 10852 26955 10854
rect 27011 10852 27017 10854
rect 26709 10832 27017 10852
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26608 9988 26660 9994
rect 26608 9930 26660 9936
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 26436 9042 26464 9862
rect 26620 9518 26648 9930
rect 26709 9820 27017 9840
rect 26709 9818 26715 9820
rect 26771 9818 26795 9820
rect 26851 9818 26875 9820
rect 26931 9818 26955 9820
rect 27011 9818 27017 9820
rect 26771 9766 26773 9818
rect 26953 9766 26955 9818
rect 26709 9764 26715 9766
rect 26771 9764 26795 9766
rect 26851 9764 26875 9766
rect 26931 9764 26955 9766
rect 27011 9764 27017 9766
rect 26709 9744 27017 9764
rect 26516 9512 26568 9518
rect 26516 9454 26568 9460
rect 26608 9512 26660 9518
rect 27080 9500 27108 11494
rect 27172 11354 27200 11630
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27264 9722 27292 11886
rect 27540 11778 27568 12582
rect 27724 12374 27752 12804
rect 27908 12714 27936 13670
rect 27896 12708 27948 12714
rect 27896 12650 27948 12656
rect 27712 12368 27764 12374
rect 27712 12310 27764 12316
rect 27896 12096 27948 12102
rect 27896 12038 27948 12044
rect 27448 11750 27568 11778
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27356 11218 27384 11630
rect 27344 11212 27396 11218
rect 27344 11154 27396 11160
rect 27448 10962 27476 11750
rect 27908 11694 27936 12038
rect 27896 11688 27948 11694
rect 27896 11630 27948 11636
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 27540 11150 27568 11562
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27632 11218 27660 11494
rect 27908 11286 27936 11630
rect 27896 11280 27948 11286
rect 27896 11222 27948 11228
rect 27620 11212 27672 11218
rect 27620 11154 27672 11160
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 27448 10934 27568 10962
rect 27436 10600 27488 10606
rect 27436 10542 27488 10548
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27252 9716 27304 9722
rect 27252 9658 27304 9664
rect 27080 9472 27292 9500
rect 26608 9454 26660 9460
rect 26528 9042 26556 9454
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26436 8430 26464 8842
rect 26528 8430 26556 8978
rect 26620 8514 26648 9454
rect 26884 9444 26936 9450
rect 26936 9404 27108 9432
rect 26884 9386 26936 9392
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 26712 8906 26740 9318
rect 27080 8906 27108 9404
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 26709 8732 27017 8752
rect 26709 8730 26715 8732
rect 26771 8730 26795 8732
rect 26851 8730 26875 8732
rect 26931 8730 26955 8732
rect 27011 8730 27017 8732
rect 26771 8678 26773 8730
rect 26953 8678 26955 8730
rect 26709 8676 26715 8678
rect 26771 8676 26795 8678
rect 26851 8676 26875 8678
rect 26931 8676 26955 8678
rect 27011 8676 27017 8678
rect 26709 8656 27017 8676
rect 26620 8498 26740 8514
rect 26620 8492 26752 8498
rect 26620 8486 26700 8492
rect 26700 8434 26752 8440
rect 27080 8430 27108 8842
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 27068 8424 27120 8430
rect 27120 8384 27200 8412
rect 27068 8366 27120 8372
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26344 7410 26372 7686
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26436 6322 26464 8366
rect 26528 7954 26556 8366
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26528 7410 26556 7890
rect 27172 7886 27200 8384
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 26709 7644 27017 7664
rect 26709 7642 26715 7644
rect 26771 7642 26795 7644
rect 26851 7642 26875 7644
rect 26931 7642 26955 7644
rect 27011 7642 27017 7644
rect 26771 7590 26773 7642
rect 26953 7590 26955 7642
rect 26709 7588 26715 7590
rect 26771 7588 26795 7590
rect 26851 7588 26875 7590
rect 26931 7588 26955 7590
rect 27011 7588 27017 7590
rect 26709 7568 27017 7588
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26528 6866 26556 7346
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26709 6556 27017 6576
rect 26709 6554 26715 6556
rect 26771 6554 26795 6556
rect 26851 6554 26875 6556
rect 26931 6554 26955 6556
rect 27011 6554 27017 6556
rect 26771 6502 26773 6554
rect 26953 6502 26955 6554
rect 26709 6500 26715 6502
rect 26771 6500 26795 6502
rect 26851 6500 26875 6502
rect 26931 6500 26955 6502
rect 27011 6500 27017 6502
rect 26709 6480 27017 6500
rect 27080 6458 27108 7278
rect 27264 6644 27292 9472
rect 27356 8634 27384 10066
rect 27448 9586 27476 10542
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27448 8974 27476 9522
rect 27540 9518 27568 10934
rect 28000 10810 28028 18770
rect 28080 16516 28132 16522
rect 28080 16458 28132 16464
rect 27988 10804 28040 10810
rect 27988 10746 28040 10752
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27540 9042 27568 9318
rect 27632 9178 27660 9862
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27896 9036 27948 9042
rect 27896 8978 27948 8984
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 27448 8362 27476 8910
rect 27540 8430 27568 8978
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27448 8022 27476 8298
rect 27908 8090 27936 8978
rect 28092 8634 28120 16458
rect 28184 15638 28212 19382
rect 28172 15632 28224 15638
rect 28172 15574 28224 15580
rect 28184 14414 28212 15574
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 28184 13870 28212 14350
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 28172 10532 28224 10538
rect 28172 10474 28224 10480
rect 28080 8628 28132 8634
rect 28080 8570 28132 8576
rect 28184 8566 28212 10474
rect 28172 8560 28224 8566
rect 28172 8502 28224 8508
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27436 8016 27488 8022
rect 27436 7958 27488 7964
rect 27448 6798 27476 7958
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27632 7206 27660 7890
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27816 7342 27844 7686
rect 27804 7336 27856 7342
rect 27804 7278 27856 7284
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27632 6866 27660 7142
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27264 6616 27476 6644
rect 27068 6452 27120 6458
rect 27068 6394 27120 6400
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 26332 6248 26384 6254
rect 26252 6208 26332 6236
rect 26332 6190 26384 6196
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 26056 5772 26108 5778
rect 26056 5714 26108 5720
rect 25240 5574 25268 5714
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 26068 5302 26096 5714
rect 26160 5710 26188 6122
rect 26157 5704 26209 5710
rect 26157 5646 26209 5652
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 25136 5160 25188 5166
rect 25136 5102 25188 5108
rect 26056 5160 26108 5166
rect 26160 5148 26188 5646
rect 26108 5120 26188 5148
rect 26240 5160 26292 5166
rect 26056 5102 26108 5108
rect 26240 5102 26292 5108
rect 26344 5114 26372 6190
rect 26424 6112 26476 6118
rect 26424 6054 26476 6060
rect 26436 5778 26464 6054
rect 26620 5914 26648 6190
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25148 4622 25176 5102
rect 26056 4752 26108 4758
rect 26056 4694 26108 4700
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25148 3602 25176 4558
rect 25228 3664 25280 3670
rect 25228 3606 25280 3612
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 25044 3528 25096 3534
rect 24964 3488 25044 3516
rect 24964 3126 24992 3488
rect 25044 3470 25096 3476
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 24952 3120 25004 3126
rect 24952 3062 25004 3068
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24676 2100 24728 2106
rect 24676 2042 24728 2048
rect 24584 1420 24636 1426
rect 24584 1362 24636 1368
rect 24780 1290 24808 2246
rect 24872 2106 24900 2586
rect 25056 2514 25084 3334
rect 25148 2990 25176 3538
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25044 2508 25096 2514
rect 25044 2450 25096 2456
rect 24860 2100 24912 2106
rect 24860 2042 24912 2048
rect 25148 1426 25176 2926
rect 25240 2514 25268 3606
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 25228 2508 25280 2514
rect 25228 2450 25280 2456
rect 25700 1834 25728 3538
rect 25872 3392 25924 3398
rect 25872 3334 25924 3340
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25688 1828 25740 1834
rect 25688 1770 25740 1776
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 25596 1420 25648 1426
rect 25596 1362 25648 1368
rect 24768 1284 24820 1290
rect 24768 1226 24820 1232
rect 25504 1216 25556 1222
rect 25504 1158 25556 1164
rect 24872 870 24992 898
rect 24032 808 24084 814
rect 24872 800 24900 870
rect 24964 814 24992 870
rect 25516 814 25544 1158
rect 25608 950 25636 1362
rect 25700 1222 25728 1770
rect 25688 1216 25740 1222
rect 25688 1158 25740 1164
rect 25596 944 25648 950
rect 25596 886 25648 892
rect 25688 944 25740 950
rect 25688 886 25740 892
rect 24952 808 25004 814
rect 24032 750 24084 756
rect 23020 468 23072 474
rect 23020 410 23072 416
rect 20168 400 20220 406
rect 20168 342 20220 348
rect 24858 0 24914 800
rect 24952 750 25004 756
rect 25504 808 25556 814
rect 25504 750 25556 756
rect 24964 474 24992 750
rect 25700 678 25728 886
rect 25792 814 25820 2246
rect 25884 1902 25912 3334
rect 25976 2990 26004 4558
rect 26068 4078 26096 4694
rect 26148 4684 26200 4690
rect 26148 4626 26200 4632
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 26068 3058 26096 4014
rect 26056 3052 26108 3058
rect 26056 2994 26108 3000
rect 26160 3040 26188 4626
rect 26252 3738 26280 5102
rect 26344 5086 26464 5114
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26240 3052 26292 3058
rect 26160 3012 26240 3040
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26068 2650 26096 2994
rect 26056 2644 26108 2650
rect 25976 2604 26056 2632
rect 25872 1896 25924 1902
rect 25872 1838 25924 1844
rect 25976 882 26004 2604
rect 26056 2586 26108 2592
rect 26160 1222 26188 3012
rect 26240 2994 26292 3000
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26148 1216 26200 1222
rect 26148 1158 26200 1164
rect 25964 876 26016 882
rect 25964 818 26016 824
rect 26160 814 26188 1158
rect 26252 814 26280 2790
rect 26344 2106 26372 4966
rect 26436 4486 26464 5086
rect 26528 4826 26556 5850
rect 26608 5772 26660 5778
rect 26608 5714 26660 5720
rect 26516 4820 26568 4826
rect 26516 4762 26568 4768
rect 26424 4480 26476 4486
rect 26424 4422 26476 4428
rect 26620 3398 26648 5714
rect 26709 5468 27017 5488
rect 26709 5466 26715 5468
rect 26771 5466 26795 5468
rect 26851 5466 26875 5468
rect 26931 5466 26955 5468
rect 27011 5466 27017 5468
rect 26771 5414 26773 5466
rect 26953 5414 26955 5466
rect 26709 5412 26715 5414
rect 26771 5412 26795 5414
rect 26851 5412 26875 5414
rect 26931 5412 26955 5414
rect 27011 5412 27017 5414
rect 26709 5392 27017 5412
rect 27080 5370 27108 6394
rect 27344 6384 27396 6390
rect 27344 6326 27396 6332
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27068 5364 27120 5370
rect 27068 5306 27120 5312
rect 26884 5228 26936 5234
rect 26884 5170 26936 5176
rect 26896 4758 26924 5170
rect 27068 5160 27120 5166
rect 27068 5102 27120 5108
rect 26884 4752 26936 4758
rect 26884 4694 26936 4700
rect 26709 4380 27017 4400
rect 26709 4378 26715 4380
rect 26771 4378 26795 4380
rect 26851 4378 26875 4380
rect 26931 4378 26955 4380
rect 27011 4378 27017 4380
rect 26771 4326 26773 4378
rect 26953 4326 26955 4378
rect 26709 4324 26715 4326
rect 26771 4324 26795 4326
rect 26851 4324 26875 4326
rect 26931 4324 26955 4326
rect 27011 4324 27017 4326
rect 26709 4304 27017 4324
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 26620 2990 26648 3334
rect 26709 3292 27017 3312
rect 26709 3290 26715 3292
rect 26771 3290 26795 3292
rect 26851 3290 26875 3292
rect 26931 3290 26955 3292
rect 27011 3290 27017 3292
rect 26771 3238 26773 3290
rect 26953 3238 26955 3290
rect 26709 3236 26715 3238
rect 26771 3236 26795 3238
rect 26851 3236 26875 3238
rect 26931 3236 26955 3238
rect 27011 3236 27017 3238
rect 26709 3216 27017 3236
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26620 2582 26648 2926
rect 27080 2854 27108 5102
rect 27172 4146 27200 6258
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 27264 5098 27292 5646
rect 27356 5148 27384 6326
rect 27448 5302 27476 6616
rect 27540 6390 27568 6734
rect 27528 6384 27580 6390
rect 27528 6326 27580 6332
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27436 5296 27488 5302
rect 27436 5238 27488 5244
rect 27436 5160 27488 5166
rect 27356 5120 27436 5148
rect 27252 5092 27304 5098
rect 27252 5034 27304 5040
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 27160 2984 27212 2990
rect 27264 2972 27292 3674
rect 27212 2944 27292 2972
rect 27160 2926 27212 2932
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 26608 2576 26660 2582
rect 26608 2518 26660 2524
rect 26709 2204 27017 2224
rect 26709 2202 26715 2204
rect 26771 2202 26795 2204
rect 26851 2202 26875 2204
rect 26931 2202 26955 2204
rect 27011 2202 27017 2204
rect 26771 2150 26773 2202
rect 26953 2150 26955 2202
rect 26709 2148 26715 2150
rect 26771 2148 26795 2150
rect 26851 2148 26875 2150
rect 26931 2148 26955 2150
rect 27011 2148 27017 2150
rect 26709 2128 27017 2148
rect 26332 2100 26384 2106
rect 26332 2042 26384 2048
rect 26424 1964 26476 1970
rect 26424 1906 26476 1912
rect 26436 1426 26464 1906
rect 26424 1420 26476 1426
rect 26424 1362 26476 1368
rect 26709 1116 27017 1136
rect 26709 1114 26715 1116
rect 26771 1114 26795 1116
rect 26851 1114 26875 1116
rect 26931 1114 26955 1116
rect 27011 1114 27017 1116
rect 26771 1062 26773 1114
rect 26953 1062 26955 1114
rect 26709 1060 26715 1062
rect 26771 1060 26795 1062
rect 26851 1060 26875 1062
rect 26931 1060 26955 1062
rect 27011 1060 27017 1062
rect 26709 1040 27017 1060
rect 27172 882 27200 2926
rect 27356 2922 27384 5120
rect 27436 5102 27488 5108
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 27448 4282 27476 4966
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 27540 4146 27568 6190
rect 27632 5778 27660 6802
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 27908 6254 27936 6598
rect 27896 6248 27948 6254
rect 27896 6190 27948 6196
rect 27620 5772 27672 5778
rect 27620 5714 27672 5720
rect 27804 5364 27856 5370
rect 27804 5306 27856 5312
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27632 4826 27660 5102
rect 27712 5024 27764 5030
rect 27712 4966 27764 4972
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27724 4758 27752 4966
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27540 3602 27568 4082
rect 27816 3738 27844 5306
rect 27988 4548 28040 4554
rect 27988 4490 28040 4496
rect 28000 4078 28028 4490
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 28276 3738 28304 22442
rect 28460 22094 28488 22578
rect 28368 22066 28488 22094
rect 28368 22030 28396 22066
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28460 21842 28488 22066
rect 28552 22030 28580 22578
rect 28644 22098 28672 23122
rect 28724 23112 28776 23118
rect 28724 23054 28776 23060
rect 28736 22710 28764 23054
rect 28724 22704 28776 22710
rect 28724 22646 28776 22652
rect 28736 22574 28764 22646
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 28736 22166 28764 22510
rect 28828 22506 28856 23462
rect 28816 22500 28868 22506
rect 28816 22442 28868 22448
rect 28724 22160 28776 22166
rect 28724 22102 28776 22108
rect 28632 22092 28684 22098
rect 29196 22094 29224 29786
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 29552 28008 29604 28014
rect 29552 27950 29604 27956
rect 29564 27538 29592 27950
rect 29748 27538 29776 28358
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29564 26450 29592 27474
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29276 26444 29328 26450
rect 29276 26386 29328 26392
rect 29552 26444 29604 26450
rect 29552 26386 29604 26392
rect 29288 25362 29316 26386
rect 29656 26330 29684 27406
rect 29748 26994 29776 27474
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 29564 26314 29684 26330
rect 29552 26308 29684 26314
rect 29604 26302 29684 26308
rect 29552 26250 29604 26256
rect 29460 25696 29512 25702
rect 29460 25638 29512 25644
rect 29472 25362 29500 25638
rect 29564 25362 29592 26250
rect 29276 25356 29328 25362
rect 29276 25298 29328 25304
rect 29460 25356 29512 25362
rect 29460 25298 29512 25304
rect 29552 25356 29604 25362
rect 29552 25298 29604 25304
rect 29736 25356 29788 25362
rect 29736 25298 29788 25304
rect 29472 24274 29500 25298
rect 29748 24614 29776 25298
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29840 24410 29868 31844
rect 30208 31142 30236 40038
rect 30472 39976 30524 39982
rect 30576 39964 30604 40326
rect 30656 40180 30708 40186
rect 30656 40122 30708 40128
rect 30524 39936 30604 39964
rect 30472 39918 30524 39924
rect 30380 39296 30432 39302
rect 30380 39238 30432 39244
rect 30392 39030 30420 39238
rect 30380 39024 30432 39030
rect 30380 38966 30432 38972
rect 30484 38894 30512 39918
rect 30564 39568 30616 39574
rect 30564 39510 30616 39516
rect 30472 38888 30524 38894
rect 30472 38830 30524 38836
rect 30380 38752 30432 38758
rect 30380 38694 30432 38700
rect 30392 37806 30420 38694
rect 30484 38554 30512 38830
rect 30472 38548 30524 38554
rect 30472 38490 30524 38496
rect 30380 37800 30432 37806
rect 30380 37742 30432 37748
rect 30576 37466 30604 39510
rect 30564 37460 30616 37466
rect 30564 37402 30616 37408
rect 30668 36038 30696 40122
rect 30944 39930 30972 41754
rect 31128 41750 31156 42094
rect 31116 41744 31168 41750
rect 31116 41686 31168 41692
rect 31024 40928 31076 40934
rect 31024 40870 31076 40876
rect 31036 40050 31064 40870
rect 31024 40044 31076 40050
rect 31024 39986 31076 39992
rect 30944 39902 31064 39930
rect 31036 38894 31064 39902
rect 31116 39024 31168 39030
rect 31116 38966 31168 38972
rect 31024 38888 31076 38894
rect 31024 38830 31076 38836
rect 31036 38434 31064 38830
rect 31128 38554 31156 38966
rect 31116 38548 31168 38554
rect 31116 38490 31168 38496
rect 31036 38406 31156 38434
rect 30748 38208 30800 38214
rect 30748 38150 30800 38156
rect 30760 37330 30788 38150
rect 31128 38010 31156 38406
rect 31116 38004 31168 38010
rect 31116 37946 31168 37952
rect 31128 37330 31156 37946
rect 30748 37324 30800 37330
rect 30748 37266 30800 37272
rect 31116 37324 31168 37330
rect 31116 37266 31168 37272
rect 30840 36576 30892 36582
rect 30840 36518 30892 36524
rect 30748 36236 30800 36242
rect 30748 36178 30800 36184
rect 30380 36032 30432 36038
rect 30380 35974 30432 35980
rect 30656 36032 30708 36038
rect 30656 35974 30708 35980
rect 30392 35562 30420 35974
rect 30380 35556 30432 35562
rect 30380 35498 30432 35504
rect 30288 35488 30340 35494
rect 30288 35430 30340 35436
rect 30564 35488 30616 35494
rect 30564 35430 30616 35436
rect 30300 34542 30328 35430
rect 30288 34536 30340 34542
rect 30288 34478 30340 34484
rect 30472 33108 30524 33114
rect 30472 33050 30524 33056
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30392 31890 30420 32302
rect 30380 31884 30432 31890
rect 30380 31826 30432 31832
rect 30196 31136 30248 31142
rect 30196 31078 30248 31084
rect 30208 30666 30236 31078
rect 30196 30660 30248 30666
rect 30196 30602 30248 30608
rect 29920 28212 29972 28218
rect 29920 28154 29972 28160
rect 29932 28014 29960 28154
rect 29920 28008 29972 28014
rect 29920 27950 29972 27956
rect 29932 27470 29960 27950
rect 30012 27940 30064 27946
rect 30012 27882 30064 27888
rect 30024 27538 30052 27882
rect 30012 27532 30064 27538
rect 30012 27474 30064 27480
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 29932 26314 29960 27406
rect 30012 26444 30064 26450
rect 30012 26386 30064 26392
rect 29920 26308 29972 26314
rect 29920 26250 29972 26256
rect 30024 25702 30052 26386
rect 30012 25696 30064 25702
rect 30012 25638 30064 25644
rect 29828 24404 29880 24410
rect 29828 24346 29880 24352
rect 29460 24268 29512 24274
rect 29460 24210 29512 24216
rect 30208 23254 30236 30602
rect 30392 30326 30420 31826
rect 30380 30320 30432 30326
rect 30380 30262 30432 30268
rect 30380 29708 30432 29714
rect 30380 29650 30432 29656
rect 30288 29028 30340 29034
rect 30288 28970 30340 28976
rect 30300 28218 30328 28970
rect 30392 28762 30420 29650
rect 30380 28756 30432 28762
rect 30380 28698 30432 28704
rect 30288 28212 30340 28218
rect 30288 28154 30340 28160
rect 30484 27690 30512 33050
rect 30576 30598 30604 35430
rect 30656 33312 30708 33318
rect 30656 33254 30708 33260
rect 30668 32298 30696 33254
rect 30656 32292 30708 32298
rect 30656 32234 30708 32240
rect 30564 30592 30616 30598
rect 30564 30534 30616 30540
rect 30576 30258 30604 30534
rect 30656 30320 30708 30326
rect 30656 30262 30708 30268
rect 30564 30252 30616 30258
rect 30564 30194 30616 30200
rect 30668 29714 30696 30262
rect 30656 29708 30708 29714
rect 30656 29650 30708 29656
rect 30668 29306 30696 29650
rect 30656 29300 30708 29306
rect 30656 29242 30708 29248
rect 30484 27662 30604 27690
rect 30472 27532 30524 27538
rect 30472 27474 30524 27480
rect 30484 26790 30512 27474
rect 30472 26784 30524 26790
rect 30472 26726 30524 26732
rect 30484 26382 30512 26726
rect 30576 26450 30604 27662
rect 30564 26444 30616 26450
rect 30564 26386 30616 26392
rect 30472 26376 30524 26382
rect 30472 26318 30524 26324
rect 30484 25362 30512 26318
rect 30472 25356 30524 25362
rect 30472 25298 30524 25304
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 30392 24750 30420 25094
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 30576 24410 30604 26386
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30288 24336 30340 24342
rect 30288 24278 30340 24284
rect 30300 23322 30328 24278
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30196 23248 30248 23254
rect 30196 23190 30248 23196
rect 29368 22432 29420 22438
rect 29368 22374 29420 22380
rect 29380 22098 29408 22374
rect 28632 22034 28684 22040
rect 29104 22066 29224 22094
rect 29368 22092 29420 22098
rect 30300 22094 30328 23258
rect 30668 22094 30696 26318
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28368 21814 28488 21842
rect 28368 21434 28396 21814
rect 28552 21706 28580 21966
rect 28460 21678 28580 21706
rect 28460 21622 28488 21678
rect 28448 21616 28500 21622
rect 28644 21570 28672 22034
rect 28724 21956 28776 21962
rect 28724 21898 28776 21904
rect 28448 21558 28500 21564
rect 28552 21542 28672 21570
rect 28552 21486 28580 21542
rect 28448 21480 28500 21486
rect 28368 21428 28448 21434
rect 28368 21422 28500 21428
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28368 21406 28488 21422
rect 28368 21010 28396 21406
rect 28552 21146 28580 21422
rect 28540 21140 28592 21146
rect 28540 21082 28592 21088
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28736 20602 28764 21898
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28908 21888 28960 21894
rect 28908 21830 28960 21836
rect 28828 21078 28856 21830
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28368 19310 28396 19654
rect 28736 19310 28764 20334
rect 28920 19854 28948 21830
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28368 16538 28396 19246
rect 28736 18630 28764 19246
rect 28816 19168 28868 19174
rect 28816 19110 28868 19116
rect 28828 18902 28856 19110
rect 28816 18896 28868 18902
rect 28816 18838 28868 18844
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 28448 17536 28500 17542
rect 28448 17478 28500 17484
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 28460 16658 28488 17478
rect 28644 17270 28672 17478
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28448 16652 28500 16658
rect 28448 16594 28500 16600
rect 28368 16510 28488 16538
rect 28356 15428 28408 15434
rect 28356 15370 28408 15376
rect 28368 15162 28396 15370
rect 28356 15156 28408 15162
rect 28356 15098 28408 15104
rect 28460 14618 28488 16510
rect 28644 16250 28672 17206
rect 28632 16244 28684 16250
rect 28632 16186 28684 16192
rect 28736 16130 28764 18566
rect 28920 18426 28948 19314
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 28908 18420 28960 18426
rect 28908 18362 28960 18368
rect 29012 18222 29040 19246
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 28816 16992 28868 16998
rect 28816 16934 28868 16940
rect 28828 16590 28856 16934
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 28920 16658 28948 16730
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 28816 16584 28868 16590
rect 28816 16526 28868 16532
rect 28644 16102 28764 16130
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28644 14482 28672 16102
rect 29012 15178 29040 18158
rect 29104 16590 29132 22066
rect 29368 22034 29420 22040
rect 30208 22066 30328 22094
rect 30576 22066 30696 22094
rect 29460 21684 29512 21690
rect 29460 21626 29512 21632
rect 29276 17196 29328 17202
rect 29276 17138 29328 17144
rect 29288 16726 29316 17138
rect 29472 17082 29500 21626
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 29380 17054 29500 17082
rect 29276 16720 29328 16726
rect 29276 16662 29328 16668
rect 29092 16584 29144 16590
rect 29092 16526 29144 16532
rect 29276 16584 29328 16590
rect 29276 16526 29328 16532
rect 29184 16516 29236 16522
rect 29184 16458 29236 16464
rect 29196 15978 29224 16458
rect 29184 15972 29236 15978
rect 29184 15914 29236 15920
rect 29196 15570 29224 15914
rect 29288 15570 29316 16526
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29276 15564 29328 15570
rect 29276 15506 29328 15512
rect 28920 15150 29040 15178
rect 28724 15088 28776 15094
rect 28776 15036 28856 15042
rect 28724 15030 28856 15036
rect 28736 15014 28856 15030
rect 28724 14612 28776 14618
rect 28724 14554 28776 14560
rect 28632 14476 28684 14482
rect 28632 14418 28684 14424
rect 28448 14340 28500 14346
rect 28448 14282 28500 14288
rect 28460 13870 28488 14282
rect 28540 14000 28592 14006
rect 28540 13942 28592 13948
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28460 13190 28488 13806
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 28460 12306 28488 13126
rect 28448 12300 28500 12306
rect 28448 12242 28500 12248
rect 28356 12164 28408 12170
rect 28356 12106 28408 12112
rect 28368 11694 28396 12106
rect 28356 11688 28408 11694
rect 28356 11630 28408 11636
rect 28448 11688 28500 11694
rect 28448 11630 28500 11636
rect 28460 11354 28488 11630
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28552 9178 28580 13942
rect 28736 13870 28764 14554
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28540 9172 28592 9178
rect 28540 9114 28592 9120
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28368 7002 28396 8026
rect 28356 6996 28408 7002
rect 28356 6938 28408 6944
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 28356 6656 28408 6662
rect 28356 6598 28408 6604
rect 28368 6458 28396 6598
rect 28356 6452 28408 6458
rect 28356 6394 28408 6400
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 28368 5914 28396 6122
rect 28460 6118 28488 6802
rect 28644 6662 28672 12174
rect 28736 11762 28764 13806
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28724 10464 28776 10470
rect 28724 10406 28776 10412
rect 28736 6798 28764 10406
rect 28828 9382 28856 15014
rect 28920 11286 28948 15150
rect 29184 14272 29236 14278
rect 29184 14214 29236 14220
rect 29000 13932 29052 13938
rect 29000 13874 29052 13880
rect 29012 12986 29040 13874
rect 29196 13462 29224 14214
rect 29184 13456 29236 13462
rect 29184 13398 29236 13404
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 29012 11354 29040 12922
rect 29092 12912 29144 12918
rect 29092 12854 29144 12860
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 28908 11008 28960 11014
rect 28908 10950 28960 10956
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28920 8498 28948 10950
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29012 9518 29040 9998
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 29012 7750 29040 9454
rect 29104 9178 29132 12854
rect 29276 10192 29328 10198
rect 29276 10134 29328 10140
rect 29092 9172 29144 9178
rect 29092 9114 29144 9120
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 7342 29040 7686
rect 29000 7336 29052 7342
rect 29000 7278 29052 7284
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28724 6452 28776 6458
rect 28724 6394 28776 6400
rect 28448 6112 28500 6118
rect 28448 6054 28500 6060
rect 28356 5908 28408 5914
rect 28356 5850 28408 5856
rect 28460 5778 28488 6054
rect 28448 5772 28500 5778
rect 28448 5714 28500 5720
rect 28736 5370 28764 6394
rect 28724 5364 28776 5370
rect 28724 5306 28776 5312
rect 29012 4690 29040 7278
rect 29104 6866 29132 8774
rect 29288 7546 29316 10134
rect 29380 9042 29408 17054
rect 29460 16720 29512 16726
rect 29460 16662 29512 16668
rect 29472 16250 29500 16662
rect 29460 16244 29512 16250
rect 29460 16186 29512 16192
rect 29564 16130 29592 21082
rect 30208 20534 30236 22066
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 30196 20528 30248 20534
rect 30196 20470 30248 20476
rect 30300 20398 30328 21354
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 29736 19168 29788 19174
rect 29736 19110 29788 19116
rect 29644 18828 29696 18834
rect 29748 18816 29776 19110
rect 29696 18788 29776 18816
rect 29644 18770 29696 18776
rect 29748 18222 29776 18788
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29748 17678 29776 18158
rect 29932 17814 29960 19654
rect 30392 19174 30420 20878
rect 30484 20466 30512 21286
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 30472 20324 30524 20330
rect 30472 20266 30524 20272
rect 30484 19378 30512 20266
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30484 18986 30512 19314
rect 30392 18958 30512 18986
rect 30288 18148 30340 18154
rect 30288 18090 30340 18096
rect 29920 17808 29972 17814
rect 29920 17750 29972 17756
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29656 16658 29684 17138
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 29472 16102 29592 16130
rect 29368 9036 29420 9042
rect 29368 8978 29420 8984
rect 29368 8900 29420 8906
rect 29368 8842 29420 8848
rect 29380 8022 29408 8842
rect 29472 8634 29500 16102
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29564 14550 29592 15438
rect 29552 14544 29604 14550
rect 29552 14486 29604 14492
rect 29656 14482 29684 16594
rect 29748 14958 29776 17614
rect 30104 17332 30156 17338
rect 30104 17274 30156 17280
rect 30116 17134 30144 17274
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 29840 16590 29868 17070
rect 30024 16810 30052 17070
rect 30024 16782 30144 16810
rect 30208 16794 30236 17682
rect 30300 17338 30328 18090
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 30024 16114 30052 16594
rect 30116 16250 30144 16782
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 30300 16658 30328 17138
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30104 16244 30156 16250
rect 30104 16186 30156 16192
rect 30012 16108 30064 16114
rect 30012 16050 30064 16056
rect 30024 15162 30052 16050
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29644 14476 29696 14482
rect 29644 14418 29696 14424
rect 29656 12782 29684 14418
rect 29748 13394 29776 14894
rect 30024 14550 30052 15098
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 29840 14006 29868 14418
rect 30116 14414 30144 16186
rect 30392 15042 30420 18958
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30484 17134 30512 18022
rect 30576 17218 30604 22066
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30668 20466 30696 21490
rect 30760 21146 30788 36178
rect 30852 31482 30880 36518
rect 30932 35080 30984 35086
rect 30932 35022 30984 35028
rect 30944 34610 30972 35022
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30944 32434 30972 34546
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 31220 31754 31248 42706
rect 31300 39976 31352 39982
rect 31300 39918 31352 39924
rect 31312 39098 31340 39918
rect 31300 39092 31352 39098
rect 31300 39034 31352 39040
rect 31484 31884 31536 31890
rect 31484 31826 31536 31832
rect 31220 31726 31340 31754
rect 30840 31476 30892 31482
rect 30840 31418 30892 31424
rect 30852 27402 30880 31418
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 31036 30734 31064 31078
rect 31024 30728 31076 30734
rect 31024 30670 31076 30676
rect 30840 27396 30892 27402
rect 30840 27338 30892 27344
rect 30932 27328 30984 27334
rect 30932 27270 30984 27276
rect 30944 26926 30972 27270
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 31036 26858 31064 30670
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 31220 28626 31248 29106
rect 31208 28620 31260 28626
rect 31208 28562 31260 28568
rect 31116 28008 31168 28014
rect 31116 27950 31168 27956
rect 31128 27674 31156 27950
rect 31116 27668 31168 27674
rect 31116 27610 31168 27616
rect 31220 26994 31248 28562
rect 31312 27538 31340 31726
rect 31300 27532 31352 27538
rect 31300 27474 31352 27480
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31024 26852 31076 26858
rect 31024 26794 31076 26800
rect 31036 26450 31064 26794
rect 31024 26444 31076 26450
rect 31024 26386 31076 26392
rect 31024 26308 31076 26314
rect 31024 26250 31076 26256
rect 31036 25838 31064 26250
rect 31220 25838 31248 26930
rect 31024 25832 31076 25838
rect 31024 25774 31076 25780
rect 31208 25832 31260 25838
rect 31208 25774 31260 25780
rect 31220 24818 31248 25774
rect 31312 25362 31340 27474
rect 31300 25356 31352 25362
rect 31300 25298 31352 25304
rect 31208 24812 31260 24818
rect 31208 24754 31260 24760
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 30852 21486 30880 24346
rect 31312 24342 31340 25298
rect 31300 24336 31352 24342
rect 31300 24278 31352 24284
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 31024 24132 31076 24138
rect 31024 24074 31076 24080
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30944 22642 30972 23598
rect 31036 23186 31064 24074
rect 31128 23322 31156 24210
rect 31116 23316 31168 23322
rect 31116 23258 31168 23264
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 31300 23180 31352 23186
rect 31300 23122 31352 23128
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30840 21480 30892 21486
rect 30840 21422 30892 21428
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 30944 21026 30972 22578
rect 31312 22098 31340 23122
rect 31300 22092 31352 22098
rect 31300 22034 31352 22040
rect 31312 21690 31340 22034
rect 31300 21684 31352 21690
rect 31300 21626 31352 21632
rect 31024 21616 31076 21622
rect 31024 21558 31076 21564
rect 30852 20998 30972 21026
rect 31036 21010 31064 21558
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31208 21480 31260 21486
rect 31128 21428 31208 21434
rect 31128 21422 31260 21428
rect 31128 21406 31248 21422
rect 31024 21004 31076 21010
rect 30852 20942 30880 20998
rect 31024 20946 31076 20952
rect 30840 20936 30892 20942
rect 30840 20878 30892 20884
rect 30932 20936 30984 20942
rect 30932 20878 30984 20884
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30668 19242 30696 20402
rect 30944 20398 30972 20878
rect 30932 20392 30984 20398
rect 30932 20334 30984 20340
rect 31036 20074 31064 20946
rect 31128 20942 31156 21406
rect 31208 21344 31260 21350
rect 31208 21286 31260 21292
rect 31220 21010 31248 21286
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 30944 20046 31064 20074
rect 31128 20058 31156 20878
rect 31116 20052 31168 20058
rect 30748 19916 30800 19922
rect 30748 19858 30800 19864
rect 30760 19514 30788 19858
rect 30748 19508 30800 19514
rect 30748 19450 30800 19456
rect 30656 19236 30708 19242
rect 30656 19178 30708 19184
rect 30668 18970 30696 19178
rect 30656 18964 30708 18970
rect 30656 18906 30708 18912
rect 30944 17882 30972 20046
rect 31116 19994 31168 20000
rect 31404 19990 31432 21490
rect 31024 19984 31076 19990
rect 31024 19926 31076 19932
rect 31392 19984 31444 19990
rect 31392 19926 31444 19932
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 30932 17876 30984 17882
rect 30932 17818 30984 17824
rect 30656 17536 30708 17542
rect 30656 17478 30708 17484
rect 30668 17338 30696 17478
rect 30656 17332 30708 17338
rect 30656 17274 30708 17280
rect 30576 17190 30788 17218
rect 30472 17128 30524 17134
rect 30472 17070 30524 17076
rect 30656 17128 30708 17134
rect 30656 17070 30708 17076
rect 30564 16788 30616 16794
rect 30564 16730 30616 16736
rect 30472 16720 30524 16726
rect 30472 16662 30524 16668
rect 30300 15014 30420 15042
rect 30300 14890 30328 15014
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30380 14884 30432 14890
rect 30380 14826 30432 14832
rect 30300 14498 30328 14826
rect 30392 14618 30420 14826
rect 30380 14612 30432 14618
rect 30380 14554 30432 14560
rect 30300 14470 30420 14498
rect 30484 14482 30512 16662
rect 30576 15706 30604 16730
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30564 14816 30616 14822
rect 30564 14758 30616 14764
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29920 14272 29972 14278
rect 29920 14214 29972 14220
rect 29828 14000 29880 14006
rect 29828 13942 29880 13948
rect 29736 13388 29788 13394
rect 29736 13330 29788 13336
rect 29932 12782 29960 14214
rect 30116 13852 30144 14350
rect 30196 14000 30248 14006
rect 30196 13942 30248 13948
rect 30024 13824 30144 13852
rect 30024 12850 30052 13824
rect 30104 13184 30156 13190
rect 30104 13126 30156 13132
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29920 12776 29972 12782
rect 29920 12718 29972 12724
rect 29564 12238 29592 12718
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 29564 11014 29592 12174
rect 29656 12170 29684 12718
rect 29932 12434 29960 12718
rect 29840 12406 29960 12434
rect 29736 12300 29788 12306
rect 29736 12242 29788 12248
rect 29644 12164 29696 12170
rect 29644 12106 29696 12112
rect 29748 11694 29776 12242
rect 29840 11898 29868 12406
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 29840 11762 29868 11834
rect 30024 11762 30052 12786
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 30012 11756 30064 11762
rect 30012 11698 30064 11704
rect 29736 11688 29788 11694
rect 29736 11630 29788 11636
rect 29644 11552 29696 11558
rect 29644 11494 29696 11500
rect 29552 11008 29604 11014
rect 29552 10950 29604 10956
rect 29564 10606 29592 10950
rect 29656 10606 29684 11494
rect 29748 10810 29776 11630
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29644 10600 29696 10606
rect 29644 10542 29696 10548
rect 29564 10062 29592 10542
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 29460 8628 29512 8634
rect 29460 8570 29512 8576
rect 29368 8016 29420 8022
rect 29368 7958 29420 7964
rect 30024 7546 30052 9658
rect 30116 9654 30144 13126
rect 30208 12782 30236 13942
rect 30392 13870 30420 14470
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30472 13864 30524 13870
rect 30472 13806 30524 13812
rect 30392 13530 30420 13806
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 12986 30328 13194
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30196 12640 30248 12646
rect 30196 12582 30248 12588
rect 30208 12374 30236 12582
rect 30300 12442 30328 12922
rect 30380 12776 30432 12782
rect 30380 12718 30432 12724
rect 30392 12442 30420 12718
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30380 12436 30432 12442
rect 30380 12378 30432 12384
rect 30196 12368 30248 12374
rect 30196 12310 30248 12316
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 30300 10198 30328 11494
rect 30484 11218 30512 13806
rect 30576 13682 30604 14758
rect 30668 13870 30696 17070
rect 30760 16674 30788 17190
rect 30852 16794 30880 17818
rect 30944 17202 30972 17818
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 31036 16794 31064 19926
rect 31300 19916 31352 19922
rect 31300 19858 31352 19864
rect 31312 18086 31340 19858
rect 31300 18080 31352 18086
rect 31300 18022 31352 18028
rect 30840 16788 30892 16794
rect 30840 16730 30892 16736
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 30760 16646 31340 16674
rect 31404 16658 31432 19926
rect 30932 15904 30984 15910
rect 30932 15846 30984 15852
rect 30944 15638 30972 15846
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 30932 15632 30984 15638
rect 30932 15574 30984 15580
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30748 14408 30800 14414
rect 30748 14350 30800 14356
rect 30760 14074 30788 14350
rect 30748 14068 30800 14074
rect 30748 14010 30800 14016
rect 30852 14006 30880 15302
rect 30840 14000 30892 14006
rect 30840 13942 30892 13948
rect 30944 13938 30972 15574
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30656 13864 30708 13870
rect 30656 13806 30708 13812
rect 30576 13654 30696 13682
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30472 11212 30524 11218
rect 30472 11154 30524 11160
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 30012 7540 30064 7546
rect 30012 7482 30064 7488
rect 29288 6866 29316 7482
rect 29092 6860 29144 6866
rect 29092 6802 29144 6808
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 29288 6458 29316 6802
rect 29276 6452 29328 6458
rect 29276 6394 29328 6400
rect 29288 5914 29316 6394
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 30024 5370 30052 7482
rect 30116 6458 30144 9590
rect 30380 9036 30432 9042
rect 30380 8978 30432 8984
rect 30392 8362 30420 8978
rect 30380 8356 30432 8362
rect 30380 8298 30432 8304
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 30104 5568 30156 5574
rect 30104 5510 30156 5516
rect 30012 5364 30064 5370
rect 30012 5306 30064 5312
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 28368 4078 28396 4422
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 27804 3732 27856 3738
rect 27804 3674 27856 3680
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 28368 3602 28396 4014
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27804 3596 27856 3602
rect 27804 3538 27856 3544
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 27344 2916 27396 2922
rect 27344 2858 27396 2864
rect 27356 2514 27384 2858
rect 27344 2508 27396 2514
rect 27344 2450 27396 2456
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 27356 1834 27384 2246
rect 27540 1834 27568 3538
rect 27816 3194 27844 3538
rect 28736 3194 28764 4082
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29000 4004 29052 4010
rect 29000 3946 29052 3952
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 28632 3052 28684 3058
rect 28632 2994 28684 3000
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 28092 2514 28120 2790
rect 28080 2508 28132 2514
rect 28080 2450 28132 2456
rect 27344 1828 27396 1834
rect 27344 1770 27396 1776
rect 27528 1828 27580 1834
rect 27528 1770 27580 1776
rect 27540 1222 27568 1770
rect 28184 1426 28212 2790
rect 28552 2650 28580 2926
rect 28540 2644 28592 2650
rect 28540 2586 28592 2592
rect 28264 2508 28316 2514
rect 28264 2450 28316 2456
rect 28276 2378 28304 2450
rect 28644 2446 28672 2994
rect 28828 2854 28856 3538
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28816 2848 28868 2854
rect 28816 2790 28868 2796
rect 28816 2508 28868 2514
rect 28920 2496 28948 2926
rect 28868 2468 28948 2496
rect 28816 2450 28868 2456
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 28264 2372 28316 2378
rect 28264 2314 28316 2320
rect 28828 2106 28856 2450
rect 28816 2100 28868 2106
rect 28816 2042 28868 2048
rect 29012 1834 29040 3946
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29000 1828 29052 1834
rect 29000 1770 29052 1776
rect 29012 1562 29040 1770
rect 29000 1556 29052 1562
rect 29000 1498 29052 1504
rect 28172 1420 28224 1426
rect 28172 1362 28224 1368
rect 27528 1216 27580 1222
rect 27528 1158 27580 1164
rect 29012 1018 29040 1498
rect 29104 1494 29132 2926
rect 29184 2916 29236 2922
rect 29184 2858 29236 2864
rect 29196 2378 29224 2858
rect 29564 2650 29592 4014
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 29184 2372 29236 2378
rect 29184 2314 29236 2320
rect 30024 2106 30052 4762
rect 30116 3194 30144 5510
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 30300 3602 30328 5238
rect 30392 4078 30420 8298
rect 30576 5914 30604 13466
rect 30668 11354 30696 13654
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30748 13184 30800 13190
rect 30748 13126 30800 13132
rect 30760 11898 30788 13126
rect 30852 12782 30880 13262
rect 30840 12776 30892 12782
rect 30892 12736 30972 12764
rect 30840 12718 30892 12724
rect 30840 12640 30892 12646
rect 30840 12582 30892 12588
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 30852 11762 30880 12582
rect 30840 11756 30892 11762
rect 30840 11698 30892 11704
rect 30944 11694 30972 12736
rect 31036 12646 31064 15642
rect 31208 15360 31260 15366
rect 31208 15302 31260 15308
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 30932 11688 30984 11694
rect 30932 11630 30984 11636
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30944 10266 30972 11630
rect 30748 10260 30800 10266
rect 30748 10202 30800 10208
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 30760 8090 30788 10202
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 30852 7478 30880 8774
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 30840 7472 30892 7478
rect 30840 7414 30892 7420
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30576 4826 30604 5850
rect 30656 5364 30708 5370
rect 30656 5306 30708 5312
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30472 4752 30524 4758
rect 30472 4694 30524 4700
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30104 3188 30156 3194
rect 30104 3130 30156 3136
rect 30104 2372 30156 2378
rect 30104 2314 30156 2320
rect 30012 2100 30064 2106
rect 30012 2042 30064 2048
rect 30024 1562 30052 2042
rect 30116 1834 30144 2314
rect 30104 1828 30156 1834
rect 30104 1770 30156 1776
rect 30012 1556 30064 1562
rect 30012 1498 30064 1504
rect 29092 1488 29144 1494
rect 29092 1430 29144 1436
rect 29000 1012 29052 1018
rect 29000 954 29052 960
rect 27160 876 27212 882
rect 27160 818 27212 824
rect 25780 808 25832 814
rect 25780 750 25832 756
rect 26148 808 26200 814
rect 26148 750 26200 756
rect 26240 808 26292 814
rect 26240 750 26292 756
rect 26700 808 26752 814
rect 30392 800 30420 3674
rect 30484 3670 30512 4694
rect 30668 4146 30696 5306
rect 30656 4140 30708 4146
rect 30656 4082 30708 4088
rect 30564 4072 30616 4078
rect 30564 4014 30616 4020
rect 30576 3738 30604 4014
rect 30564 3732 30616 3738
rect 30564 3674 30616 3680
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30760 2774 30788 6734
rect 30944 4146 30972 8434
rect 31036 6610 31064 12582
rect 31128 11694 31156 14418
rect 31220 14414 31248 15302
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 31208 13388 31260 13394
rect 31208 13330 31260 13336
rect 31116 11688 31168 11694
rect 31116 11630 31168 11636
rect 31116 11552 31168 11558
rect 31116 11494 31168 11500
rect 31128 11218 31156 11494
rect 31116 11212 31168 11218
rect 31116 11154 31168 11160
rect 31116 7336 31168 7342
rect 31116 7278 31168 7284
rect 31128 7002 31156 7278
rect 31116 6996 31168 7002
rect 31116 6938 31168 6944
rect 31036 6582 31156 6610
rect 31024 6452 31076 6458
rect 31024 6394 31076 6400
rect 31036 4826 31064 6394
rect 31128 5914 31156 6582
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 31128 5370 31156 5850
rect 31116 5364 31168 5370
rect 31116 5306 31168 5312
rect 31024 4820 31076 4826
rect 31024 4762 31076 4768
rect 31220 4758 31248 13330
rect 31312 6866 31340 16646
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31496 14618 31524 31826
rect 31588 21554 31616 45970
rect 31668 34060 31720 34066
rect 31668 34002 31720 34008
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31576 21412 31628 21418
rect 31576 21354 31628 21360
rect 31484 14612 31536 14618
rect 31484 14554 31536 14560
rect 31300 6860 31352 6866
rect 31300 6802 31352 6808
rect 31312 5166 31340 6802
rect 31588 6458 31616 21354
rect 31680 20602 31708 34002
rect 31668 20596 31720 20602
rect 31668 20538 31720 20544
rect 31576 6452 31628 6458
rect 31576 6394 31628 6400
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 31208 4752 31260 4758
rect 31208 4694 31260 4700
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30484 2746 30788 2774
rect 30484 1426 30512 2746
rect 30944 2650 30972 4082
rect 31312 3194 31340 5102
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 31036 2530 31064 3130
rect 30944 2502 31064 2530
rect 30944 1766 30972 2502
rect 30932 1760 30984 1766
rect 30932 1702 30984 1708
rect 30472 1420 30524 1426
rect 30472 1362 30524 1368
rect 30944 814 30972 1702
rect 30932 808 30984 814
rect 26700 750 26752 756
rect 25688 672 25740 678
rect 25688 614 25740 620
rect 26148 672 26200 678
rect 26148 614 26200 620
rect 26160 474 26188 614
rect 24952 468 25004 474
rect 24952 410 25004 416
rect 26148 468 26200 474
rect 26148 410 26200 416
rect 26712 406 26740 750
rect 26700 400 26752 406
rect 26700 342 26752 348
rect 30378 0 30434 800
rect 30932 750 30984 756
<< via2 >>
rect 11259 48442 11315 48444
rect 11339 48442 11395 48444
rect 11419 48442 11475 48444
rect 11499 48442 11555 48444
rect 11259 48390 11305 48442
rect 11305 48390 11315 48442
rect 11339 48390 11369 48442
rect 11369 48390 11381 48442
rect 11381 48390 11395 48442
rect 11419 48390 11433 48442
rect 11433 48390 11445 48442
rect 11445 48390 11475 48442
rect 11499 48390 11509 48442
rect 11509 48390 11555 48442
rect 11259 48388 11315 48390
rect 11339 48388 11395 48390
rect 11419 48388 11475 48390
rect 11499 48388 11555 48390
rect 21563 48442 21619 48444
rect 21643 48442 21699 48444
rect 21723 48442 21779 48444
rect 21803 48442 21859 48444
rect 21563 48390 21609 48442
rect 21609 48390 21619 48442
rect 21643 48390 21673 48442
rect 21673 48390 21685 48442
rect 21685 48390 21699 48442
rect 21723 48390 21737 48442
rect 21737 48390 21749 48442
rect 21749 48390 21779 48442
rect 21803 48390 21813 48442
rect 21813 48390 21859 48442
rect 21563 48388 21619 48390
rect 21643 48388 21699 48390
rect 21723 48388 21779 48390
rect 21803 48388 21859 48390
rect 6108 47898 6164 47900
rect 6188 47898 6244 47900
rect 6268 47898 6324 47900
rect 6348 47898 6404 47900
rect 6108 47846 6154 47898
rect 6154 47846 6164 47898
rect 6188 47846 6218 47898
rect 6218 47846 6230 47898
rect 6230 47846 6244 47898
rect 6268 47846 6282 47898
rect 6282 47846 6294 47898
rect 6294 47846 6324 47898
rect 6348 47846 6358 47898
rect 6358 47846 6404 47898
rect 6108 47844 6164 47846
rect 6188 47844 6244 47846
rect 6268 47844 6324 47846
rect 6348 47844 6404 47846
rect 6108 46810 6164 46812
rect 6188 46810 6244 46812
rect 6268 46810 6324 46812
rect 6348 46810 6404 46812
rect 6108 46758 6154 46810
rect 6154 46758 6164 46810
rect 6188 46758 6218 46810
rect 6218 46758 6230 46810
rect 6230 46758 6244 46810
rect 6268 46758 6282 46810
rect 6282 46758 6294 46810
rect 6294 46758 6324 46810
rect 6348 46758 6358 46810
rect 6358 46758 6404 46810
rect 6108 46756 6164 46758
rect 6188 46756 6244 46758
rect 6268 46756 6324 46758
rect 6348 46756 6404 46758
rect 6108 45722 6164 45724
rect 6188 45722 6244 45724
rect 6268 45722 6324 45724
rect 6348 45722 6404 45724
rect 6108 45670 6154 45722
rect 6154 45670 6164 45722
rect 6188 45670 6218 45722
rect 6218 45670 6230 45722
rect 6230 45670 6244 45722
rect 6268 45670 6282 45722
rect 6282 45670 6294 45722
rect 6294 45670 6324 45722
rect 6348 45670 6358 45722
rect 6358 45670 6404 45722
rect 6108 45668 6164 45670
rect 6188 45668 6244 45670
rect 6268 45668 6324 45670
rect 6348 45668 6404 45670
rect 6108 44634 6164 44636
rect 6188 44634 6244 44636
rect 6268 44634 6324 44636
rect 6348 44634 6404 44636
rect 6108 44582 6154 44634
rect 6154 44582 6164 44634
rect 6188 44582 6218 44634
rect 6218 44582 6230 44634
rect 6230 44582 6244 44634
rect 6268 44582 6282 44634
rect 6282 44582 6294 44634
rect 6294 44582 6324 44634
rect 6348 44582 6358 44634
rect 6358 44582 6404 44634
rect 6108 44580 6164 44582
rect 6188 44580 6244 44582
rect 6268 44580 6324 44582
rect 6348 44580 6404 44582
rect 6108 43546 6164 43548
rect 6188 43546 6244 43548
rect 6268 43546 6324 43548
rect 6348 43546 6404 43548
rect 6108 43494 6154 43546
rect 6154 43494 6164 43546
rect 6188 43494 6218 43546
rect 6218 43494 6230 43546
rect 6230 43494 6244 43546
rect 6268 43494 6282 43546
rect 6282 43494 6294 43546
rect 6294 43494 6324 43546
rect 6348 43494 6358 43546
rect 6358 43494 6404 43546
rect 6108 43492 6164 43494
rect 6188 43492 6244 43494
rect 6268 43492 6324 43494
rect 6348 43492 6404 43494
rect 6108 42458 6164 42460
rect 6188 42458 6244 42460
rect 6268 42458 6324 42460
rect 6348 42458 6404 42460
rect 6108 42406 6154 42458
rect 6154 42406 6164 42458
rect 6188 42406 6218 42458
rect 6218 42406 6230 42458
rect 6230 42406 6244 42458
rect 6268 42406 6282 42458
rect 6282 42406 6294 42458
rect 6294 42406 6324 42458
rect 6348 42406 6358 42458
rect 6358 42406 6404 42458
rect 6108 42404 6164 42406
rect 6188 42404 6244 42406
rect 6268 42404 6324 42406
rect 6348 42404 6404 42406
rect 6108 41370 6164 41372
rect 6188 41370 6244 41372
rect 6268 41370 6324 41372
rect 6348 41370 6404 41372
rect 6108 41318 6154 41370
rect 6154 41318 6164 41370
rect 6188 41318 6218 41370
rect 6218 41318 6230 41370
rect 6230 41318 6244 41370
rect 6268 41318 6282 41370
rect 6282 41318 6294 41370
rect 6294 41318 6324 41370
rect 6348 41318 6358 41370
rect 6358 41318 6404 41370
rect 6108 41316 6164 41318
rect 6188 41316 6244 41318
rect 6268 41316 6324 41318
rect 6348 41316 6404 41318
rect 6108 40282 6164 40284
rect 6188 40282 6244 40284
rect 6268 40282 6324 40284
rect 6348 40282 6404 40284
rect 6108 40230 6154 40282
rect 6154 40230 6164 40282
rect 6188 40230 6218 40282
rect 6218 40230 6230 40282
rect 6230 40230 6244 40282
rect 6268 40230 6282 40282
rect 6282 40230 6294 40282
rect 6294 40230 6324 40282
rect 6348 40230 6358 40282
rect 6358 40230 6404 40282
rect 6108 40228 6164 40230
rect 6188 40228 6244 40230
rect 6268 40228 6324 40230
rect 6348 40228 6404 40230
rect 6108 39194 6164 39196
rect 6188 39194 6244 39196
rect 6268 39194 6324 39196
rect 6348 39194 6404 39196
rect 6108 39142 6154 39194
rect 6154 39142 6164 39194
rect 6188 39142 6218 39194
rect 6218 39142 6230 39194
rect 6230 39142 6244 39194
rect 6268 39142 6282 39194
rect 6282 39142 6294 39194
rect 6294 39142 6324 39194
rect 6348 39142 6358 39194
rect 6358 39142 6404 39194
rect 6108 39140 6164 39142
rect 6188 39140 6244 39142
rect 6268 39140 6324 39142
rect 6348 39140 6404 39142
rect 6108 38106 6164 38108
rect 6188 38106 6244 38108
rect 6268 38106 6324 38108
rect 6348 38106 6404 38108
rect 6108 38054 6154 38106
rect 6154 38054 6164 38106
rect 6188 38054 6218 38106
rect 6218 38054 6230 38106
rect 6230 38054 6244 38106
rect 6268 38054 6282 38106
rect 6282 38054 6294 38106
rect 6294 38054 6324 38106
rect 6348 38054 6358 38106
rect 6358 38054 6404 38106
rect 6108 38052 6164 38054
rect 6188 38052 6244 38054
rect 6268 38052 6324 38054
rect 6348 38052 6404 38054
rect 6108 37018 6164 37020
rect 6188 37018 6244 37020
rect 6268 37018 6324 37020
rect 6348 37018 6404 37020
rect 6108 36966 6154 37018
rect 6154 36966 6164 37018
rect 6188 36966 6218 37018
rect 6218 36966 6230 37018
rect 6230 36966 6244 37018
rect 6268 36966 6282 37018
rect 6282 36966 6294 37018
rect 6294 36966 6324 37018
rect 6348 36966 6358 37018
rect 6358 36966 6404 37018
rect 6108 36964 6164 36966
rect 6188 36964 6244 36966
rect 6268 36964 6324 36966
rect 6348 36964 6404 36966
rect 6108 35930 6164 35932
rect 6188 35930 6244 35932
rect 6268 35930 6324 35932
rect 6348 35930 6404 35932
rect 6108 35878 6154 35930
rect 6154 35878 6164 35930
rect 6188 35878 6218 35930
rect 6218 35878 6230 35930
rect 6230 35878 6244 35930
rect 6268 35878 6282 35930
rect 6282 35878 6294 35930
rect 6294 35878 6324 35930
rect 6348 35878 6358 35930
rect 6358 35878 6404 35930
rect 6108 35876 6164 35878
rect 6188 35876 6244 35878
rect 6268 35876 6324 35878
rect 6348 35876 6404 35878
rect 6108 34842 6164 34844
rect 6188 34842 6244 34844
rect 6268 34842 6324 34844
rect 6348 34842 6404 34844
rect 6108 34790 6154 34842
rect 6154 34790 6164 34842
rect 6188 34790 6218 34842
rect 6218 34790 6230 34842
rect 6230 34790 6244 34842
rect 6268 34790 6282 34842
rect 6282 34790 6294 34842
rect 6294 34790 6324 34842
rect 6348 34790 6358 34842
rect 6358 34790 6404 34842
rect 6108 34788 6164 34790
rect 6188 34788 6244 34790
rect 6268 34788 6324 34790
rect 6348 34788 6404 34790
rect 6108 33754 6164 33756
rect 6188 33754 6244 33756
rect 6268 33754 6324 33756
rect 6348 33754 6404 33756
rect 6108 33702 6154 33754
rect 6154 33702 6164 33754
rect 6188 33702 6218 33754
rect 6218 33702 6230 33754
rect 6230 33702 6244 33754
rect 6268 33702 6282 33754
rect 6282 33702 6294 33754
rect 6294 33702 6324 33754
rect 6348 33702 6358 33754
rect 6358 33702 6404 33754
rect 6108 33700 6164 33702
rect 6188 33700 6244 33702
rect 6268 33700 6324 33702
rect 6348 33700 6404 33702
rect 6108 32666 6164 32668
rect 6188 32666 6244 32668
rect 6268 32666 6324 32668
rect 6348 32666 6404 32668
rect 6108 32614 6154 32666
rect 6154 32614 6164 32666
rect 6188 32614 6218 32666
rect 6218 32614 6230 32666
rect 6230 32614 6244 32666
rect 6268 32614 6282 32666
rect 6282 32614 6294 32666
rect 6294 32614 6324 32666
rect 6348 32614 6358 32666
rect 6358 32614 6404 32666
rect 6108 32612 6164 32614
rect 6188 32612 6244 32614
rect 6268 32612 6324 32614
rect 6348 32612 6404 32614
rect 6108 31578 6164 31580
rect 6188 31578 6244 31580
rect 6268 31578 6324 31580
rect 6348 31578 6404 31580
rect 6108 31526 6154 31578
rect 6154 31526 6164 31578
rect 6188 31526 6218 31578
rect 6218 31526 6230 31578
rect 6230 31526 6244 31578
rect 6268 31526 6282 31578
rect 6282 31526 6294 31578
rect 6294 31526 6324 31578
rect 6348 31526 6358 31578
rect 6358 31526 6404 31578
rect 6108 31524 6164 31526
rect 6188 31524 6244 31526
rect 6268 31524 6324 31526
rect 6348 31524 6404 31526
rect 6108 30490 6164 30492
rect 6188 30490 6244 30492
rect 6268 30490 6324 30492
rect 6348 30490 6404 30492
rect 6108 30438 6154 30490
rect 6154 30438 6164 30490
rect 6188 30438 6218 30490
rect 6218 30438 6230 30490
rect 6230 30438 6244 30490
rect 6268 30438 6282 30490
rect 6282 30438 6294 30490
rect 6294 30438 6324 30490
rect 6348 30438 6358 30490
rect 6358 30438 6404 30490
rect 6108 30436 6164 30438
rect 6188 30436 6244 30438
rect 6268 30436 6324 30438
rect 6348 30436 6404 30438
rect 6108 29402 6164 29404
rect 6188 29402 6244 29404
rect 6268 29402 6324 29404
rect 6348 29402 6404 29404
rect 6108 29350 6154 29402
rect 6154 29350 6164 29402
rect 6188 29350 6218 29402
rect 6218 29350 6230 29402
rect 6230 29350 6244 29402
rect 6268 29350 6282 29402
rect 6282 29350 6294 29402
rect 6294 29350 6324 29402
rect 6348 29350 6358 29402
rect 6358 29350 6404 29402
rect 6108 29348 6164 29350
rect 6188 29348 6244 29350
rect 6268 29348 6324 29350
rect 6348 29348 6404 29350
rect 6108 28314 6164 28316
rect 6188 28314 6244 28316
rect 6268 28314 6324 28316
rect 6348 28314 6404 28316
rect 6108 28262 6154 28314
rect 6154 28262 6164 28314
rect 6188 28262 6218 28314
rect 6218 28262 6230 28314
rect 6230 28262 6244 28314
rect 6268 28262 6282 28314
rect 6282 28262 6294 28314
rect 6294 28262 6324 28314
rect 6348 28262 6358 28314
rect 6358 28262 6404 28314
rect 6108 28260 6164 28262
rect 6188 28260 6244 28262
rect 6268 28260 6324 28262
rect 6348 28260 6404 28262
rect 6108 27226 6164 27228
rect 6188 27226 6244 27228
rect 6268 27226 6324 27228
rect 6348 27226 6404 27228
rect 6108 27174 6154 27226
rect 6154 27174 6164 27226
rect 6188 27174 6218 27226
rect 6218 27174 6230 27226
rect 6230 27174 6244 27226
rect 6268 27174 6282 27226
rect 6282 27174 6294 27226
rect 6294 27174 6324 27226
rect 6348 27174 6358 27226
rect 6358 27174 6404 27226
rect 6108 27172 6164 27174
rect 6188 27172 6244 27174
rect 6268 27172 6324 27174
rect 6348 27172 6404 27174
rect 6108 26138 6164 26140
rect 6188 26138 6244 26140
rect 6268 26138 6324 26140
rect 6348 26138 6404 26140
rect 6108 26086 6154 26138
rect 6154 26086 6164 26138
rect 6188 26086 6218 26138
rect 6218 26086 6230 26138
rect 6230 26086 6244 26138
rect 6268 26086 6282 26138
rect 6282 26086 6294 26138
rect 6294 26086 6324 26138
rect 6348 26086 6358 26138
rect 6358 26086 6404 26138
rect 6108 26084 6164 26086
rect 6188 26084 6244 26086
rect 6268 26084 6324 26086
rect 6348 26084 6404 26086
rect 6108 25050 6164 25052
rect 6188 25050 6244 25052
rect 6268 25050 6324 25052
rect 6348 25050 6404 25052
rect 6108 24998 6154 25050
rect 6154 24998 6164 25050
rect 6188 24998 6218 25050
rect 6218 24998 6230 25050
rect 6230 24998 6244 25050
rect 6268 24998 6282 25050
rect 6282 24998 6294 25050
rect 6294 24998 6324 25050
rect 6348 24998 6358 25050
rect 6358 24998 6404 25050
rect 6108 24996 6164 24998
rect 6188 24996 6244 24998
rect 6268 24996 6324 24998
rect 6348 24996 6404 24998
rect 6108 23962 6164 23964
rect 6188 23962 6244 23964
rect 6268 23962 6324 23964
rect 6348 23962 6404 23964
rect 6108 23910 6154 23962
rect 6154 23910 6164 23962
rect 6188 23910 6218 23962
rect 6218 23910 6230 23962
rect 6230 23910 6244 23962
rect 6268 23910 6282 23962
rect 6282 23910 6294 23962
rect 6294 23910 6324 23962
rect 6348 23910 6358 23962
rect 6358 23910 6404 23962
rect 6108 23908 6164 23910
rect 6188 23908 6244 23910
rect 6268 23908 6324 23910
rect 6348 23908 6404 23910
rect 6108 22874 6164 22876
rect 6188 22874 6244 22876
rect 6268 22874 6324 22876
rect 6348 22874 6404 22876
rect 6108 22822 6154 22874
rect 6154 22822 6164 22874
rect 6188 22822 6218 22874
rect 6218 22822 6230 22874
rect 6230 22822 6244 22874
rect 6268 22822 6282 22874
rect 6282 22822 6294 22874
rect 6294 22822 6324 22874
rect 6348 22822 6358 22874
rect 6358 22822 6404 22874
rect 6108 22820 6164 22822
rect 6188 22820 6244 22822
rect 6268 22820 6324 22822
rect 6348 22820 6404 22822
rect 6108 21786 6164 21788
rect 6188 21786 6244 21788
rect 6268 21786 6324 21788
rect 6348 21786 6404 21788
rect 6108 21734 6154 21786
rect 6154 21734 6164 21786
rect 6188 21734 6218 21786
rect 6218 21734 6230 21786
rect 6230 21734 6244 21786
rect 6268 21734 6282 21786
rect 6282 21734 6294 21786
rect 6294 21734 6324 21786
rect 6348 21734 6358 21786
rect 6358 21734 6404 21786
rect 6108 21732 6164 21734
rect 6188 21732 6244 21734
rect 6268 21732 6324 21734
rect 6348 21732 6404 21734
rect 6108 20698 6164 20700
rect 6188 20698 6244 20700
rect 6268 20698 6324 20700
rect 6348 20698 6404 20700
rect 6108 20646 6154 20698
rect 6154 20646 6164 20698
rect 6188 20646 6218 20698
rect 6218 20646 6230 20698
rect 6230 20646 6244 20698
rect 6268 20646 6282 20698
rect 6282 20646 6294 20698
rect 6294 20646 6324 20698
rect 6348 20646 6358 20698
rect 6358 20646 6404 20698
rect 6108 20644 6164 20646
rect 6188 20644 6244 20646
rect 6268 20644 6324 20646
rect 6348 20644 6404 20646
rect 6108 19610 6164 19612
rect 6188 19610 6244 19612
rect 6268 19610 6324 19612
rect 6348 19610 6404 19612
rect 6108 19558 6154 19610
rect 6154 19558 6164 19610
rect 6188 19558 6218 19610
rect 6218 19558 6230 19610
rect 6230 19558 6244 19610
rect 6268 19558 6282 19610
rect 6282 19558 6294 19610
rect 6294 19558 6324 19610
rect 6348 19558 6358 19610
rect 6358 19558 6404 19610
rect 6108 19556 6164 19558
rect 6188 19556 6244 19558
rect 6268 19556 6324 19558
rect 6348 19556 6404 19558
rect 6108 18522 6164 18524
rect 6188 18522 6244 18524
rect 6268 18522 6324 18524
rect 6348 18522 6404 18524
rect 6108 18470 6154 18522
rect 6154 18470 6164 18522
rect 6188 18470 6218 18522
rect 6218 18470 6230 18522
rect 6230 18470 6244 18522
rect 6268 18470 6282 18522
rect 6282 18470 6294 18522
rect 6294 18470 6324 18522
rect 6348 18470 6358 18522
rect 6358 18470 6404 18522
rect 6108 18468 6164 18470
rect 6188 18468 6244 18470
rect 6268 18468 6324 18470
rect 6348 18468 6404 18470
rect 6108 17434 6164 17436
rect 6188 17434 6244 17436
rect 6268 17434 6324 17436
rect 6348 17434 6404 17436
rect 6108 17382 6154 17434
rect 6154 17382 6164 17434
rect 6188 17382 6218 17434
rect 6218 17382 6230 17434
rect 6230 17382 6244 17434
rect 6268 17382 6282 17434
rect 6282 17382 6294 17434
rect 6294 17382 6324 17434
rect 6348 17382 6358 17434
rect 6358 17382 6404 17434
rect 6108 17380 6164 17382
rect 6188 17380 6244 17382
rect 6268 17380 6324 17382
rect 6348 17380 6404 17382
rect 6108 16346 6164 16348
rect 6188 16346 6244 16348
rect 6268 16346 6324 16348
rect 6348 16346 6404 16348
rect 6108 16294 6154 16346
rect 6154 16294 6164 16346
rect 6188 16294 6218 16346
rect 6218 16294 6230 16346
rect 6230 16294 6244 16346
rect 6268 16294 6282 16346
rect 6282 16294 6294 16346
rect 6294 16294 6324 16346
rect 6348 16294 6358 16346
rect 6358 16294 6404 16346
rect 6108 16292 6164 16294
rect 6188 16292 6244 16294
rect 6268 16292 6324 16294
rect 6348 16292 6404 16294
rect 6108 15258 6164 15260
rect 6188 15258 6244 15260
rect 6268 15258 6324 15260
rect 6348 15258 6404 15260
rect 6108 15206 6154 15258
rect 6154 15206 6164 15258
rect 6188 15206 6218 15258
rect 6218 15206 6230 15258
rect 6230 15206 6244 15258
rect 6268 15206 6282 15258
rect 6282 15206 6294 15258
rect 6294 15206 6324 15258
rect 6348 15206 6358 15258
rect 6358 15206 6404 15258
rect 6108 15204 6164 15206
rect 6188 15204 6244 15206
rect 6268 15204 6324 15206
rect 6348 15204 6404 15206
rect 6108 14170 6164 14172
rect 6188 14170 6244 14172
rect 6268 14170 6324 14172
rect 6348 14170 6404 14172
rect 6108 14118 6154 14170
rect 6154 14118 6164 14170
rect 6188 14118 6218 14170
rect 6218 14118 6230 14170
rect 6230 14118 6244 14170
rect 6268 14118 6282 14170
rect 6282 14118 6294 14170
rect 6294 14118 6324 14170
rect 6348 14118 6358 14170
rect 6358 14118 6404 14170
rect 6108 14116 6164 14118
rect 6188 14116 6244 14118
rect 6268 14116 6324 14118
rect 6348 14116 6404 14118
rect 6108 13082 6164 13084
rect 6188 13082 6244 13084
rect 6268 13082 6324 13084
rect 6348 13082 6404 13084
rect 6108 13030 6154 13082
rect 6154 13030 6164 13082
rect 6188 13030 6218 13082
rect 6218 13030 6230 13082
rect 6230 13030 6244 13082
rect 6268 13030 6282 13082
rect 6282 13030 6294 13082
rect 6294 13030 6324 13082
rect 6348 13030 6358 13082
rect 6358 13030 6404 13082
rect 6108 13028 6164 13030
rect 6188 13028 6244 13030
rect 6268 13028 6324 13030
rect 6348 13028 6404 13030
rect 11259 47354 11315 47356
rect 11339 47354 11395 47356
rect 11419 47354 11475 47356
rect 11499 47354 11555 47356
rect 11259 47302 11305 47354
rect 11305 47302 11315 47354
rect 11339 47302 11369 47354
rect 11369 47302 11381 47354
rect 11381 47302 11395 47354
rect 11419 47302 11433 47354
rect 11433 47302 11445 47354
rect 11445 47302 11475 47354
rect 11499 47302 11509 47354
rect 11509 47302 11555 47354
rect 11259 47300 11315 47302
rect 11339 47300 11395 47302
rect 11419 47300 11475 47302
rect 11499 47300 11555 47302
rect 11259 46266 11315 46268
rect 11339 46266 11395 46268
rect 11419 46266 11475 46268
rect 11499 46266 11555 46268
rect 11259 46214 11305 46266
rect 11305 46214 11315 46266
rect 11339 46214 11369 46266
rect 11369 46214 11381 46266
rect 11381 46214 11395 46266
rect 11419 46214 11433 46266
rect 11433 46214 11445 46266
rect 11445 46214 11475 46266
rect 11499 46214 11509 46266
rect 11509 46214 11555 46266
rect 11259 46212 11315 46214
rect 11339 46212 11395 46214
rect 11419 46212 11475 46214
rect 11499 46212 11555 46214
rect 11259 45178 11315 45180
rect 11339 45178 11395 45180
rect 11419 45178 11475 45180
rect 11499 45178 11555 45180
rect 11259 45126 11305 45178
rect 11305 45126 11315 45178
rect 11339 45126 11369 45178
rect 11369 45126 11381 45178
rect 11381 45126 11395 45178
rect 11419 45126 11433 45178
rect 11433 45126 11445 45178
rect 11445 45126 11475 45178
rect 11499 45126 11509 45178
rect 11509 45126 11555 45178
rect 11259 45124 11315 45126
rect 11339 45124 11395 45126
rect 11419 45124 11475 45126
rect 11499 45124 11555 45126
rect 11259 44090 11315 44092
rect 11339 44090 11395 44092
rect 11419 44090 11475 44092
rect 11499 44090 11555 44092
rect 11259 44038 11305 44090
rect 11305 44038 11315 44090
rect 11339 44038 11369 44090
rect 11369 44038 11381 44090
rect 11381 44038 11395 44090
rect 11419 44038 11433 44090
rect 11433 44038 11445 44090
rect 11445 44038 11475 44090
rect 11499 44038 11509 44090
rect 11509 44038 11555 44090
rect 11259 44036 11315 44038
rect 11339 44036 11395 44038
rect 11419 44036 11475 44038
rect 11499 44036 11555 44038
rect 11259 43002 11315 43004
rect 11339 43002 11395 43004
rect 11419 43002 11475 43004
rect 11499 43002 11555 43004
rect 11259 42950 11305 43002
rect 11305 42950 11315 43002
rect 11339 42950 11369 43002
rect 11369 42950 11381 43002
rect 11381 42950 11395 43002
rect 11419 42950 11433 43002
rect 11433 42950 11445 43002
rect 11445 42950 11475 43002
rect 11499 42950 11509 43002
rect 11509 42950 11555 43002
rect 11259 42948 11315 42950
rect 11339 42948 11395 42950
rect 11419 42948 11475 42950
rect 11499 42948 11555 42950
rect 6108 11994 6164 11996
rect 6188 11994 6244 11996
rect 6268 11994 6324 11996
rect 6348 11994 6404 11996
rect 6108 11942 6154 11994
rect 6154 11942 6164 11994
rect 6188 11942 6218 11994
rect 6218 11942 6230 11994
rect 6230 11942 6244 11994
rect 6268 11942 6282 11994
rect 6282 11942 6294 11994
rect 6294 11942 6324 11994
rect 6348 11942 6358 11994
rect 6358 11942 6404 11994
rect 6108 11940 6164 11942
rect 6188 11940 6244 11942
rect 6268 11940 6324 11942
rect 6348 11940 6404 11942
rect 6108 10906 6164 10908
rect 6188 10906 6244 10908
rect 6268 10906 6324 10908
rect 6348 10906 6404 10908
rect 6108 10854 6154 10906
rect 6154 10854 6164 10906
rect 6188 10854 6218 10906
rect 6218 10854 6230 10906
rect 6230 10854 6244 10906
rect 6268 10854 6282 10906
rect 6282 10854 6294 10906
rect 6294 10854 6324 10906
rect 6348 10854 6358 10906
rect 6358 10854 6404 10906
rect 6108 10852 6164 10854
rect 6188 10852 6244 10854
rect 6268 10852 6324 10854
rect 6348 10852 6404 10854
rect 6108 9818 6164 9820
rect 6188 9818 6244 9820
rect 6268 9818 6324 9820
rect 6348 9818 6404 9820
rect 6108 9766 6154 9818
rect 6154 9766 6164 9818
rect 6188 9766 6218 9818
rect 6218 9766 6230 9818
rect 6230 9766 6244 9818
rect 6268 9766 6282 9818
rect 6282 9766 6294 9818
rect 6294 9766 6324 9818
rect 6348 9766 6358 9818
rect 6358 9766 6404 9818
rect 6108 9764 6164 9766
rect 6188 9764 6244 9766
rect 6268 9764 6324 9766
rect 6348 9764 6404 9766
rect 6108 8730 6164 8732
rect 6188 8730 6244 8732
rect 6268 8730 6324 8732
rect 6348 8730 6404 8732
rect 6108 8678 6154 8730
rect 6154 8678 6164 8730
rect 6188 8678 6218 8730
rect 6218 8678 6230 8730
rect 6230 8678 6244 8730
rect 6268 8678 6282 8730
rect 6282 8678 6294 8730
rect 6294 8678 6324 8730
rect 6348 8678 6358 8730
rect 6358 8678 6404 8730
rect 6108 8676 6164 8678
rect 6188 8676 6244 8678
rect 6268 8676 6324 8678
rect 6348 8676 6404 8678
rect 6108 7642 6164 7644
rect 6188 7642 6244 7644
rect 6268 7642 6324 7644
rect 6348 7642 6404 7644
rect 6108 7590 6154 7642
rect 6154 7590 6164 7642
rect 6188 7590 6218 7642
rect 6218 7590 6230 7642
rect 6230 7590 6244 7642
rect 6268 7590 6282 7642
rect 6282 7590 6294 7642
rect 6294 7590 6324 7642
rect 6348 7590 6358 7642
rect 6358 7590 6404 7642
rect 6108 7588 6164 7590
rect 6188 7588 6244 7590
rect 6268 7588 6324 7590
rect 6348 7588 6404 7590
rect 6108 6554 6164 6556
rect 6188 6554 6244 6556
rect 6268 6554 6324 6556
rect 6348 6554 6404 6556
rect 6108 6502 6154 6554
rect 6154 6502 6164 6554
rect 6188 6502 6218 6554
rect 6218 6502 6230 6554
rect 6230 6502 6244 6554
rect 6268 6502 6282 6554
rect 6282 6502 6294 6554
rect 6294 6502 6324 6554
rect 6348 6502 6358 6554
rect 6358 6502 6404 6554
rect 6108 6500 6164 6502
rect 6188 6500 6244 6502
rect 6268 6500 6324 6502
rect 6348 6500 6404 6502
rect 6108 5466 6164 5468
rect 6188 5466 6244 5468
rect 6268 5466 6324 5468
rect 6348 5466 6404 5468
rect 6108 5414 6154 5466
rect 6154 5414 6164 5466
rect 6188 5414 6218 5466
rect 6218 5414 6230 5466
rect 6230 5414 6244 5466
rect 6268 5414 6282 5466
rect 6282 5414 6294 5466
rect 6294 5414 6324 5466
rect 6348 5414 6358 5466
rect 6358 5414 6404 5466
rect 6108 5412 6164 5414
rect 6188 5412 6244 5414
rect 6268 5412 6324 5414
rect 6348 5412 6404 5414
rect 6108 4378 6164 4380
rect 6188 4378 6244 4380
rect 6268 4378 6324 4380
rect 6348 4378 6404 4380
rect 6108 4326 6154 4378
rect 6154 4326 6164 4378
rect 6188 4326 6218 4378
rect 6218 4326 6230 4378
rect 6230 4326 6244 4378
rect 6268 4326 6282 4378
rect 6282 4326 6294 4378
rect 6294 4326 6324 4378
rect 6348 4326 6358 4378
rect 6358 4326 6404 4378
rect 6108 4324 6164 4326
rect 6188 4324 6244 4326
rect 6268 4324 6324 4326
rect 6348 4324 6404 4326
rect 6108 3290 6164 3292
rect 6188 3290 6244 3292
rect 6268 3290 6324 3292
rect 6348 3290 6404 3292
rect 6108 3238 6154 3290
rect 6154 3238 6164 3290
rect 6188 3238 6218 3290
rect 6218 3238 6230 3290
rect 6230 3238 6244 3290
rect 6268 3238 6282 3290
rect 6282 3238 6294 3290
rect 6294 3238 6324 3290
rect 6348 3238 6358 3290
rect 6358 3238 6404 3290
rect 6108 3236 6164 3238
rect 6188 3236 6244 3238
rect 6268 3236 6324 3238
rect 6348 3236 6404 3238
rect 6108 2202 6164 2204
rect 6188 2202 6244 2204
rect 6268 2202 6324 2204
rect 6348 2202 6404 2204
rect 6108 2150 6154 2202
rect 6154 2150 6164 2202
rect 6188 2150 6218 2202
rect 6218 2150 6230 2202
rect 6230 2150 6244 2202
rect 6268 2150 6282 2202
rect 6282 2150 6294 2202
rect 6294 2150 6324 2202
rect 6348 2150 6358 2202
rect 6358 2150 6404 2202
rect 6108 2148 6164 2150
rect 6188 2148 6244 2150
rect 6268 2148 6324 2150
rect 6348 2148 6404 2150
rect 11259 41914 11315 41916
rect 11339 41914 11395 41916
rect 11419 41914 11475 41916
rect 11499 41914 11555 41916
rect 11259 41862 11305 41914
rect 11305 41862 11315 41914
rect 11339 41862 11369 41914
rect 11369 41862 11381 41914
rect 11381 41862 11395 41914
rect 11419 41862 11433 41914
rect 11433 41862 11445 41914
rect 11445 41862 11475 41914
rect 11499 41862 11509 41914
rect 11509 41862 11555 41914
rect 11259 41860 11315 41862
rect 11339 41860 11395 41862
rect 11419 41860 11475 41862
rect 11499 41860 11555 41862
rect 11259 40826 11315 40828
rect 11339 40826 11395 40828
rect 11419 40826 11475 40828
rect 11499 40826 11555 40828
rect 11259 40774 11305 40826
rect 11305 40774 11315 40826
rect 11339 40774 11369 40826
rect 11369 40774 11381 40826
rect 11381 40774 11395 40826
rect 11419 40774 11433 40826
rect 11433 40774 11445 40826
rect 11445 40774 11475 40826
rect 11499 40774 11509 40826
rect 11509 40774 11555 40826
rect 11259 40772 11315 40774
rect 11339 40772 11395 40774
rect 11419 40772 11475 40774
rect 11499 40772 11555 40774
rect 11259 39738 11315 39740
rect 11339 39738 11395 39740
rect 11419 39738 11475 39740
rect 11499 39738 11555 39740
rect 11259 39686 11305 39738
rect 11305 39686 11315 39738
rect 11339 39686 11369 39738
rect 11369 39686 11381 39738
rect 11381 39686 11395 39738
rect 11419 39686 11433 39738
rect 11433 39686 11445 39738
rect 11445 39686 11475 39738
rect 11499 39686 11509 39738
rect 11509 39686 11555 39738
rect 11259 39684 11315 39686
rect 11339 39684 11395 39686
rect 11419 39684 11475 39686
rect 11499 39684 11555 39686
rect 11259 38650 11315 38652
rect 11339 38650 11395 38652
rect 11419 38650 11475 38652
rect 11499 38650 11555 38652
rect 11259 38598 11305 38650
rect 11305 38598 11315 38650
rect 11339 38598 11369 38650
rect 11369 38598 11381 38650
rect 11381 38598 11395 38650
rect 11419 38598 11433 38650
rect 11433 38598 11445 38650
rect 11445 38598 11475 38650
rect 11499 38598 11509 38650
rect 11509 38598 11555 38650
rect 11259 38596 11315 38598
rect 11339 38596 11395 38598
rect 11419 38596 11475 38598
rect 11499 38596 11555 38598
rect 11259 37562 11315 37564
rect 11339 37562 11395 37564
rect 11419 37562 11475 37564
rect 11499 37562 11555 37564
rect 11259 37510 11305 37562
rect 11305 37510 11315 37562
rect 11339 37510 11369 37562
rect 11369 37510 11381 37562
rect 11381 37510 11395 37562
rect 11419 37510 11433 37562
rect 11433 37510 11445 37562
rect 11445 37510 11475 37562
rect 11499 37510 11509 37562
rect 11509 37510 11555 37562
rect 11259 37508 11315 37510
rect 11339 37508 11395 37510
rect 11419 37508 11475 37510
rect 11499 37508 11555 37510
rect 11259 36474 11315 36476
rect 11339 36474 11395 36476
rect 11419 36474 11475 36476
rect 11499 36474 11555 36476
rect 11259 36422 11305 36474
rect 11305 36422 11315 36474
rect 11339 36422 11369 36474
rect 11369 36422 11381 36474
rect 11381 36422 11395 36474
rect 11419 36422 11433 36474
rect 11433 36422 11445 36474
rect 11445 36422 11475 36474
rect 11499 36422 11509 36474
rect 11509 36422 11555 36474
rect 11259 36420 11315 36422
rect 11339 36420 11395 36422
rect 11419 36420 11475 36422
rect 11499 36420 11555 36422
rect 11259 35386 11315 35388
rect 11339 35386 11395 35388
rect 11419 35386 11475 35388
rect 11499 35386 11555 35388
rect 11259 35334 11305 35386
rect 11305 35334 11315 35386
rect 11339 35334 11369 35386
rect 11369 35334 11381 35386
rect 11381 35334 11395 35386
rect 11419 35334 11433 35386
rect 11433 35334 11445 35386
rect 11445 35334 11475 35386
rect 11499 35334 11509 35386
rect 11509 35334 11555 35386
rect 11259 35332 11315 35334
rect 11339 35332 11395 35334
rect 11419 35332 11475 35334
rect 11499 35332 11555 35334
rect 11259 34298 11315 34300
rect 11339 34298 11395 34300
rect 11419 34298 11475 34300
rect 11499 34298 11555 34300
rect 11259 34246 11305 34298
rect 11305 34246 11315 34298
rect 11339 34246 11369 34298
rect 11369 34246 11381 34298
rect 11381 34246 11395 34298
rect 11419 34246 11433 34298
rect 11433 34246 11445 34298
rect 11445 34246 11475 34298
rect 11499 34246 11509 34298
rect 11509 34246 11555 34298
rect 11259 34244 11315 34246
rect 11339 34244 11395 34246
rect 11419 34244 11475 34246
rect 11499 34244 11555 34246
rect 11259 33210 11315 33212
rect 11339 33210 11395 33212
rect 11419 33210 11475 33212
rect 11499 33210 11555 33212
rect 11259 33158 11305 33210
rect 11305 33158 11315 33210
rect 11339 33158 11369 33210
rect 11369 33158 11381 33210
rect 11381 33158 11395 33210
rect 11419 33158 11433 33210
rect 11433 33158 11445 33210
rect 11445 33158 11475 33210
rect 11499 33158 11509 33210
rect 11509 33158 11555 33210
rect 11259 33156 11315 33158
rect 11339 33156 11395 33158
rect 11419 33156 11475 33158
rect 11499 33156 11555 33158
rect 11259 32122 11315 32124
rect 11339 32122 11395 32124
rect 11419 32122 11475 32124
rect 11499 32122 11555 32124
rect 11259 32070 11305 32122
rect 11305 32070 11315 32122
rect 11339 32070 11369 32122
rect 11369 32070 11381 32122
rect 11381 32070 11395 32122
rect 11419 32070 11433 32122
rect 11433 32070 11445 32122
rect 11445 32070 11475 32122
rect 11499 32070 11509 32122
rect 11509 32070 11555 32122
rect 11259 32068 11315 32070
rect 11339 32068 11395 32070
rect 11419 32068 11475 32070
rect 11499 32068 11555 32070
rect 11259 31034 11315 31036
rect 11339 31034 11395 31036
rect 11419 31034 11475 31036
rect 11499 31034 11555 31036
rect 11259 30982 11305 31034
rect 11305 30982 11315 31034
rect 11339 30982 11369 31034
rect 11369 30982 11381 31034
rect 11381 30982 11395 31034
rect 11419 30982 11433 31034
rect 11433 30982 11445 31034
rect 11445 30982 11475 31034
rect 11499 30982 11509 31034
rect 11509 30982 11555 31034
rect 11259 30980 11315 30982
rect 11339 30980 11395 30982
rect 11419 30980 11475 30982
rect 11499 30980 11555 30982
rect 11259 29946 11315 29948
rect 11339 29946 11395 29948
rect 11419 29946 11475 29948
rect 11499 29946 11555 29948
rect 11259 29894 11305 29946
rect 11305 29894 11315 29946
rect 11339 29894 11369 29946
rect 11369 29894 11381 29946
rect 11381 29894 11395 29946
rect 11419 29894 11433 29946
rect 11433 29894 11445 29946
rect 11445 29894 11475 29946
rect 11499 29894 11509 29946
rect 11509 29894 11555 29946
rect 11259 29892 11315 29894
rect 11339 29892 11395 29894
rect 11419 29892 11475 29894
rect 11499 29892 11555 29894
rect 11259 28858 11315 28860
rect 11339 28858 11395 28860
rect 11419 28858 11475 28860
rect 11499 28858 11555 28860
rect 11259 28806 11305 28858
rect 11305 28806 11315 28858
rect 11339 28806 11369 28858
rect 11369 28806 11381 28858
rect 11381 28806 11395 28858
rect 11419 28806 11433 28858
rect 11433 28806 11445 28858
rect 11445 28806 11475 28858
rect 11499 28806 11509 28858
rect 11509 28806 11555 28858
rect 11259 28804 11315 28806
rect 11339 28804 11395 28806
rect 11419 28804 11475 28806
rect 11499 28804 11555 28806
rect 11259 27770 11315 27772
rect 11339 27770 11395 27772
rect 11419 27770 11475 27772
rect 11499 27770 11555 27772
rect 11259 27718 11305 27770
rect 11305 27718 11315 27770
rect 11339 27718 11369 27770
rect 11369 27718 11381 27770
rect 11381 27718 11395 27770
rect 11419 27718 11433 27770
rect 11433 27718 11445 27770
rect 11445 27718 11475 27770
rect 11499 27718 11509 27770
rect 11509 27718 11555 27770
rect 11259 27716 11315 27718
rect 11339 27716 11395 27718
rect 11419 27716 11475 27718
rect 11499 27716 11555 27718
rect 11259 26682 11315 26684
rect 11339 26682 11395 26684
rect 11419 26682 11475 26684
rect 11499 26682 11555 26684
rect 11259 26630 11305 26682
rect 11305 26630 11315 26682
rect 11339 26630 11369 26682
rect 11369 26630 11381 26682
rect 11381 26630 11395 26682
rect 11419 26630 11433 26682
rect 11433 26630 11445 26682
rect 11445 26630 11475 26682
rect 11499 26630 11509 26682
rect 11509 26630 11555 26682
rect 11259 26628 11315 26630
rect 11339 26628 11395 26630
rect 11419 26628 11475 26630
rect 11499 26628 11555 26630
rect 11259 25594 11315 25596
rect 11339 25594 11395 25596
rect 11419 25594 11475 25596
rect 11499 25594 11555 25596
rect 11259 25542 11305 25594
rect 11305 25542 11315 25594
rect 11339 25542 11369 25594
rect 11369 25542 11381 25594
rect 11381 25542 11395 25594
rect 11419 25542 11433 25594
rect 11433 25542 11445 25594
rect 11445 25542 11475 25594
rect 11499 25542 11509 25594
rect 11509 25542 11555 25594
rect 11259 25540 11315 25542
rect 11339 25540 11395 25542
rect 11419 25540 11475 25542
rect 11499 25540 11555 25542
rect 11259 24506 11315 24508
rect 11339 24506 11395 24508
rect 11419 24506 11475 24508
rect 11499 24506 11555 24508
rect 11259 24454 11305 24506
rect 11305 24454 11315 24506
rect 11339 24454 11369 24506
rect 11369 24454 11381 24506
rect 11381 24454 11395 24506
rect 11419 24454 11433 24506
rect 11433 24454 11445 24506
rect 11445 24454 11475 24506
rect 11499 24454 11509 24506
rect 11509 24454 11555 24506
rect 11259 24452 11315 24454
rect 11339 24452 11395 24454
rect 11419 24452 11475 24454
rect 11499 24452 11555 24454
rect 11259 23418 11315 23420
rect 11339 23418 11395 23420
rect 11419 23418 11475 23420
rect 11499 23418 11555 23420
rect 11259 23366 11305 23418
rect 11305 23366 11315 23418
rect 11339 23366 11369 23418
rect 11369 23366 11381 23418
rect 11381 23366 11395 23418
rect 11419 23366 11433 23418
rect 11433 23366 11445 23418
rect 11445 23366 11475 23418
rect 11499 23366 11509 23418
rect 11509 23366 11555 23418
rect 11259 23364 11315 23366
rect 11339 23364 11395 23366
rect 11419 23364 11475 23366
rect 11499 23364 11555 23366
rect 11259 22330 11315 22332
rect 11339 22330 11395 22332
rect 11419 22330 11475 22332
rect 11499 22330 11555 22332
rect 11259 22278 11305 22330
rect 11305 22278 11315 22330
rect 11339 22278 11369 22330
rect 11369 22278 11381 22330
rect 11381 22278 11395 22330
rect 11419 22278 11433 22330
rect 11433 22278 11445 22330
rect 11445 22278 11475 22330
rect 11499 22278 11509 22330
rect 11509 22278 11555 22330
rect 11259 22276 11315 22278
rect 11339 22276 11395 22278
rect 11419 22276 11475 22278
rect 11499 22276 11555 22278
rect 11259 21242 11315 21244
rect 11339 21242 11395 21244
rect 11419 21242 11475 21244
rect 11499 21242 11555 21244
rect 11259 21190 11305 21242
rect 11305 21190 11315 21242
rect 11339 21190 11369 21242
rect 11369 21190 11381 21242
rect 11381 21190 11395 21242
rect 11419 21190 11433 21242
rect 11433 21190 11445 21242
rect 11445 21190 11475 21242
rect 11499 21190 11509 21242
rect 11509 21190 11555 21242
rect 11259 21188 11315 21190
rect 11339 21188 11395 21190
rect 11419 21188 11475 21190
rect 11499 21188 11555 21190
rect 11259 20154 11315 20156
rect 11339 20154 11395 20156
rect 11419 20154 11475 20156
rect 11499 20154 11555 20156
rect 11259 20102 11305 20154
rect 11305 20102 11315 20154
rect 11339 20102 11369 20154
rect 11369 20102 11381 20154
rect 11381 20102 11395 20154
rect 11419 20102 11433 20154
rect 11433 20102 11445 20154
rect 11445 20102 11475 20154
rect 11499 20102 11509 20154
rect 11509 20102 11555 20154
rect 11259 20100 11315 20102
rect 11339 20100 11395 20102
rect 11419 20100 11475 20102
rect 11499 20100 11555 20102
rect 11259 19066 11315 19068
rect 11339 19066 11395 19068
rect 11419 19066 11475 19068
rect 11499 19066 11555 19068
rect 11259 19014 11305 19066
rect 11305 19014 11315 19066
rect 11339 19014 11369 19066
rect 11369 19014 11381 19066
rect 11381 19014 11395 19066
rect 11419 19014 11433 19066
rect 11433 19014 11445 19066
rect 11445 19014 11475 19066
rect 11499 19014 11509 19066
rect 11509 19014 11555 19066
rect 11259 19012 11315 19014
rect 11339 19012 11395 19014
rect 11419 19012 11475 19014
rect 11499 19012 11555 19014
rect 11259 17978 11315 17980
rect 11339 17978 11395 17980
rect 11419 17978 11475 17980
rect 11499 17978 11555 17980
rect 11259 17926 11305 17978
rect 11305 17926 11315 17978
rect 11339 17926 11369 17978
rect 11369 17926 11381 17978
rect 11381 17926 11395 17978
rect 11419 17926 11433 17978
rect 11433 17926 11445 17978
rect 11445 17926 11475 17978
rect 11499 17926 11509 17978
rect 11509 17926 11555 17978
rect 11259 17924 11315 17926
rect 11339 17924 11395 17926
rect 11419 17924 11475 17926
rect 11499 17924 11555 17926
rect 11259 16890 11315 16892
rect 11339 16890 11395 16892
rect 11419 16890 11475 16892
rect 11499 16890 11555 16892
rect 11259 16838 11305 16890
rect 11305 16838 11315 16890
rect 11339 16838 11369 16890
rect 11369 16838 11381 16890
rect 11381 16838 11395 16890
rect 11419 16838 11433 16890
rect 11433 16838 11445 16890
rect 11445 16838 11475 16890
rect 11499 16838 11509 16890
rect 11509 16838 11555 16890
rect 11259 16836 11315 16838
rect 11339 16836 11395 16838
rect 11419 16836 11475 16838
rect 11499 16836 11555 16838
rect 11259 15802 11315 15804
rect 11339 15802 11395 15804
rect 11419 15802 11475 15804
rect 11499 15802 11555 15804
rect 11259 15750 11305 15802
rect 11305 15750 11315 15802
rect 11339 15750 11369 15802
rect 11369 15750 11381 15802
rect 11381 15750 11395 15802
rect 11419 15750 11433 15802
rect 11433 15750 11445 15802
rect 11445 15750 11475 15802
rect 11499 15750 11509 15802
rect 11509 15750 11555 15802
rect 11259 15748 11315 15750
rect 11339 15748 11395 15750
rect 11419 15748 11475 15750
rect 11499 15748 11555 15750
rect 11259 14714 11315 14716
rect 11339 14714 11395 14716
rect 11419 14714 11475 14716
rect 11499 14714 11555 14716
rect 11259 14662 11305 14714
rect 11305 14662 11315 14714
rect 11339 14662 11369 14714
rect 11369 14662 11381 14714
rect 11381 14662 11395 14714
rect 11419 14662 11433 14714
rect 11433 14662 11445 14714
rect 11445 14662 11475 14714
rect 11499 14662 11509 14714
rect 11509 14662 11555 14714
rect 11259 14660 11315 14662
rect 11339 14660 11395 14662
rect 11419 14660 11475 14662
rect 11499 14660 11555 14662
rect 11259 13626 11315 13628
rect 11339 13626 11395 13628
rect 11419 13626 11475 13628
rect 11499 13626 11555 13628
rect 11259 13574 11305 13626
rect 11305 13574 11315 13626
rect 11339 13574 11369 13626
rect 11369 13574 11381 13626
rect 11381 13574 11395 13626
rect 11419 13574 11433 13626
rect 11433 13574 11445 13626
rect 11445 13574 11475 13626
rect 11499 13574 11509 13626
rect 11509 13574 11555 13626
rect 11259 13572 11315 13574
rect 11339 13572 11395 13574
rect 11419 13572 11475 13574
rect 11499 13572 11555 13574
rect 6108 1114 6164 1116
rect 6188 1114 6244 1116
rect 6268 1114 6324 1116
rect 6348 1114 6404 1116
rect 6108 1062 6154 1114
rect 6154 1062 6164 1114
rect 6188 1062 6218 1114
rect 6218 1062 6230 1114
rect 6230 1062 6244 1114
rect 6268 1062 6282 1114
rect 6282 1062 6294 1114
rect 6294 1062 6324 1114
rect 6348 1062 6358 1114
rect 6358 1062 6404 1114
rect 6108 1060 6164 1062
rect 6188 1060 6244 1062
rect 6268 1060 6324 1062
rect 6348 1060 6404 1062
rect 11259 12538 11315 12540
rect 11339 12538 11395 12540
rect 11419 12538 11475 12540
rect 11499 12538 11555 12540
rect 11259 12486 11305 12538
rect 11305 12486 11315 12538
rect 11339 12486 11369 12538
rect 11369 12486 11381 12538
rect 11381 12486 11395 12538
rect 11419 12486 11433 12538
rect 11433 12486 11445 12538
rect 11445 12486 11475 12538
rect 11499 12486 11509 12538
rect 11509 12486 11555 12538
rect 11259 12484 11315 12486
rect 11339 12484 11395 12486
rect 11419 12484 11475 12486
rect 11499 12484 11555 12486
rect 11259 11450 11315 11452
rect 11339 11450 11395 11452
rect 11419 11450 11475 11452
rect 11499 11450 11555 11452
rect 11259 11398 11305 11450
rect 11305 11398 11315 11450
rect 11339 11398 11369 11450
rect 11369 11398 11381 11450
rect 11381 11398 11395 11450
rect 11419 11398 11433 11450
rect 11433 11398 11445 11450
rect 11445 11398 11475 11450
rect 11499 11398 11509 11450
rect 11509 11398 11555 11450
rect 11259 11396 11315 11398
rect 11339 11396 11395 11398
rect 11419 11396 11475 11398
rect 11499 11396 11555 11398
rect 11259 10362 11315 10364
rect 11339 10362 11395 10364
rect 11419 10362 11475 10364
rect 11499 10362 11555 10364
rect 11259 10310 11305 10362
rect 11305 10310 11315 10362
rect 11339 10310 11369 10362
rect 11369 10310 11381 10362
rect 11381 10310 11395 10362
rect 11419 10310 11433 10362
rect 11433 10310 11445 10362
rect 11445 10310 11475 10362
rect 11499 10310 11509 10362
rect 11509 10310 11555 10362
rect 11259 10308 11315 10310
rect 11339 10308 11395 10310
rect 11419 10308 11475 10310
rect 11499 10308 11555 10310
rect 11259 9274 11315 9276
rect 11339 9274 11395 9276
rect 11419 9274 11475 9276
rect 11499 9274 11555 9276
rect 11259 9222 11305 9274
rect 11305 9222 11315 9274
rect 11339 9222 11369 9274
rect 11369 9222 11381 9274
rect 11381 9222 11395 9274
rect 11419 9222 11433 9274
rect 11433 9222 11445 9274
rect 11445 9222 11475 9274
rect 11499 9222 11509 9274
rect 11509 9222 11555 9274
rect 11259 9220 11315 9222
rect 11339 9220 11395 9222
rect 11419 9220 11475 9222
rect 11499 9220 11555 9222
rect 11259 8186 11315 8188
rect 11339 8186 11395 8188
rect 11419 8186 11475 8188
rect 11499 8186 11555 8188
rect 11259 8134 11305 8186
rect 11305 8134 11315 8186
rect 11339 8134 11369 8186
rect 11369 8134 11381 8186
rect 11381 8134 11395 8186
rect 11419 8134 11433 8186
rect 11433 8134 11445 8186
rect 11445 8134 11475 8186
rect 11499 8134 11509 8186
rect 11509 8134 11555 8186
rect 11259 8132 11315 8134
rect 11339 8132 11395 8134
rect 11419 8132 11475 8134
rect 11499 8132 11555 8134
rect 11259 7098 11315 7100
rect 11339 7098 11395 7100
rect 11419 7098 11475 7100
rect 11499 7098 11555 7100
rect 11259 7046 11305 7098
rect 11305 7046 11315 7098
rect 11339 7046 11369 7098
rect 11369 7046 11381 7098
rect 11381 7046 11395 7098
rect 11419 7046 11433 7098
rect 11433 7046 11445 7098
rect 11445 7046 11475 7098
rect 11499 7046 11509 7098
rect 11509 7046 11555 7098
rect 11259 7044 11315 7046
rect 11339 7044 11395 7046
rect 11419 7044 11475 7046
rect 11499 7044 11555 7046
rect 11259 6010 11315 6012
rect 11339 6010 11395 6012
rect 11419 6010 11475 6012
rect 11499 6010 11555 6012
rect 11259 5958 11305 6010
rect 11305 5958 11315 6010
rect 11339 5958 11369 6010
rect 11369 5958 11381 6010
rect 11381 5958 11395 6010
rect 11419 5958 11433 6010
rect 11433 5958 11445 6010
rect 11445 5958 11475 6010
rect 11499 5958 11509 6010
rect 11509 5958 11555 6010
rect 11259 5956 11315 5958
rect 11339 5956 11395 5958
rect 11419 5956 11475 5958
rect 11499 5956 11555 5958
rect 11259 4922 11315 4924
rect 11339 4922 11395 4924
rect 11419 4922 11475 4924
rect 11499 4922 11555 4924
rect 11259 4870 11305 4922
rect 11305 4870 11315 4922
rect 11339 4870 11369 4922
rect 11369 4870 11381 4922
rect 11381 4870 11395 4922
rect 11419 4870 11433 4922
rect 11433 4870 11445 4922
rect 11445 4870 11475 4922
rect 11499 4870 11509 4922
rect 11509 4870 11555 4922
rect 11259 4868 11315 4870
rect 11339 4868 11395 4870
rect 11419 4868 11475 4870
rect 11499 4868 11555 4870
rect 11259 3834 11315 3836
rect 11339 3834 11395 3836
rect 11419 3834 11475 3836
rect 11499 3834 11555 3836
rect 11259 3782 11305 3834
rect 11305 3782 11315 3834
rect 11339 3782 11369 3834
rect 11369 3782 11381 3834
rect 11381 3782 11395 3834
rect 11419 3782 11433 3834
rect 11433 3782 11445 3834
rect 11445 3782 11475 3834
rect 11499 3782 11509 3834
rect 11509 3782 11555 3834
rect 11259 3780 11315 3782
rect 11339 3780 11395 3782
rect 11419 3780 11475 3782
rect 11499 3780 11555 3782
rect 11259 2746 11315 2748
rect 11339 2746 11395 2748
rect 11419 2746 11475 2748
rect 11499 2746 11555 2748
rect 11259 2694 11305 2746
rect 11305 2694 11315 2746
rect 11339 2694 11369 2746
rect 11369 2694 11381 2746
rect 11381 2694 11395 2746
rect 11419 2694 11433 2746
rect 11433 2694 11445 2746
rect 11445 2694 11475 2746
rect 11499 2694 11509 2746
rect 11509 2694 11555 2746
rect 11259 2692 11315 2694
rect 11339 2692 11395 2694
rect 11419 2692 11475 2694
rect 11499 2692 11555 2694
rect 11259 1658 11315 1660
rect 11339 1658 11395 1660
rect 11419 1658 11475 1660
rect 11499 1658 11555 1660
rect 11259 1606 11305 1658
rect 11305 1606 11315 1658
rect 11339 1606 11369 1658
rect 11369 1606 11381 1658
rect 11381 1606 11395 1658
rect 11419 1606 11433 1658
rect 11433 1606 11445 1658
rect 11445 1606 11475 1658
rect 11499 1606 11509 1658
rect 11509 1606 11555 1658
rect 11259 1604 11315 1606
rect 11339 1604 11395 1606
rect 11419 1604 11475 1606
rect 11499 1604 11555 1606
rect 16411 47898 16467 47900
rect 16491 47898 16547 47900
rect 16571 47898 16627 47900
rect 16651 47898 16707 47900
rect 16411 47846 16457 47898
rect 16457 47846 16467 47898
rect 16491 47846 16521 47898
rect 16521 47846 16533 47898
rect 16533 47846 16547 47898
rect 16571 47846 16585 47898
rect 16585 47846 16597 47898
rect 16597 47846 16627 47898
rect 16651 47846 16661 47898
rect 16661 47846 16707 47898
rect 16411 47844 16467 47846
rect 16491 47844 16547 47846
rect 16571 47844 16627 47846
rect 16651 47844 16707 47846
rect 16411 46810 16467 46812
rect 16491 46810 16547 46812
rect 16571 46810 16627 46812
rect 16651 46810 16707 46812
rect 16411 46758 16457 46810
rect 16457 46758 16467 46810
rect 16491 46758 16521 46810
rect 16521 46758 16533 46810
rect 16533 46758 16547 46810
rect 16571 46758 16585 46810
rect 16585 46758 16597 46810
rect 16597 46758 16627 46810
rect 16651 46758 16661 46810
rect 16661 46758 16707 46810
rect 16411 46756 16467 46758
rect 16491 46756 16547 46758
rect 16571 46756 16627 46758
rect 16651 46756 16707 46758
rect 16411 45722 16467 45724
rect 16491 45722 16547 45724
rect 16571 45722 16627 45724
rect 16651 45722 16707 45724
rect 16411 45670 16457 45722
rect 16457 45670 16467 45722
rect 16491 45670 16521 45722
rect 16521 45670 16533 45722
rect 16533 45670 16547 45722
rect 16571 45670 16585 45722
rect 16585 45670 16597 45722
rect 16597 45670 16627 45722
rect 16651 45670 16661 45722
rect 16661 45670 16707 45722
rect 16411 45668 16467 45670
rect 16491 45668 16547 45670
rect 16571 45668 16627 45670
rect 16651 45668 16707 45670
rect 16411 44634 16467 44636
rect 16491 44634 16547 44636
rect 16571 44634 16627 44636
rect 16651 44634 16707 44636
rect 16411 44582 16457 44634
rect 16457 44582 16467 44634
rect 16491 44582 16521 44634
rect 16521 44582 16533 44634
rect 16533 44582 16547 44634
rect 16571 44582 16585 44634
rect 16585 44582 16597 44634
rect 16597 44582 16627 44634
rect 16651 44582 16661 44634
rect 16661 44582 16707 44634
rect 16411 44580 16467 44582
rect 16491 44580 16547 44582
rect 16571 44580 16627 44582
rect 16651 44580 16707 44582
rect 16411 43546 16467 43548
rect 16491 43546 16547 43548
rect 16571 43546 16627 43548
rect 16651 43546 16707 43548
rect 16411 43494 16457 43546
rect 16457 43494 16467 43546
rect 16491 43494 16521 43546
rect 16521 43494 16533 43546
rect 16533 43494 16547 43546
rect 16571 43494 16585 43546
rect 16585 43494 16597 43546
rect 16597 43494 16627 43546
rect 16651 43494 16661 43546
rect 16661 43494 16707 43546
rect 16411 43492 16467 43494
rect 16491 43492 16547 43494
rect 16571 43492 16627 43494
rect 16651 43492 16707 43494
rect 16411 42458 16467 42460
rect 16491 42458 16547 42460
rect 16571 42458 16627 42460
rect 16651 42458 16707 42460
rect 16411 42406 16457 42458
rect 16457 42406 16467 42458
rect 16491 42406 16521 42458
rect 16521 42406 16533 42458
rect 16533 42406 16547 42458
rect 16571 42406 16585 42458
rect 16585 42406 16597 42458
rect 16597 42406 16627 42458
rect 16651 42406 16661 42458
rect 16661 42406 16707 42458
rect 16411 42404 16467 42406
rect 16491 42404 16547 42406
rect 16571 42404 16627 42406
rect 16651 42404 16707 42406
rect 16411 41370 16467 41372
rect 16491 41370 16547 41372
rect 16571 41370 16627 41372
rect 16651 41370 16707 41372
rect 16411 41318 16457 41370
rect 16457 41318 16467 41370
rect 16491 41318 16521 41370
rect 16521 41318 16533 41370
rect 16533 41318 16547 41370
rect 16571 41318 16585 41370
rect 16585 41318 16597 41370
rect 16597 41318 16627 41370
rect 16651 41318 16661 41370
rect 16661 41318 16707 41370
rect 16411 41316 16467 41318
rect 16491 41316 16547 41318
rect 16571 41316 16627 41318
rect 16651 41316 16707 41318
rect 16411 40282 16467 40284
rect 16491 40282 16547 40284
rect 16571 40282 16627 40284
rect 16651 40282 16707 40284
rect 16411 40230 16457 40282
rect 16457 40230 16467 40282
rect 16491 40230 16521 40282
rect 16521 40230 16533 40282
rect 16533 40230 16547 40282
rect 16571 40230 16585 40282
rect 16585 40230 16597 40282
rect 16597 40230 16627 40282
rect 16651 40230 16661 40282
rect 16661 40230 16707 40282
rect 16411 40228 16467 40230
rect 16491 40228 16547 40230
rect 16571 40228 16627 40230
rect 16651 40228 16707 40230
rect 16411 39194 16467 39196
rect 16491 39194 16547 39196
rect 16571 39194 16627 39196
rect 16651 39194 16707 39196
rect 16411 39142 16457 39194
rect 16457 39142 16467 39194
rect 16491 39142 16521 39194
rect 16521 39142 16533 39194
rect 16533 39142 16547 39194
rect 16571 39142 16585 39194
rect 16585 39142 16597 39194
rect 16597 39142 16627 39194
rect 16651 39142 16661 39194
rect 16661 39142 16707 39194
rect 16411 39140 16467 39142
rect 16491 39140 16547 39142
rect 16571 39140 16627 39142
rect 16651 39140 16707 39142
rect 16411 38106 16467 38108
rect 16491 38106 16547 38108
rect 16571 38106 16627 38108
rect 16651 38106 16707 38108
rect 16411 38054 16457 38106
rect 16457 38054 16467 38106
rect 16491 38054 16521 38106
rect 16521 38054 16533 38106
rect 16533 38054 16547 38106
rect 16571 38054 16585 38106
rect 16585 38054 16597 38106
rect 16597 38054 16627 38106
rect 16651 38054 16661 38106
rect 16661 38054 16707 38106
rect 16411 38052 16467 38054
rect 16491 38052 16547 38054
rect 16571 38052 16627 38054
rect 16651 38052 16707 38054
rect 16411 37018 16467 37020
rect 16491 37018 16547 37020
rect 16571 37018 16627 37020
rect 16651 37018 16707 37020
rect 16411 36966 16457 37018
rect 16457 36966 16467 37018
rect 16491 36966 16521 37018
rect 16521 36966 16533 37018
rect 16533 36966 16547 37018
rect 16571 36966 16585 37018
rect 16585 36966 16597 37018
rect 16597 36966 16627 37018
rect 16651 36966 16661 37018
rect 16661 36966 16707 37018
rect 16411 36964 16467 36966
rect 16491 36964 16547 36966
rect 16571 36964 16627 36966
rect 16651 36964 16707 36966
rect 16411 35930 16467 35932
rect 16491 35930 16547 35932
rect 16571 35930 16627 35932
rect 16651 35930 16707 35932
rect 16411 35878 16457 35930
rect 16457 35878 16467 35930
rect 16491 35878 16521 35930
rect 16521 35878 16533 35930
rect 16533 35878 16547 35930
rect 16571 35878 16585 35930
rect 16585 35878 16597 35930
rect 16597 35878 16627 35930
rect 16651 35878 16661 35930
rect 16661 35878 16707 35930
rect 16411 35876 16467 35878
rect 16491 35876 16547 35878
rect 16571 35876 16627 35878
rect 16651 35876 16707 35878
rect 16411 34842 16467 34844
rect 16491 34842 16547 34844
rect 16571 34842 16627 34844
rect 16651 34842 16707 34844
rect 16411 34790 16457 34842
rect 16457 34790 16467 34842
rect 16491 34790 16521 34842
rect 16521 34790 16533 34842
rect 16533 34790 16547 34842
rect 16571 34790 16585 34842
rect 16585 34790 16597 34842
rect 16597 34790 16627 34842
rect 16651 34790 16661 34842
rect 16661 34790 16707 34842
rect 16411 34788 16467 34790
rect 16491 34788 16547 34790
rect 16571 34788 16627 34790
rect 16651 34788 16707 34790
rect 16411 33754 16467 33756
rect 16491 33754 16547 33756
rect 16571 33754 16627 33756
rect 16651 33754 16707 33756
rect 16411 33702 16457 33754
rect 16457 33702 16467 33754
rect 16491 33702 16521 33754
rect 16521 33702 16533 33754
rect 16533 33702 16547 33754
rect 16571 33702 16585 33754
rect 16585 33702 16597 33754
rect 16597 33702 16627 33754
rect 16651 33702 16661 33754
rect 16661 33702 16707 33754
rect 16411 33700 16467 33702
rect 16491 33700 16547 33702
rect 16571 33700 16627 33702
rect 16651 33700 16707 33702
rect 16411 32666 16467 32668
rect 16491 32666 16547 32668
rect 16571 32666 16627 32668
rect 16651 32666 16707 32668
rect 16411 32614 16457 32666
rect 16457 32614 16467 32666
rect 16491 32614 16521 32666
rect 16521 32614 16533 32666
rect 16533 32614 16547 32666
rect 16571 32614 16585 32666
rect 16585 32614 16597 32666
rect 16597 32614 16627 32666
rect 16651 32614 16661 32666
rect 16661 32614 16707 32666
rect 16411 32612 16467 32614
rect 16491 32612 16547 32614
rect 16571 32612 16627 32614
rect 16651 32612 16707 32614
rect 16411 31578 16467 31580
rect 16491 31578 16547 31580
rect 16571 31578 16627 31580
rect 16651 31578 16707 31580
rect 16411 31526 16457 31578
rect 16457 31526 16467 31578
rect 16491 31526 16521 31578
rect 16521 31526 16533 31578
rect 16533 31526 16547 31578
rect 16571 31526 16585 31578
rect 16585 31526 16597 31578
rect 16597 31526 16627 31578
rect 16651 31526 16661 31578
rect 16661 31526 16707 31578
rect 16411 31524 16467 31526
rect 16491 31524 16547 31526
rect 16571 31524 16627 31526
rect 16651 31524 16707 31526
rect 16411 30490 16467 30492
rect 16491 30490 16547 30492
rect 16571 30490 16627 30492
rect 16651 30490 16707 30492
rect 16411 30438 16457 30490
rect 16457 30438 16467 30490
rect 16491 30438 16521 30490
rect 16521 30438 16533 30490
rect 16533 30438 16547 30490
rect 16571 30438 16585 30490
rect 16585 30438 16597 30490
rect 16597 30438 16627 30490
rect 16651 30438 16661 30490
rect 16661 30438 16707 30490
rect 16411 30436 16467 30438
rect 16491 30436 16547 30438
rect 16571 30436 16627 30438
rect 16651 30436 16707 30438
rect 16411 29402 16467 29404
rect 16491 29402 16547 29404
rect 16571 29402 16627 29404
rect 16651 29402 16707 29404
rect 16411 29350 16457 29402
rect 16457 29350 16467 29402
rect 16491 29350 16521 29402
rect 16521 29350 16533 29402
rect 16533 29350 16547 29402
rect 16571 29350 16585 29402
rect 16585 29350 16597 29402
rect 16597 29350 16627 29402
rect 16651 29350 16661 29402
rect 16661 29350 16707 29402
rect 16411 29348 16467 29350
rect 16491 29348 16547 29350
rect 16571 29348 16627 29350
rect 16651 29348 16707 29350
rect 16411 28314 16467 28316
rect 16491 28314 16547 28316
rect 16571 28314 16627 28316
rect 16651 28314 16707 28316
rect 16411 28262 16457 28314
rect 16457 28262 16467 28314
rect 16491 28262 16521 28314
rect 16521 28262 16533 28314
rect 16533 28262 16547 28314
rect 16571 28262 16585 28314
rect 16585 28262 16597 28314
rect 16597 28262 16627 28314
rect 16651 28262 16661 28314
rect 16661 28262 16707 28314
rect 16411 28260 16467 28262
rect 16491 28260 16547 28262
rect 16571 28260 16627 28262
rect 16651 28260 16707 28262
rect 16411 27226 16467 27228
rect 16491 27226 16547 27228
rect 16571 27226 16627 27228
rect 16651 27226 16707 27228
rect 16411 27174 16457 27226
rect 16457 27174 16467 27226
rect 16491 27174 16521 27226
rect 16521 27174 16533 27226
rect 16533 27174 16547 27226
rect 16571 27174 16585 27226
rect 16585 27174 16597 27226
rect 16597 27174 16627 27226
rect 16651 27174 16661 27226
rect 16661 27174 16707 27226
rect 16411 27172 16467 27174
rect 16491 27172 16547 27174
rect 16571 27172 16627 27174
rect 16651 27172 16707 27174
rect 16411 26138 16467 26140
rect 16491 26138 16547 26140
rect 16571 26138 16627 26140
rect 16651 26138 16707 26140
rect 16411 26086 16457 26138
rect 16457 26086 16467 26138
rect 16491 26086 16521 26138
rect 16521 26086 16533 26138
rect 16533 26086 16547 26138
rect 16571 26086 16585 26138
rect 16585 26086 16597 26138
rect 16597 26086 16627 26138
rect 16651 26086 16661 26138
rect 16661 26086 16707 26138
rect 16411 26084 16467 26086
rect 16491 26084 16547 26086
rect 16571 26084 16627 26086
rect 16651 26084 16707 26086
rect 16411 25050 16467 25052
rect 16491 25050 16547 25052
rect 16571 25050 16627 25052
rect 16651 25050 16707 25052
rect 16411 24998 16457 25050
rect 16457 24998 16467 25050
rect 16491 24998 16521 25050
rect 16521 24998 16533 25050
rect 16533 24998 16547 25050
rect 16571 24998 16585 25050
rect 16585 24998 16597 25050
rect 16597 24998 16627 25050
rect 16651 24998 16661 25050
rect 16661 24998 16707 25050
rect 16411 24996 16467 24998
rect 16491 24996 16547 24998
rect 16571 24996 16627 24998
rect 16651 24996 16707 24998
rect 11259 570 11315 572
rect 11339 570 11395 572
rect 11419 570 11475 572
rect 11499 570 11555 572
rect 11259 518 11305 570
rect 11305 518 11315 570
rect 11339 518 11369 570
rect 11369 518 11381 570
rect 11381 518 11395 570
rect 11419 518 11433 570
rect 11433 518 11445 570
rect 11445 518 11475 570
rect 11499 518 11509 570
rect 11509 518 11555 570
rect 11259 516 11315 518
rect 11339 516 11395 518
rect 11419 516 11475 518
rect 11499 516 11555 518
rect 16411 23962 16467 23964
rect 16491 23962 16547 23964
rect 16571 23962 16627 23964
rect 16651 23962 16707 23964
rect 16411 23910 16457 23962
rect 16457 23910 16467 23962
rect 16491 23910 16521 23962
rect 16521 23910 16533 23962
rect 16533 23910 16547 23962
rect 16571 23910 16585 23962
rect 16585 23910 16597 23962
rect 16597 23910 16627 23962
rect 16651 23910 16661 23962
rect 16661 23910 16707 23962
rect 16411 23908 16467 23910
rect 16491 23908 16547 23910
rect 16571 23908 16627 23910
rect 16651 23908 16707 23910
rect 16411 22874 16467 22876
rect 16491 22874 16547 22876
rect 16571 22874 16627 22876
rect 16651 22874 16707 22876
rect 16411 22822 16457 22874
rect 16457 22822 16467 22874
rect 16491 22822 16521 22874
rect 16521 22822 16533 22874
rect 16533 22822 16547 22874
rect 16571 22822 16585 22874
rect 16585 22822 16597 22874
rect 16597 22822 16627 22874
rect 16651 22822 16661 22874
rect 16661 22822 16707 22874
rect 16411 22820 16467 22822
rect 16491 22820 16547 22822
rect 16571 22820 16627 22822
rect 16651 22820 16707 22822
rect 16411 21786 16467 21788
rect 16491 21786 16547 21788
rect 16571 21786 16627 21788
rect 16651 21786 16707 21788
rect 16411 21734 16457 21786
rect 16457 21734 16467 21786
rect 16491 21734 16521 21786
rect 16521 21734 16533 21786
rect 16533 21734 16547 21786
rect 16571 21734 16585 21786
rect 16585 21734 16597 21786
rect 16597 21734 16627 21786
rect 16651 21734 16661 21786
rect 16661 21734 16707 21786
rect 16411 21732 16467 21734
rect 16491 21732 16547 21734
rect 16571 21732 16627 21734
rect 16651 21732 16707 21734
rect 16411 20698 16467 20700
rect 16491 20698 16547 20700
rect 16571 20698 16627 20700
rect 16651 20698 16707 20700
rect 16411 20646 16457 20698
rect 16457 20646 16467 20698
rect 16491 20646 16521 20698
rect 16521 20646 16533 20698
rect 16533 20646 16547 20698
rect 16571 20646 16585 20698
rect 16585 20646 16597 20698
rect 16597 20646 16627 20698
rect 16651 20646 16661 20698
rect 16661 20646 16707 20698
rect 16411 20644 16467 20646
rect 16491 20644 16547 20646
rect 16571 20644 16627 20646
rect 16651 20644 16707 20646
rect 16411 19610 16467 19612
rect 16491 19610 16547 19612
rect 16571 19610 16627 19612
rect 16651 19610 16707 19612
rect 16411 19558 16457 19610
rect 16457 19558 16467 19610
rect 16491 19558 16521 19610
rect 16521 19558 16533 19610
rect 16533 19558 16547 19610
rect 16571 19558 16585 19610
rect 16585 19558 16597 19610
rect 16597 19558 16627 19610
rect 16651 19558 16661 19610
rect 16661 19558 16707 19610
rect 16411 19556 16467 19558
rect 16491 19556 16547 19558
rect 16571 19556 16627 19558
rect 16651 19556 16707 19558
rect 16411 18522 16467 18524
rect 16491 18522 16547 18524
rect 16571 18522 16627 18524
rect 16651 18522 16707 18524
rect 16411 18470 16457 18522
rect 16457 18470 16467 18522
rect 16491 18470 16521 18522
rect 16521 18470 16533 18522
rect 16533 18470 16547 18522
rect 16571 18470 16585 18522
rect 16585 18470 16597 18522
rect 16597 18470 16627 18522
rect 16651 18470 16661 18522
rect 16661 18470 16707 18522
rect 16411 18468 16467 18470
rect 16491 18468 16547 18470
rect 16571 18468 16627 18470
rect 16651 18468 16707 18470
rect 16411 17434 16467 17436
rect 16491 17434 16547 17436
rect 16571 17434 16627 17436
rect 16651 17434 16707 17436
rect 16411 17382 16457 17434
rect 16457 17382 16467 17434
rect 16491 17382 16521 17434
rect 16521 17382 16533 17434
rect 16533 17382 16547 17434
rect 16571 17382 16585 17434
rect 16585 17382 16597 17434
rect 16597 17382 16627 17434
rect 16651 17382 16661 17434
rect 16661 17382 16707 17434
rect 16411 17380 16467 17382
rect 16491 17380 16547 17382
rect 16571 17380 16627 17382
rect 16651 17380 16707 17382
rect 16411 16346 16467 16348
rect 16491 16346 16547 16348
rect 16571 16346 16627 16348
rect 16651 16346 16707 16348
rect 16411 16294 16457 16346
rect 16457 16294 16467 16346
rect 16491 16294 16521 16346
rect 16521 16294 16533 16346
rect 16533 16294 16547 16346
rect 16571 16294 16585 16346
rect 16585 16294 16597 16346
rect 16597 16294 16627 16346
rect 16651 16294 16661 16346
rect 16661 16294 16707 16346
rect 16411 16292 16467 16294
rect 16491 16292 16547 16294
rect 16571 16292 16627 16294
rect 16651 16292 16707 16294
rect 16411 15258 16467 15260
rect 16491 15258 16547 15260
rect 16571 15258 16627 15260
rect 16651 15258 16707 15260
rect 16411 15206 16457 15258
rect 16457 15206 16467 15258
rect 16491 15206 16521 15258
rect 16521 15206 16533 15258
rect 16533 15206 16547 15258
rect 16571 15206 16585 15258
rect 16585 15206 16597 15258
rect 16597 15206 16627 15258
rect 16651 15206 16661 15258
rect 16661 15206 16707 15258
rect 16411 15204 16467 15206
rect 16491 15204 16547 15206
rect 16571 15204 16627 15206
rect 16651 15204 16707 15206
rect 16411 14170 16467 14172
rect 16491 14170 16547 14172
rect 16571 14170 16627 14172
rect 16651 14170 16707 14172
rect 16411 14118 16457 14170
rect 16457 14118 16467 14170
rect 16491 14118 16521 14170
rect 16521 14118 16533 14170
rect 16533 14118 16547 14170
rect 16571 14118 16585 14170
rect 16585 14118 16597 14170
rect 16597 14118 16627 14170
rect 16651 14118 16661 14170
rect 16661 14118 16707 14170
rect 16411 14116 16467 14118
rect 16491 14116 16547 14118
rect 16571 14116 16627 14118
rect 16651 14116 16707 14118
rect 16411 13082 16467 13084
rect 16491 13082 16547 13084
rect 16571 13082 16627 13084
rect 16651 13082 16707 13084
rect 16411 13030 16457 13082
rect 16457 13030 16467 13082
rect 16491 13030 16521 13082
rect 16521 13030 16533 13082
rect 16533 13030 16547 13082
rect 16571 13030 16585 13082
rect 16585 13030 16597 13082
rect 16597 13030 16627 13082
rect 16651 13030 16661 13082
rect 16661 13030 16707 13082
rect 16411 13028 16467 13030
rect 16491 13028 16547 13030
rect 16571 13028 16627 13030
rect 16651 13028 16707 13030
rect 16411 11994 16467 11996
rect 16491 11994 16547 11996
rect 16571 11994 16627 11996
rect 16651 11994 16707 11996
rect 16411 11942 16457 11994
rect 16457 11942 16467 11994
rect 16491 11942 16521 11994
rect 16521 11942 16533 11994
rect 16533 11942 16547 11994
rect 16571 11942 16585 11994
rect 16585 11942 16597 11994
rect 16597 11942 16627 11994
rect 16651 11942 16661 11994
rect 16661 11942 16707 11994
rect 16411 11940 16467 11942
rect 16491 11940 16547 11942
rect 16571 11940 16627 11942
rect 16651 11940 16707 11942
rect 16411 10906 16467 10908
rect 16491 10906 16547 10908
rect 16571 10906 16627 10908
rect 16651 10906 16707 10908
rect 16411 10854 16457 10906
rect 16457 10854 16467 10906
rect 16491 10854 16521 10906
rect 16521 10854 16533 10906
rect 16533 10854 16547 10906
rect 16571 10854 16585 10906
rect 16585 10854 16597 10906
rect 16597 10854 16627 10906
rect 16651 10854 16661 10906
rect 16661 10854 16707 10906
rect 16411 10852 16467 10854
rect 16491 10852 16547 10854
rect 16571 10852 16627 10854
rect 16651 10852 16707 10854
rect 16411 9818 16467 9820
rect 16491 9818 16547 9820
rect 16571 9818 16627 9820
rect 16651 9818 16707 9820
rect 16411 9766 16457 9818
rect 16457 9766 16467 9818
rect 16491 9766 16521 9818
rect 16521 9766 16533 9818
rect 16533 9766 16547 9818
rect 16571 9766 16585 9818
rect 16585 9766 16597 9818
rect 16597 9766 16627 9818
rect 16651 9766 16661 9818
rect 16661 9766 16707 9818
rect 16411 9764 16467 9766
rect 16491 9764 16547 9766
rect 16571 9764 16627 9766
rect 16651 9764 16707 9766
rect 16411 8730 16467 8732
rect 16491 8730 16547 8732
rect 16571 8730 16627 8732
rect 16651 8730 16707 8732
rect 16411 8678 16457 8730
rect 16457 8678 16467 8730
rect 16491 8678 16521 8730
rect 16521 8678 16533 8730
rect 16533 8678 16547 8730
rect 16571 8678 16585 8730
rect 16585 8678 16597 8730
rect 16597 8678 16627 8730
rect 16651 8678 16661 8730
rect 16661 8678 16707 8730
rect 16411 8676 16467 8678
rect 16491 8676 16547 8678
rect 16571 8676 16627 8678
rect 16651 8676 16707 8678
rect 16411 7642 16467 7644
rect 16491 7642 16547 7644
rect 16571 7642 16627 7644
rect 16651 7642 16707 7644
rect 16411 7590 16457 7642
rect 16457 7590 16467 7642
rect 16491 7590 16521 7642
rect 16521 7590 16533 7642
rect 16533 7590 16547 7642
rect 16571 7590 16585 7642
rect 16585 7590 16597 7642
rect 16597 7590 16627 7642
rect 16651 7590 16661 7642
rect 16661 7590 16707 7642
rect 16411 7588 16467 7590
rect 16491 7588 16547 7590
rect 16571 7588 16627 7590
rect 16651 7588 16707 7590
rect 16411 6554 16467 6556
rect 16491 6554 16547 6556
rect 16571 6554 16627 6556
rect 16651 6554 16707 6556
rect 16411 6502 16457 6554
rect 16457 6502 16467 6554
rect 16491 6502 16521 6554
rect 16521 6502 16533 6554
rect 16533 6502 16547 6554
rect 16571 6502 16585 6554
rect 16585 6502 16597 6554
rect 16597 6502 16627 6554
rect 16651 6502 16661 6554
rect 16661 6502 16707 6554
rect 16411 6500 16467 6502
rect 16491 6500 16547 6502
rect 16571 6500 16627 6502
rect 16651 6500 16707 6502
rect 16411 5466 16467 5468
rect 16491 5466 16547 5468
rect 16571 5466 16627 5468
rect 16651 5466 16707 5468
rect 16411 5414 16457 5466
rect 16457 5414 16467 5466
rect 16491 5414 16521 5466
rect 16521 5414 16533 5466
rect 16533 5414 16547 5466
rect 16571 5414 16585 5466
rect 16585 5414 16597 5466
rect 16597 5414 16627 5466
rect 16651 5414 16661 5466
rect 16661 5414 16707 5466
rect 16411 5412 16467 5414
rect 16491 5412 16547 5414
rect 16571 5412 16627 5414
rect 16651 5412 16707 5414
rect 16411 4378 16467 4380
rect 16491 4378 16547 4380
rect 16571 4378 16627 4380
rect 16651 4378 16707 4380
rect 16411 4326 16457 4378
rect 16457 4326 16467 4378
rect 16491 4326 16521 4378
rect 16521 4326 16533 4378
rect 16533 4326 16547 4378
rect 16571 4326 16585 4378
rect 16585 4326 16597 4378
rect 16597 4326 16627 4378
rect 16651 4326 16661 4378
rect 16661 4326 16707 4378
rect 16411 4324 16467 4326
rect 16491 4324 16547 4326
rect 16571 4324 16627 4326
rect 16651 4324 16707 4326
rect 16411 3290 16467 3292
rect 16491 3290 16547 3292
rect 16571 3290 16627 3292
rect 16651 3290 16707 3292
rect 16411 3238 16457 3290
rect 16457 3238 16467 3290
rect 16491 3238 16521 3290
rect 16521 3238 16533 3290
rect 16533 3238 16547 3290
rect 16571 3238 16585 3290
rect 16585 3238 16597 3290
rect 16597 3238 16627 3290
rect 16651 3238 16661 3290
rect 16661 3238 16707 3290
rect 16411 3236 16467 3238
rect 16491 3236 16547 3238
rect 16571 3236 16627 3238
rect 16651 3236 16707 3238
rect 16411 2202 16467 2204
rect 16491 2202 16547 2204
rect 16571 2202 16627 2204
rect 16651 2202 16707 2204
rect 16411 2150 16457 2202
rect 16457 2150 16467 2202
rect 16491 2150 16521 2202
rect 16521 2150 16533 2202
rect 16533 2150 16547 2202
rect 16571 2150 16585 2202
rect 16585 2150 16597 2202
rect 16597 2150 16627 2202
rect 16651 2150 16661 2202
rect 16661 2150 16707 2202
rect 16411 2148 16467 2150
rect 16491 2148 16547 2150
rect 16571 2148 16627 2150
rect 16651 2148 16707 2150
rect 21563 47354 21619 47356
rect 21643 47354 21699 47356
rect 21723 47354 21779 47356
rect 21803 47354 21859 47356
rect 21563 47302 21609 47354
rect 21609 47302 21619 47354
rect 21643 47302 21673 47354
rect 21673 47302 21685 47354
rect 21685 47302 21699 47354
rect 21723 47302 21737 47354
rect 21737 47302 21749 47354
rect 21749 47302 21779 47354
rect 21803 47302 21813 47354
rect 21813 47302 21859 47354
rect 21563 47300 21619 47302
rect 21643 47300 21699 47302
rect 21723 47300 21779 47302
rect 21803 47300 21859 47302
rect 16411 1114 16467 1116
rect 16491 1114 16547 1116
rect 16571 1114 16627 1116
rect 16651 1114 16707 1116
rect 16411 1062 16457 1114
rect 16457 1062 16467 1114
rect 16491 1062 16521 1114
rect 16521 1062 16533 1114
rect 16533 1062 16547 1114
rect 16571 1062 16585 1114
rect 16585 1062 16597 1114
rect 16597 1062 16627 1114
rect 16651 1062 16661 1114
rect 16661 1062 16707 1114
rect 16411 1060 16467 1062
rect 16491 1060 16547 1062
rect 16571 1060 16627 1062
rect 16651 1060 16707 1062
rect 21563 46266 21619 46268
rect 21643 46266 21699 46268
rect 21723 46266 21779 46268
rect 21803 46266 21859 46268
rect 21563 46214 21609 46266
rect 21609 46214 21619 46266
rect 21643 46214 21673 46266
rect 21673 46214 21685 46266
rect 21685 46214 21699 46266
rect 21723 46214 21737 46266
rect 21737 46214 21749 46266
rect 21749 46214 21779 46266
rect 21803 46214 21813 46266
rect 21813 46214 21859 46266
rect 21563 46212 21619 46214
rect 21643 46212 21699 46214
rect 21723 46212 21779 46214
rect 21803 46212 21859 46214
rect 21563 45178 21619 45180
rect 21643 45178 21699 45180
rect 21723 45178 21779 45180
rect 21803 45178 21859 45180
rect 21563 45126 21609 45178
rect 21609 45126 21619 45178
rect 21643 45126 21673 45178
rect 21673 45126 21685 45178
rect 21685 45126 21699 45178
rect 21723 45126 21737 45178
rect 21737 45126 21749 45178
rect 21749 45126 21779 45178
rect 21803 45126 21813 45178
rect 21813 45126 21859 45178
rect 21563 45124 21619 45126
rect 21643 45124 21699 45126
rect 21723 45124 21779 45126
rect 21803 45124 21859 45126
rect 21563 44090 21619 44092
rect 21643 44090 21699 44092
rect 21723 44090 21779 44092
rect 21803 44090 21859 44092
rect 21563 44038 21609 44090
rect 21609 44038 21619 44090
rect 21643 44038 21673 44090
rect 21673 44038 21685 44090
rect 21685 44038 21699 44090
rect 21723 44038 21737 44090
rect 21737 44038 21749 44090
rect 21749 44038 21779 44090
rect 21803 44038 21813 44090
rect 21813 44038 21859 44090
rect 21563 44036 21619 44038
rect 21643 44036 21699 44038
rect 21723 44036 21779 44038
rect 21803 44036 21859 44038
rect 21563 43002 21619 43004
rect 21643 43002 21699 43004
rect 21723 43002 21779 43004
rect 21803 43002 21859 43004
rect 21563 42950 21609 43002
rect 21609 42950 21619 43002
rect 21643 42950 21673 43002
rect 21673 42950 21685 43002
rect 21685 42950 21699 43002
rect 21723 42950 21737 43002
rect 21737 42950 21749 43002
rect 21749 42950 21779 43002
rect 21803 42950 21813 43002
rect 21813 42950 21859 43002
rect 21563 42948 21619 42950
rect 21643 42948 21699 42950
rect 21723 42948 21779 42950
rect 21803 42948 21859 42950
rect 21563 41914 21619 41916
rect 21643 41914 21699 41916
rect 21723 41914 21779 41916
rect 21803 41914 21859 41916
rect 21563 41862 21609 41914
rect 21609 41862 21619 41914
rect 21643 41862 21673 41914
rect 21673 41862 21685 41914
rect 21685 41862 21699 41914
rect 21723 41862 21737 41914
rect 21737 41862 21749 41914
rect 21749 41862 21779 41914
rect 21803 41862 21813 41914
rect 21813 41862 21859 41914
rect 21563 41860 21619 41862
rect 21643 41860 21699 41862
rect 21723 41860 21779 41862
rect 21803 41860 21859 41862
rect 21563 40826 21619 40828
rect 21643 40826 21699 40828
rect 21723 40826 21779 40828
rect 21803 40826 21859 40828
rect 21563 40774 21609 40826
rect 21609 40774 21619 40826
rect 21643 40774 21673 40826
rect 21673 40774 21685 40826
rect 21685 40774 21699 40826
rect 21723 40774 21737 40826
rect 21737 40774 21749 40826
rect 21749 40774 21779 40826
rect 21803 40774 21813 40826
rect 21813 40774 21859 40826
rect 21563 40772 21619 40774
rect 21643 40772 21699 40774
rect 21723 40772 21779 40774
rect 21803 40772 21859 40774
rect 21563 39738 21619 39740
rect 21643 39738 21699 39740
rect 21723 39738 21779 39740
rect 21803 39738 21859 39740
rect 21563 39686 21609 39738
rect 21609 39686 21619 39738
rect 21643 39686 21673 39738
rect 21673 39686 21685 39738
rect 21685 39686 21699 39738
rect 21723 39686 21737 39738
rect 21737 39686 21749 39738
rect 21749 39686 21779 39738
rect 21803 39686 21813 39738
rect 21813 39686 21859 39738
rect 21563 39684 21619 39686
rect 21643 39684 21699 39686
rect 21723 39684 21779 39686
rect 21803 39684 21859 39686
rect 21563 38650 21619 38652
rect 21643 38650 21699 38652
rect 21723 38650 21779 38652
rect 21803 38650 21859 38652
rect 21563 38598 21609 38650
rect 21609 38598 21619 38650
rect 21643 38598 21673 38650
rect 21673 38598 21685 38650
rect 21685 38598 21699 38650
rect 21723 38598 21737 38650
rect 21737 38598 21749 38650
rect 21749 38598 21779 38650
rect 21803 38598 21813 38650
rect 21813 38598 21859 38650
rect 21563 38596 21619 38598
rect 21643 38596 21699 38598
rect 21723 38596 21779 38598
rect 21803 38596 21859 38598
rect 21563 37562 21619 37564
rect 21643 37562 21699 37564
rect 21723 37562 21779 37564
rect 21803 37562 21859 37564
rect 21563 37510 21609 37562
rect 21609 37510 21619 37562
rect 21643 37510 21673 37562
rect 21673 37510 21685 37562
rect 21685 37510 21699 37562
rect 21723 37510 21737 37562
rect 21737 37510 21749 37562
rect 21749 37510 21779 37562
rect 21803 37510 21813 37562
rect 21813 37510 21859 37562
rect 21563 37508 21619 37510
rect 21643 37508 21699 37510
rect 21723 37508 21779 37510
rect 21803 37508 21859 37510
rect 21563 36474 21619 36476
rect 21643 36474 21699 36476
rect 21723 36474 21779 36476
rect 21803 36474 21859 36476
rect 21563 36422 21609 36474
rect 21609 36422 21619 36474
rect 21643 36422 21673 36474
rect 21673 36422 21685 36474
rect 21685 36422 21699 36474
rect 21723 36422 21737 36474
rect 21737 36422 21749 36474
rect 21749 36422 21779 36474
rect 21803 36422 21813 36474
rect 21813 36422 21859 36474
rect 21563 36420 21619 36422
rect 21643 36420 21699 36422
rect 21723 36420 21779 36422
rect 21803 36420 21859 36422
rect 26715 47898 26771 47900
rect 26795 47898 26851 47900
rect 26875 47898 26931 47900
rect 26955 47898 27011 47900
rect 26715 47846 26761 47898
rect 26761 47846 26771 47898
rect 26795 47846 26825 47898
rect 26825 47846 26837 47898
rect 26837 47846 26851 47898
rect 26875 47846 26889 47898
rect 26889 47846 26901 47898
rect 26901 47846 26931 47898
rect 26955 47846 26965 47898
rect 26965 47846 27011 47898
rect 26715 47844 26771 47846
rect 26795 47844 26851 47846
rect 26875 47844 26931 47846
rect 26955 47844 27011 47846
rect 26715 46810 26771 46812
rect 26795 46810 26851 46812
rect 26875 46810 26931 46812
rect 26955 46810 27011 46812
rect 26715 46758 26761 46810
rect 26761 46758 26771 46810
rect 26795 46758 26825 46810
rect 26825 46758 26837 46810
rect 26837 46758 26851 46810
rect 26875 46758 26889 46810
rect 26889 46758 26901 46810
rect 26901 46758 26931 46810
rect 26955 46758 26965 46810
rect 26965 46758 27011 46810
rect 26715 46756 26771 46758
rect 26795 46756 26851 46758
rect 26875 46756 26931 46758
rect 26955 46756 27011 46758
rect 21563 35386 21619 35388
rect 21643 35386 21699 35388
rect 21723 35386 21779 35388
rect 21803 35386 21859 35388
rect 21563 35334 21609 35386
rect 21609 35334 21619 35386
rect 21643 35334 21673 35386
rect 21673 35334 21685 35386
rect 21685 35334 21699 35386
rect 21723 35334 21737 35386
rect 21737 35334 21749 35386
rect 21749 35334 21779 35386
rect 21803 35334 21813 35386
rect 21813 35334 21859 35386
rect 21563 35332 21619 35334
rect 21643 35332 21699 35334
rect 21723 35332 21779 35334
rect 21803 35332 21859 35334
rect 21563 34298 21619 34300
rect 21643 34298 21699 34300
rect 21723 34298 21779 34300
rect 21803 34298 21859 34300
rect 21563 34246 21609 34298
rect 21609 34246 21619 34298
rect 21643 34246 21673 34298
rect 21673 34246 21685 34298
rect 21685 34246 21699 34298
rect 21723 34246 21737 34298
rect 21737 34246 21749 34298
rect 21749 34246 21779 34298
rect 21803 34246 21813 34298
rect 21813 34246 21859 34298
rect 21563 34244 21619 34246
rect 21643 34244 21699 34246
rect 21723 34244 21779 34246
rect 21803 34244 21859 34246
rect 21563 33210 21619 33212
rect 21643 33210 21699 33212
rect 21723 33210 21779 33212
rect 21803 33210 21859 33212
rect 21563 33158 21609 33210
rect 21609 33158 21619 33210
rect 21643 33158 21673 33210
rect 21673 33158 21685 33210
rect 21685 33158 21699 33210
rect 21723 33158 21737 33210
rect 21737 33158 21749 33210
rect 21749 33158 21779 33210
rect 21803 33158 21813 33210
rect 21813 33158 21859 33210
rect 21563 33156 21619 33158
rect 21643 33156 21699 33158
rect 21723 33156 21779 33158
rect 21803 33156 21859 33158
rect 21563 32122 21619 32124
rect 21643 32122 21699 32124
rect 21723 32122 21779 32124
rect 21803 32122 21859 32124
rect 21563 32070 21609 32122
rect 21609 32070 21619 32122
rect 21643 32070 21673 32122
rect 21673 32070 21685 32122
rect 21685 32070 21699 32122
rect 21723 32070 21737 32122
rect 21737 32070 21749 32122
rect 21749 32070 21779 32122
rect 21803 32070 21813 32122
rect 21813 32070 21859 32122
rect 21563 32068 21619 32070
rect 21643 32068 21699 32070
rect 21723 32068 21779 32070
rect 21803 32068 21859 32070
rect 21563 31034 21619 31036
rect 21643 31034 21699 31036
rect 21723 31034 21779 31036
rect 21803 31034 21859 31036
rect 21563 30982 21609 31034
rect 21609 30982 21619 31034
rect 21643 30982 21673 31034
rect 21673 30982 21685 31034
rect 21685 30982 21699 31034
rect 21723 30982 21737 31034
rect 21737 30982 21749 31034
rect 21749 30982 21779 31034
rect 21803 30982 21813 31034
rect 21813 30982 21859 31034
rect 21563 30980 21619 30982
rect 21643 30980 21699 30982
rect 21723 30980 21779 30982
rect 21803 30980 21859 30982
rect 21563 29946 21619 29948
rect 21643 29946 21699 29948
rect 21723 29946 21779 29948
rect 21803 29946 21859 29948
rect 21563 29894 21609 29946
rect 21609 29894 21619 29946
rect 21643 29894 21673 29946
rect 21673 29894 21685 29946
rect 21685 29894 21699 29946
rect 21723 29894 21737 29946
rect 21737 29894 21749 29946
rect 21749 29894 21779 29946
rect 21803 29894 21813 29946
rect 21813 29894 21859 29946
rect 21563 29892 21619 29894
rect 21643 29892 21699 29894
rect 21723 29892 21779 29894
rect 21803 29892 21859 29894
rect 21563 28858 21619 28860
rect 21643 28858 21699 28860
rect 21723 28858 21779 28860
rect 21803 28858 21859 28860
rect 21563 28806 21609 28858
rect 21609 28806 21619 28858
rect 21643 28806 21673 28858
rect 21673 28806 21685 28858
rect 21685 28806 21699 28858
rect 21723 28806 21737 28858
rect 21737 28806 21749 28858
rect 21749 28806 21779 28858
rect 21803 28806 21813 28858
rect 21813 28806 21859 28858
rect 21563 28804 21619 28806
rect 21643 28804 21699 28806
rect 21723 28804 21779 28806
rect 21803 28804 21859 28806
rect 21563 27770 21619 27772
rect 21643 27770 21699 27772
rect 21723 27770 21779 27772
rect 21803 27770 21859 27772
rect 21563 27718 21609 27770
rect 21609 27718 21619 27770
rect 21643 27718 21673 27770
rect 21673 27718 21685 27770
rect 21685 27718 21699 27770
rect 21723 27718 21737 27770
rect 21737 27718 21749 27770
rect 21749 27718 21779 27770
rect 21803 27718 21813 27770
rect 21813 27718 21859 27770
rect 21563 27716 21619 27718
rect 21643 27716 21699 27718
rect 21723 27716 21779 27718
rect 21803 27716 21859 27718
rect 21563 26682 21619 26684
rect 21643 26682 21699 26684
rect 21723 26682 21779 26684
rect 21803 26682 21859 26684
rect 21563 26630 21609 26682
rect 21609 26630 21619 26682
rect 21643 26630 21673 26682
rect 21673 26630 21685 26682
rect 21685 26630 21699 26682
rect 21723 26630 21737 26682
rect 21737 26630 21749 26682
rect 21749 26630 21779 26682
rect 21803 26630 21813 26682
rect 21813 26630 21859 26682
rect 21563 26628 21619 26630
rect 21643 26628 21699 26630
rect 21723 26628 21779 26630
rect 21803 26628 21859 26630
rect 21563 25594 21619 25596
rect 21643 25594 21699 25596
rect 21723 25594 21779 25596
rect 21803 25594 21859 25596
rect 21563 25542 21609 25594
rect 21609 25542 21619 25594
rect 21643 25542 21673 25594
rect 21673 25542 21685 25594
rect 21685 25542 21699 25594
rect 21723 25542 21737 25594
rect 21737 25542 21749 25594
rect 21749 25542 21779 25594
rect 21803 25542 21813 25594
rect 21813 25542 21859 25594
rect 21563 25540 21619 25542
rect 21643 25540 21699 25542
rect 21723 25540 21779 25542
rect 21803 25540 21859 25542
rect 21563 24506 21619 24508
rect 21643 24506 21699 24508
rect 21723 24506 21779 24508
rect 21803 24506 21859 24508
rect 21563 24454 21609 24506
rect 21609 24454 21619 24506
rect 21643 24454 21673 24506
rect 21673 24454 21685 24506
rect 21685 24454 21699 24506
rect 21723 24454 21737 24506
rect 21737 24454 21749 24506
rect 21749 24454 21779 24506
rect 21803 24454 21813 24506
rect 21813 24454 21859 24506
rect 21563 24452 21619 24454
rect 21643 24452 21699 24454
rect 21723 24452 21779 24454
rect 21803 24452 21859 24454
rect 21563 23418 21619 23420
rect 21643 23418 21699 23420
rect 21723 23418 21779 23420
rect 21803 23418 21859 23420
rect 21563 23366 21609 23418
rect 21609 23366 21619 23418
rect 21643 23366 21673 23418
rect 21673 23366 21685 23418
rect 21685 23366 21699 23418
rect 21723 23366 21737 23418
rect 21737 23366 21749 23418
rect 21749 23366 21779 23418
rect 21803 23366 21813 23418
rect 21813 23366 21859 23418
rect 21563 23364 21619 23366
rect 21643 23364 21699 23366
rect 21723 23364 21779 23366
rect 21803 23364 21859 23366
rect 21563 22330 21619 22332
rect 21643 22330 21699 22332
rect 21723 22330 21779 22332
rect 21803 22330 21859 22332
rect 21563 22278 21609 22330
rect 21609 22278 21619 22330
rect 21643 22278 21673 22330
rect 21673 22278 21685 22330
rect 21685 22278 21699 22330
rect 21723 22278 21737 22330
rect 21737 22278 21749 22330
rect 21749 22278 21779 22330
rect 21803 22278 21813 22330
rect 21813 22278 21859 22330
rect 21563 22276 21619 22278
rect 21643 22276 21699 22278
rect 21723 22276 21779 22278
rect 21803 22276 21859 22278
rect 21563 21242 21619 21244
rect 21643 21242 21699 21244
rect 21723 21242 21779 21244
rect 21803 21242 21859 21244
rect 21563 21190 21609 21242
rect 21609 21190 21619 21242
rect 21643 21190 21673 21242
rect 21673 21190 21685 21242
rect 21685 21190 21699 21242
rect 21723 21190 21737 21242
rect 21737 21190 21749 21242
rect 21749 21190 21779 21242
rect 21803 21190 21813 21242
rect 21813 21190 21859 21242
rect 21563 21188 21619 21190
rect 21643 21188 21699 21190
rect 21723 21188 21779 21190
rect 21803 21188 21859 21190
rect 21563 20154 21619 20156
rect 21643 20154 21699 20156
rect 21723 20154 21779 20156
rect 21803 20154 21859 20156
rect 21563 20102 21609 20154
rect 21609 20102 21619 20154
rect 21643 20102 21673 20154
rect 21673 20102 21685 20154
rect 21685 20102 21699 20154
rect 21723 20102 21737 20154
rect 21737 20102 21749 20154
rect 21749 20102 21779 20154
rect 21803 20102 21813 20154
rect 21813 20102 21859 20154
rect 21563 20100 21619 20102
rect 21643 20100 21699 20102
rect 21723 20100 21779 20102
rect 21803 20100 21859 20102
rect 21563 19066 21619 19068
rect 21643 19066 21699 19068
rect 21723 19066 21779 19068
rect 21803 19066 21859 19068
rect 21563 19014 21609 19066
rect 21609 19014 21619 19066
rect 21643 19014 21673 19066
rect 21673 19014 21685 19066
rect 21685 19014 21699 19066
rect 21723 19014 21737 19066
rect 21737 19014 21749 19066
rect 21749 19014 21779 19066
rect 21803 19014 21813 19066
rect 21813 19014 21859 19066
rect 21563 19012 21619 19014
rect 21643 19012 21699 19014
rect 21723 19012 21779 19014
rect 21803 19012 21859 19014
rect 21563 17978 21619 17980
rect 21643 17978 21699 17980
rect 21723 17978 21779 17980
rect 21803 17978 21859 17980
rect 21563 17926 21609 17978
rect 21609 17926 21619 17978
rect 21643 17926 21673 17978
rect 21673 17926 21685 17978
rect 21685 17926 21699 17978
rect 21723 17926 21737 17978
rect 21737 17926 21749 17978
rect 21749 17926 21779 17978
rect 21803 17926 21813 17978
rect 21813 17926 21859 17978
rect 21563 17924 21619 17926
rect 21643 17924 21699 17926
rect 21723 17924 21779 17926
rect 21803 17924 21859 17926
rect 21563 16890 21619 16892
rect 21643 16890 21699 16892
rect 21723 16890 21779 16892
rect 21803 16890 21859 16892
rect 21563 16838 21609 16890
rect 21609 16838 21619 16890
rect 21643 16838 21673 16890
rect 21673 16838 21685 16890
rect 21685 16838 21699 16890
rect 21723 16838 21737 16890
rect 21737 16838 21749 16890
rect 21749 16838 21779 16890
rect 21803 16838 21813 16890
rect 21813 16838 21859 16890
rect 21563 16836 21619 16838
rect 21643 16836 21699 16838
rect 21723 16836 21779 16838
rect 21803 16836 21859 16838
rect 21563 15802 21619 15804
rect 21643 15802 21699 15804
rect 21723 15802 21779 15804
rect 21803 15802 21859 15804
rect 21563 15750 21609 15802
rect 21609 15750 21619 15802
rect 21643 15750 21673 15802
rect 21673 15750 21685 15802
rect 21685 15750 21699 15802
rect 21723 15750 21737 15802
rect 21737 15750 21749 15802
rect 21749 15750 21779 15802
rect 21803 15750 21813 15802
rect 21813 15750 21859 15802
rect 21563 15748 21619 15750
rect 21643 15748 21699 15750
rect 21723 15748 21779 15750
rect 21803 15748 21859 15750
rect 21563 14714 21619 14716
rect 21643 14714 21699 14716
rect 21723 14714 21779 14716
rect 21803 14714 21859 14716
rect 21563 14662 21609 14714
rect 21609 14662 21619 14714
rect 21643 14662 21673 14714
rect 21673 14662 21685 14714
rect 21685 14662 21699 14714
rect 21723 14662 21737 14714
rect 21737 14662 21749 14714
rect 21749 14662 21779 14714
rect 21803 14662 21813 14714
rect 21813 14662 21859 14714
rect 21563 14660 21619 14662
rect 21643 14660 21699 14662
rect 21723 14660 21779 14662
rect 21803 14660 21859 14662
rect 21563 13626 21619 13628
rect 21643 13626 21699 13628
rect 21723 13626 21779 13628
rect 21803 13626 21859 13628
rect 21563 13574 21609 13626
rect 21609 13574 21619 13626
rect 21643 13574 21673 13626
rect 21673 13574 21685 13626
rect 21685 13574 21699 13626
rect 21723 13574 21737 13626
rect 21737 13574 21749 13626
rect 21749 13574 21779 13626
rect 21803 13574 21813 13626
rect 21813 13574 21859 13626
rect 21563 13572 21619 13574
rect 21643 13572 21699 13574
rect 21723 13572 21779 13574
rect 21803 13572 21859 13574
rect 21563 12538 21619 12540
rect 21643 12538 21699 12540
rect 21723 12538 21779 12540
rect 21803 12538 21859 12540
rect 21563 12486 21609 12538
rect 21609 12486 21619 12538
rect 21643 12486 21673 12538
rect 21673 12486 21685 12538
rect 21685 12486 21699 12538
rect 21723 12486 21737 12538
rect 21737 12486 21749 12538
rect 21749 12486 21779 12538
rect 21803 12486 21813 12538
rect 21813 12486 21859 12538
rect 21563 12484 21619 12486
rect 21643 12484 21699 12486
rect 21723 12484 21779 12486
rect 21803 12484 21859 12486
rect 21563 11450 21619 11452
rect 21643 11450 21699 11452
rect 21723 11450 21779 11452
rect 21803 11450 21859 11452
rect 21563 11398 21609 11450
rect 21609 11398 21619 11450
rect 21643 11398 21673 11450
rect 21673 11398 21685 11450
rect 21685 11398 21699 11450
rect 21723 11398 21737 11450
rect 21737 11398 21749 11450
rect 21749 11398 21779 11450
rect 21803 11398 21813 11450
rect 21813 11398 21859 11450
rect 21563 11396 21619 11398
rect 21643 11396 21699 11398
rect 21723 11396 21779 11398
rect 21803 11396 21859 11398
rect 21563 10362 21619 10364
rect 21643 10362 21699 10364
rect 21723 10362 21779 10364
rect 21803 10362 21859 10364
rect 21563 10310 21609 10362
rect 21609 10310 21619 10362
rect 21643 10310 21673 10362
rect 21673 10310 21685 10362
rect 21685 10310 21699 10362
rect 21723 10310 21737 10362
rect 21737 10310 21749 10362
rect 21749 10310 21779 10362
rect 21803 10310 21813 10362
rect 21813 10310 21859 10362
rect 21563 10308 21619 10310
rect 21643 10308 21699 10310
rect 21723 10308 21779 10310
rect 21803 10308 21859 10310
rect 26715 45722 26771 45724
rect 26795 45722 26851 45724
rect 26875 45722 26931 45724
rect 26955 45722 27011 45724
rect 26715 45670 26761 45722
rect 26761 45670 26771 45722
rect 26795 45670 26825 45722
rect 26825 45670 26837 45722
rect 26837 45670 26851 45722
rect 26875 45670 26889 45722
rect 26889 45670 26901 45722
rect 26901 45670 26931 45722
rect 26955 45670 26965 45722
rect 26965 45670 27011 45722
rect 26715 45668 26771 45670
rect 26795 45668 26851 45670
rect 26875 45668 26931 45670
rect 26955 45668 27011 45670
rect 26715 44634 26771 44636
rect 26795 44634 26851 44636
rect 26875 44634 26931 44636
rect 26955 44634 27011 44636
rect 26715 44582 26761 44634
rect 26761 44582 26771 44634
rect 26795 44582 26825 44634
rect 26825 44582 26837 44634
rect 26837 44582 26851 44634
rect 26875 44582 26889 44634
rect 26889 44582 26901 44634
rect 26901 44582 26931 44634
rect 26955 44582 26965 44634
rect 26965 44582 27011 44634
rect 26715 44580 26771 44582
rect 26795 44580 26851 44582
rect 26875 44580 26931 44582
rect 26955 44580 27011 44582
rect 21563 9274 21619 9276
rect 21643 9274 21699 9276
rect 21723 9274 21779 9276
rect 21803 9274 21859 9276
rect 21563 9222 21609 9274
rect 21609 9222 21619 9274
rect 21643 9222 21673 9274
rect 21673 9222 21685 9274
rect 21685 9222 21699 9274
rect 21723 9222 21737 9274
rect 21737 9222 21749 9274
rect 21749 9222 21779 9274
rect 21803 9222 21813 9274
rect 21813 9222 21859 9274
rect 21563 9220 21619 9222
rect 21643 9220 21699 9222
rect 21723 9220 21779 9222
rect 21803 9220 21859 9222
rect 21563 8186 21619 8188
rect 21643 8186 21699 8188
rect 21723 8186 21779 8188
rect 21803 8186 21859 8188
rect 21563 8134 21609 8186
rect 21609 8134 21619 8186
rect 21643 8134 21673 8186
rect 21673 8134 21685 8186
rect 21685 8134 21699 8186
rect 21723 8134 21737 8186
rect 21737 8134 21749 8186
rect 21749 8134 21779 8186
rect 21803 8134 21813 8186
rect 21813 8134 21859 8186
rect 21563 8132 21619 8134
rect 21643 8132 21699 8134
rect 21723 8132 21779 8134
rect 21803 8132 21859 8134
rect 21563 7098 21619 7100
rect 21643 7098 21699 7100
rect 21723 7098 21779 7100
rect 21803 7098 21859 7100
rect 21563 7046 21609 7098
rect 21609 7046 21619 7098
rect 21643 7046 21673 7098
rect 21673 7046 21685 7098
rect 21685 7046 21699 7098
rect 21723 7046 21737 7098
rect 21737 7046 21749 7098
rect 21749 7046 21779 7098
rect 21803 7046 21813 7098
rect 21813 7046 21859 7098
rect 21563 7044 21619 7046
rect 21643 7044 21699 7046
rect 21723 7044 21779 7046
rect 21803 7044 21859 7046
rect 21563 6010 21619 6012
rect 21643 6010 21699 6012
rect 21723 6010 21779 6012
rect 21803 6010 21859 6012
rect 21563 5958 21609 6010
rect 21609 5958 21619 6010
rect 21643 5958 21673 6010
rect 21673 5958 21685 6010
rect 21685 5958 21699 6010
rect 21723 5958 21737 6010
rect 21737 5958 21749 6010
rect 21749 5958 21779 6010
rect 21803 5958 21813 6010
rect 21813 5958 21859 6010
rect 21563 5956 21619 5958
rect 21643 5956 21699 5958
rect 21723 5956 21779 5958
rect 21803 5956 21859 5958
rect 21563 4922 21619 4924
rect 21643 4922 21699 4924
rect 21723 4922 21779 4924
rect 21803 4922 21859 4924
rect 21563 4870 21609 4922
rect 21609 4870 21619 4922
rect 21643 4870 21673 4922
rect 21673 4870 21685 4922
rect 21685 4870 21699 4922
rect 21723 4870 21737 4922
rect 21737 4870 21749 4922
rect 21749 4870 21779 4922
rect 21803 4870 21813 4922
rect 21813 4870 21859 4922
rect 21563 4868 21619 4870
rect 21643 4868 21699 4870
rect 21723 4868 21779 4870
rect 21803 4868 21859 4870
rect 21563 3834 21619 3836
rect 21643 3834 21699 3836
rect 21723 3834 21779 3836
rect 21803 3834 21859 3836
rect 21563 3782 21609 3834
rect 21609 3782 21619 3834
rect 21643 3782 21673 3834
rect 21673 3782 21685 3834
rect 21685 3782 21699 3834
rect 21723 3782 21737 3834
rect 21737 3782 21749 3834
rect 21749 3782 21779 3834
rect 21803 3782 21813 3834
rect 21813 3782 21859 3834
rect 21563 3780 21619 3782
rect 21643 3780 21699 3782
rect 21723 3780 21779 3782
rect 21803 3780 21859 3782
rect 21563 2746 21619 2748
rect 21643 2746 21699 2748
rect 21723 2746 21779 2748
rect 21803 2746 21859 2748
rect 21563 2694 21609 2746
rect 21609 2694 21619 2746
rect 21643 2694 21673 2746
rect 21673 2694 21685 2746
rect 21685 2694 21699 2746
rect 21723 2694 21737 2746
rect 21737 2694 21749 2746
rect 21749 2694 21779 2746
rect 21803 2694 21813 2746
rect 21813 2694 21859 2746
rect 21563 2692 21619 2694
rect 21643 2692 21699 2694
rect 21723 2692 21779 2694
rect 21803 2692 21859 2694
rect 21563 1658 21619 1660
rect 21643 1658 21699 1660
rect 21723 1658 21779 1660
rect 21803 1658 21859 1660
rect 21563 1606 21609 1658
rect 21609 1606 21619 1658
rect 21643 1606 21673 1658
rect 21673 1606 21685 1658
rect 21685 1606 21699 1658
rect 21723 1606 21737 1658
rect 21737 1606 21749 1658
rect 21749 1606 21779 1658
rect 21803 1606 21813 1658
rect 21813 1606 21859 1658
rect 21563 1604 21619 1606
rect 21643 1604 21699 1606
rect 21723 1604 21779 1606
rect 21803 1604 21859 1606
rect 26715 43546 26771 43548
rect 26795 43546 26851 43548
rect 26875 43546 26931 43548
rect 26955 43546 27011 43548
rect 26715 43494 26761 43546
rect 26761 43494 26771 43546
rect 26795 43494 26825 43546
rect 26825 43494 26837 43546
rect 26837 43494 26851 43546
rect 26875 43494 26889 43546
rect 26889 43494 26901 43546
rect 26901 43494 26931 43546
rect 26955 43494 26965 43546
rect 26965 43494 27011 43546
rect 26715 43492 26771 43494
rect 26795 43492 26851 43494
rect 26875 43492 26931 43494
rect 26955 43492 27011 43494
rect 26715 42458 26771 42460
rect 26795 42458 26851 42460
rect 26875 42458 26931 42460
rect 26955 42458 27011 42460
rect 26715 42406 26761 42458
rect 26761 42406 26771 42458
rect 26795 42406 26825 42458
rect 26825 42406 26837 42458
rect 26837 42406 26851 42458
rect 26875 42406 26889 42458
rect 26889 42406 26901 42458
rect 26901 42406 26931 42458
rect 26955 42406 26965 42458
rect 26965 42406 27011 42458
rect 26715 42404 26771 42406
rect 26795 42404 26851 42406
rect 26875 42404 26931 42406
rect 26955 42404 27011 42406
rect 26715 41370 26771 41372
rect 26795 41370 26851 41372
rect 26875 41370 26931 41372
rect 26955 41370 27011 41372
rect 26715 41318 26761 41370
rect 26761 41318 26771 41370
rect 26795 41318 26825 41370
rect 26825 41318 26837 41370
rect 26837 41318 26851 41370
rect 26875 41318 26889 41370
rect 26889 41318 26901 41370
rect 26901 41318 26931 41370
rect 26955 41318 26965 41370
rect 26965 41318 27011 41370
rect 26715 41316 26771 41318
rect 26795 41316 26851 41318
rect 26875 41316 26931 41318
rect 26955 41316 27011 41318
rect 26715 40282 26771 40284
rect 26795 40282 26851 40284
rect 26875 40282 26931 40284
rect 26955 40282 27011 40284
rect 26715 40230 26761 40282
rect 26761 40230 26771 40282
rect 26795 40230 26825 40282
rect 26825 40230 26837 40282
rect 26837 40230 26851 40282
rect 26875 40230 26889 40282
rect 26889 40230 26901 40282
rect 26901 40230 26931 40282
rect 26955 40230 26965 40282
rect 26965 40230 27011 40282
rect 26715 40228 26771 40230
rect 26795 40228 26851 40230
rect 26875 40228 26931 40230
rect 26955 40228 27011 40230
rect 26715 39194 26771 39196
rect 26795 39194 26851 39196
rect 26875 39194 26931 39196
rect 26955 39194 27011 39196
rect 26715 39142 26761 39194
rect 26761 39142 26771 39194
rect 26795 39142 26825 39194
rect 26825 39142 26837 39194
rect 26837 39142 26851 39194
rect 26875 39142 26889 39194
rect 26889 39142 26901 39194
rect 26901 39142 26931 39194
rect 26955 39142 26965 39194
rect 26965 39142 27011 39194
rect 26715 39140 26771 39142
rect 26795 39140 26851 39142
rect 26875 39140 26931 39142
rect 26955 39140 27011 39142
rect 26715 38106 26771 38108
rect 26795 38106 26851 38108
rect 26875 38106 26931 38108
rect 26955 38106 27011 38108
rect 26715 38054 26761 38106
rect 26761 38054 26771 38106
rect 26795 38054 26825 38106
rect 26825 38054 26837 38106
rect 26837 38054 26851 38106
rect 26875 38054 26889 38106
rect 26889 38054 26901 38106
rect 26901 38054 26931 38106
rect 26955 38054 26965 38106
rect 26965 38054 27011 38106
rect 26715 38052 26771 38054
rect 26795 38052 26851 38054
rect 26875 38052 26931 38054
rect 26955 38052 27011 38054
rect 26715 37018 26771 37020
rect 26795 37018 26851 37020
rect 26875 37018 26931 37020
rect 26955 37018 27011 37020
rect 26715 36966 26761 37018
rect 26761 36966 26771 37018
rect 26795 36966 26825 37018
rect 26825 36966 26837 37018
rect 26837 36966 26851 37018
rect 26875 36966 26889 37018
rect 26889 36966 26901 37018
rect 26901 36966 26931 37018
rect 26955 36966 26965 37018
rect 26965 36966 27011 37018
rect 26715 36964 26771 36966
rect 26795 36964 26851 36966
rect 26875 36964 26931 36966
rect 26955 36964 27011 36966
rect 26715 35930 26771 35932
rect 26795 35930 26851 35932
rect 26875 35930 26931 35932
rect 26955 35930 27011 35932
rect 26715 35878 26761 35930
rect 26761 35878 26771 35930
rect 26795 35878 26825 35930
rect 26825 35878 26837 35930
rect 26837 35878 26851 35930
rect 26875 35878 26889 35930
rect 26889 35878 26901 35930
rect 26901 35878 26931 35930
rect 26955 35878 26965 35930
rect 26965 35878 27011 35930
rect 26715 35876 26771 35878
rect 26795 35876 26851 35878
rect 26875 35876 26931 35878
rect 26955 35876 27011 35878
rect 26715 34842 26771 34844
rect 26795 34842 26851 34844
rect 26875 34842 26931 34844
rect 26955 34842 27011 34844
rect 26715 34790 26761 34842
rect 26761 34790 26771 34842
rect 26795 34790 26825 34842
rect 26825 34790 26837 34842
rect 26837 34790 26851 34842
rect 26875 34790 26889 34842
rect 26889 34790 26901 34842
rect 26901 34790 26931 34842
rect 26955 34790 26965 34842
rect 26965 34790 27011 34842
rect 26715 34788 26771 34790
rect 26795 34788 26851 34790
rect 26875 34788 26931 34790
rect 26955 34788 27011 34790
rect 26715 33754 26771 33756
rect 26795 33754 26851 33756
rect 26875 33754 26931 33756
rect 26955 33754 27011 33756
rect 26715 33702 26761 33754
rect 26761 33702 26771 33754
rect 26795 33702 26825 33754
rect 26825 33702 26837 33754
rect 26837 33702 26851 33754
rect 26875 33702 26889 33754
rect 26889 33702 26901 33754
rect 26901 33702 26931 33754
rect 26955 33702 26965 33754
rect 26965 33702 27011 33754
rect 26715 33700 26771 33702
rect 26795 33700 26851 33702
rect 26875 33700 26931 33702
rect 26955 33700 27011 33702
rect 26715 32666 26771 32668
rect 26795 32666 26851 32668
rect 26875 32666 26931 32668
rect 26955 32666 27011 32668
rect 26715 32614 26761 32666
rect 26761 32614 26771 32666
rect 26795 32614 26825 32666
rect 26825 32614 26837 32666
rect 26837 32614 26851 32666
rect 26875 32614 26889 32666
rect 26889 32614 26901 32666
rect 26901 32614 26931 32666
rect 26955 32614 26965 32666
rect 26965 32614 27011 32666
rect 26715 32612 26771 32614
rect 26795 32612 26851 32614
rect 26875 32612 26931 32614
rect 26955 32612 27011 32614
rect 26715 31578 26771 31580
rect 26795 31578 26851 31580
rect 26875 31578 26931 31580
rect 26955 31578 27011 31580
rect 26715 31526 26761 31578
rect 26761 31526 26771 31578
rect 26795 31526 26825 31578
rect 26825 31526 26837 31578
rect 26837 31526 26851 31578
rect 26875 31526 26889 31578
rect 26889 31526 26901 31578
rect 26901 31526 26931 31578
rect 26955 31526 26965 31578
rect 26965 31526 27011 31578
rect 26715 31524 26771 31526
rect 26795 31524 26851 31526
rect 26875 31524 26931 31526
rect 26955 31524 27011 31526
rect 21563 570 21619 572
rect 21643 570 21699 572
rect 21723 570 21779 572
rect 21803 570 21859 572
rect 21563 518 21609 570
rect 21609 518 21619 570
rect 21643 518 21673 570
rect 21673 518 21685 570
rect 21685 518 21699 570
rect 21723 518 21737 570
rect 21737 518 21749 570
rect 21749 518 21779 570
rect 21803 518 21813 570
rect 21813 518 21859 570
rect 21563 516 21619 518
rect 21643 516 21699 518
rect 21723 516 21779 518
rect 21803 516 21859 518
rect 26715 30490 26771 30492
rect 26795 30490 26851 30492
rect 26875 30490 26931 30492
rect 26955 30490 27011 30492
rect 26715 30438 26761 30490
rect 26761 30438 26771 30490
rect 26795 30438 26825 30490
rect 26825 30438 26837 30490
rect 26837 30438 26851 30490
rect 26875 30438 26889 30490
rect 26889 30438 26901 30490
rect 26901 30438 26931 30490
rect 26955 30438 26965 30490
rect 26965 30438 27011 30490
rect 26715 30436 26771 30438
rect 26795 30436 26851 30438
rect 26875 30436 26931 30438
rect 26955 30436 27011 30438
rect 26715 29402 26771 29404
rect 26795 29402 26851 29404
rect 26875 29402 26931 29404
rect 26955 29402 27011 29404
rect 26715 29350 26761 29402
rect 26761 29350 26771 29402
rect 26795 29350 26825 29402
rect 26825 29350 26837 29402
rect 26837 29350 26851 29402
rect 26875 29350 26889 29402
rect 26889 29350 26901 29402
rect 26901 29350 26931 29402
rect 26955 29350 26965 29402
rect 26965 29350 27011 29402
rect 26715 29348 26771 29350
rect 26795 29348 26851 29350
rect 26875 29348 26931 29350
rect 26955 29348 27011 29350
rect 26715 28314 26771 28316
rect 26795 28314 26851 28316
rect 26875 28314 26931 28316
rect 26955 28314 27011 28316
rect 26715 28262 26761 28314
rect 26761 28262 26771 28314
rect 26795 28262 26825 28314
rect 26825 28262 26837 28314
rect 26837 28262 26851 28314
rect 26875 28262 26889 28314
rect 26889 28262 26901 28314
rect 26901 28262 26931 28314
rect 26955 28262 26965 28314
rect 26965 28262 27011 28314
rect 26715 28260 26771 28262
rect 26795 28260 26851 28262
rect 26875 28260 26931 28262
rect 26955 28260 27011 28262
rect 26715 27226 26771 27228
rect 26795 27226 26851 27228
rect 26875 27226 26931 27228
rect 26955 27226 27011 27228
rect 26715 27174 26761 27226
rect 26761 27174 26771 27226
rect 26795 27174 26825 27226
rect 26825 27174 26837 27226
rect 26837 27174 26851 27226
rect 26875 27174 26889 27226
rect 26889 27174 26901 27226
rect 26901 27174 26931 27226
rect 26955 27174 26965 27226
rect 26965 27174 27011 27226
rect 26715 27172 26771 27174
rect 26795 27172 26851 27174
rect 26875 27172 26931 27174
rect 26955 27172 27011 27174
rect 26715 26138 26771 26140
rect 26795 26138 26851 26140
rect 26875 26138 26931 26140
rect 26955 26138 27011 26140
rect 26715 26086 26761 26138
rect 26761 26086 26771 26138
rect 26795 26086 26825 26138
rect 26825 26086 26837 26138
rect 26837 26086 26851 26138
rect 26875 26086 26889 26138
rect 26889 26086 26901 26138
rect 26901 26086 26931 26138
rect 26955 26086 26965 26138
rect 26965 26086 27011 26138
rect 26715 26084 26771 26086
rect 26795 26084 26851 26086
rect 26875 26084 26931 26086
rect 26955 26084 27011 26086
rect 26715 25050 26771 25052
rect 26795 25050 26851 25052
rect 26875 25050 26931 25052
rect 26955 25050 27011 25052
rect 26715 24998 26761 25050
rect 26761 24998 26771 25050
rect 26795 24998 26825 25050
rect 26825 24998 26837 25050
rect 26837 24998 26851 25050
rect 26875 24998 26889 25050
rect 26889 24998 26901 25050
rect 26901 24998 26931 25050
rect 26955 24998 26965 25050
rect 26965 24998 27011 25050
rect 26715 24996 26771 24998
rect 26795 24996 26851 24998
rect 26875 24996 26931 24998
rect 26955 24996 27011 24998
rect 26715 23962 26771 23964
rect 26795 23962 26851 23964
rect 26875 23962 26931 23964
rect 26955 23962 27011 23964
rect 26715 23910 26761 23962
rect 26761 23910 26771 23962
rect 26795 23910 26825 23962
rect 26825 23910 26837 23962
rect 26837 23910 26851 23962
rect 26875 23910 26889 23962
rect 26889 23910 26901 23962
rect 26901 23910 26931 23962
rect 26955 23910 26965 23962
rect 26965 23910 27011 23962
rect 26715 23908 26771 23910
rect 26795 23908 26851 23910
rect 26875 23908 26931 23910
rect 26955 23908 27011 23910
rect 26715 22874 26771 22876
rect 26795 22874 26851 22876
rect 26875 22874 26931 22876
rect 26955 22874 27011 22876
rect 26715 22822 26761 22874
rect 26761 22822 26771 22874
rect 26795 22822 26825 22874
rect 26825 22822 26837 22874
rect 26837 22822 26851 22874
rect 26875 22822 26889 22874
rect 26889 22822 26901 22874
rect 26901 22822 26931 22874
rect 26955 22822 26965 22874
rect 26965 22822 27011 22874
rect 26715 22820 26771 22822
rect 26795 22820 26851 22822
rect 26875 22820 26931 22822
rect 26955 22820 27011 22822
rect 26715 21786 26771 21788
rect 26795 21786 26851 21788
rect 26875 21786 26931 21788
rect 26955 21786 27011 21788
rect 26715 21734 26761 21786
rect 26761 21734 26771 21786
rect 26795 21734 26825 21786
rect 26825 21734 26837 21786
rect 26837 21734 26851 21786
rect 26875 21734 26889 21786
rect 26889 21734 26901 21786
rect 26901 21734 26931 21786
rect 26955 21734 26965 21786
rect 26965 21734 27011 21786
rect 26715 21732 26771 21734
rect 26795 21732 26851 21734
rect 26875 21732 26931 21734
rect 26955 21732 27011 21734
rect 26715 20698 26771 20700
rect 26795 20698 26851 20700
rect 26875 20698 26931 20700
rect 26955 20698 27011 20700
rect 26715 20646 26761 20698
rect 26761 20646 26771 20698
rect 26795 20646 26825 20698
rect 26825 20646 26837 20698
rect 26837 20646 26851 20698
rect 26875 20646 26889 20698
rect 26889 20646 26901 20698
rect 26901 20646 26931 20698
rect 26955 20646 26965 20698
rect 26965 20646 27011 20698
rect 26715 20644 26771 20646
rect 26795 20644 26851 20646
rect 26875 20644 26931 20646
rect 26955 20644 27011 20646
rect 26715 19610 26771 19612
rect 26795 19610 26851 19612
rect 26875 19610 26931 19612
rect 26955 19610 27011 19612
rect 26715 19558 26761 19610
rect 26761 19558 26771 19610
rect 26795 19558 26825 19610
rect 26825 19558 26837 19610
rect 26837 19558 26851 19610
rect 26875 19558 26889 19610
rect 26889 19558 26901 19610
rect 26901 19558 26931 19610
rect 26955 19558 26965 19610
rect 26965 19558 27011 19610
rect 26715 19556 26771 19558
rect 26795 19556 26851 19558
rect 26875 19556 26931 19558
rect 26955 19556 27011 19558
rect 26715 18522 26771 18524
rect 26795 18522 26851 18524
rect 26875 18522 26931 18524
rect 26955 18522 27011 18524
rect 26715 18470 26761 18522
rect 26761 18470 26771 18522
rect 26795 18470 26825 18522
rect 26825 18470 26837 18522
rect 26837 18470 26851 18522
rect 26875 18470 26889 18522
rect 26889 18470 26901 18522
rect 26901 18470 26931 18522
rect 26955 18470 26965 18522
rect 26965 18470 27011 18522
rect 26715 18468 26771 18470
rect 26795 18468 26851 18470
rect 26875 18468 26931 18470
rect 26955 18468 27011 18470
rect 26715 17434 26771 17436
rect 26795 17434 26851 17436
rect 26875 17434 26931 17436
rect 26955 17434 27011 17436
rect 26715 17382 26761 17434
rect 26761 17382 26771 17434
rect 26795 17382 26825 17434
rect 26825 17382 26837 17434
rect 26837 17382 26851 17434
rect 26875 17382 26889 17434
rect 26889 17382 26901 17434
rect 26901 17382 26931 17434
rect 26955 17382 26965 17434
rect 26965 17382 27011 17434
rect 26715 17380 26771 17382
rect 26795 17380 26851 17382
rect 26875 17380 26931 17382
rect 26955 17380 27011 17382
rect 26715 16346 26771 16348
rect 26795 16346 26851 16348
rect 26875 16346 26931 16348
rect 26955 16346 27011 16348
rect 26715 16294 26761 16346
rect 26761 16294 26771 16346
rect 26795 16294 26825 16346
rect 26825 16294 26837 16346
rect 26837 16294 26851 16346
rect 26875 16294 26889 16346
rect 26889 16294 26901 16346
rect 26901 16294 26931 16346
rect 26955 16294 26965 16346
rect 26965 16294 27011 16346
rect 26715 16292 26771 16294
rect 26795 16292 26851 16294
rect 26875 16292 26931 16294
rect 26955 16292 27011 16294
rect 26715 15258 26771 15260
rect 26795 15258 26851 15260
rect 26875 15258 26931 15260
rect 26955 15258 27011 15260
rect 26715 15206 26761 15258
rect 26761 15206 26771 15258
rect 26795 15206 26825 15258
rect 26825 15206 26837 15258
rect 26837 15206 26851 15258
rect 26875 15206 26889 15258
rect 26889 15206 26901 15258
rect 26901 15206 26931 15258
rect 26955 15206 26965 15258
rect 26965 15206 27011 15258
rect 26715 15204 26771 15206
rect 26795 15204 26851 15206
rect 26875 15204 26931 15206
rect 26955 15204 27011 15206
rect 26715 14170 26771 14172
rect 26795 14170 26851 14172
rect 26875 14170 26931 14172
rect 26955 14170 27011 14172
rect 26715 14118 26761 14170
rect 26761 14118 26771 14170
rect 26795 14118 26825 14170
rect 26825 14118 26837 14170
rect 26837 14118 26851 14170
rect 26875 14118 26889 14170
rect 26889 14118 26901 14170
rect 26901 14118 26931 14170
rect 26955 14118 26965 14170
rect 26965 14118 27011 14170
rect 26715 14116 26771 14118
rect 26795 14116 26851 14118
rect 26875 14116 26931 14118
rect 26955 14116 27011 14118
rect 26715 13082 26771 13084
rect 26795 13082 26851 13084
rect 26875 13082 26931 13084
rect 26955 13082 27011 13084
rect 26715 13030 26761 13082
rect 26761 13030 26771 13082
rect 26795 13030 26825 13082
rect 26825 13030 26837 13082
rect 26837 13030 26851 13082
rect 26875 13030 26889 13082
rect 26889 13030 26901 13082
rect 26901 13030 26931 13082
rect 26955 13030 26965 13082
rect 26965 13030 27011 13082
rect 26715 13028 26771 13030
rect 26795 13028 26851 13030
rect 26875 13028 26931 13030
rect 26955 13028 27011 13030
rect 26715 11994 26771 11996
rect 26795 11994 26851 11996
rect 26875 11994 26931 11996
rect 26955 11994 27011 11996
rect 26715 11942 26761 11994
rect 26761 11942 26771 11994
rect 26795 11942 26825 11994
rect 26825 11942 26837 11994
rect 26837 11942 26851 11994
rect 26875 11942 26889 11994
rect 26889 11942 26901 11994
rect 26901 11942 26931 11994
rect 26955 11942 26965 11994
rect 26965 11942 27011 11994
rect 26715 11940 26771 11942
rect 26795 11940 26851 11942
rect 26875 11940 26931 11942
rect 26955 11940 27011 11942
rect 26715 10906 26771 10908
rect 26795 10906 26851 10908
rect 26875 10906 26931 10908
rect 26955 10906 27011 10908
rect 26715 10854 26761 10906
rect 26761 10854 26771 10906
rect 26795 10854 26825 10906
rect 26825 10854 26837 10906
rect 26837 10854 26851 10906
rect 26875 10854 26889 10906
rect 26889 10854 26901 10906
rect 26901 10854 26931 10906
rect 26955 10854 26965 10906
rect 26965 10854 27011 10906
rect 26715 10852 26771 10854
rect 26795 10852 26851 10854
rect 26875 10852 26931 10854
rect 26955 10852 27011 10854
rect 26715 9818 26771 9820
rect 26795 9818 26851 9820
rect 26875 9818 26931 9820
rect 26955 9818 27011 9820
rect 26715 9766 26761 9818
rect 26761 9766 26771 9818
rect 26795 9766 26825 9818
rect 26825 9766 26837 9818
rect 26837 9766 26851 9818
rect 26875 9766 26889 9818
rect 26889 9766 26901 9818
rect 26901 9766 26931 9818
rect 26955 9766 26965 9818
rect 26965 9766 27011 9818
rect 26715 9764 26771 9766
rect 26795 9764 26851 9766
rect 26875 9764 26931 9766
rect 26955 9764 27011 9766
rect 26715 8730 26771 8732
rect 26795 8730 26851 8732
rect 26875 8730 26931 8732
rect 26955 8730 27011 8732
rect 26715 8678 26761 8730
rect 26761 8678 26771 8730
rect 26795 8678 26825 8730
rect 26825 8678 26837 8730
rect 26837 8678 26851 8730
rect 26875 8678 26889 8730
rect 26889 8678 26901 8730
rect 26901 8678 26931 8730
rect 26955 8678 26965 8730
rect 26965 8678 27011 8730
rect 26715 8676 26771 8678
rect 26795 8676 26851 8678
rect 26875 8676 26931 8678
rect 26955 8676 27011 8678
rect 26715 7642 26771 7644
rect 26795 7642 26851 7644
rect 26875 7642 26931 7644
rect 26955 7642 27011 7644
rect 26715 7590 26761 7642
rect 26761 7590 26771 7642
rect 26795 7590 26825 7642
rect 26825 7590 26837 7642
rect 26837 7590 26851 7642
rect 26875 7590 26889 7642
rect 26889 7590 26901 7642
rect 26901 7590 26931 7642
rect 26955 7590 26965 7642
rect 26965 7590 27011 7642
rect 26715 7588 26771 7590
rect 26795 7588 26851 7590
rect 26875 7588 26931 7590
rect 26955 7588 27011 7590
rect 26715 6554 26771 6556
rect 26795 6554 26851 6556
rect 26875 6554 26931 6556
rect 26955 6554 27011 6556
rect 26715 6502 26761 6554
rect 26761 6502 26771 6554
rect 26795 6502 26825 6554
rect 26825 6502 26837 6554
rect 26837 6502 26851 6554
rect 26875 6502 26889 6554
rect 26889 6502 26901 6554
rect 26901 6502 26931 6554
rect 26955 6502 26965 6554
rect 26965 6502 27011 6554
rect 26715 6500 26771 6502
rect 26795 6500 26851 6502
rect 26875 6500 26931 6502
rect 26955 6500 27011 6502
rect 26715 5466 26771 5468
rect 26795 5466 26851 5468
rect 26875 5466 26931 5468
rect 26955 5466 27011 5468
rect 26715 5414 26761 5466
rect 26761 5414 26771 5466
rect 26795 5414 26825 5466
rect 26825 5414 26837 5466
rect 26837 5414 26851 5466
rect 26875 5414 26889 5466
rect 26889 5414 26901 5466
rect 26901 5414 26931 5466
rect 26955 5414 26965 5466
rect 26965 5414 27011 5466
rect 26715 5412 26771 5414
rect 26795 5412 26851 5414
rect 26875 5412 26931 5414
rect 26955 5412 27011 5414
rect 26715 4378 26771 4380
rect 26795 4378 26851 4380
rect 26875 4378 26931 4380
rect 26955 4378 27011 4380
rect 26715 4326 26761 4378
rect 26761 4326 26771 4378
rect 26795 4326 26825 4378
rect 26825 4326 26837 4378
rect 26837 4326 26851 4378
rect 26875 4326 26889 4378
rect 26889 4326 26901 4378
rect 26901 4326 26931 4378
rect 26955 4326 26965 4378
rect 26965 4326 27011 4378
rect 26715 4324 26771 4326
rect 26795 4324 26851 4326
rect 26875 4324 26931 4326
rect 26955 4324 27011 4326
rect 26715 3290 26771 3292
rect 26795 3290 26851 3292
rect 26875 3290 26931 3292
rect 26955 3290 27011 3292
rect 26715 3238 26761 3290
rect 26761 3238 26771 3290
rect 26795 3238 26825 3290
rect 26825 3238 26837 3290
rect 26837 3238 26851 3290
rect 26875 3238 26889 3290
rect 26889 3238 26901 3290
rect 26901 3238 26931 3290
rect 26955 3238 26965 3290
rect 26965 3238 27011 3290
rect 26715 3236 26771 3238
rect 26795 3236 26851 3238
rect 26875 3236 26931 3238
rect 26955 3236 27011 3238
rect 26715 2202 26771 2204
rect 26795 2202 26851 2204
rect 26875 2202 26931 2204
rect 26955 2202 27011 2204
rect 26715 2150 26761 2202
rect 26761 2150 26771 2202
rect 26795 2150 26825 2202
rect 26825 2150 26837 2202
rect 26837 2150 26851 2202
rect 26875 2150 26889 2202
rect 26889 2150 26901 2202
rect 26901 2150 26931 2202
rect 26955 2150 26965 2202
rect 26965 2150 27011 2202
rect 26715 2148 26771 2150
rect 26795 2148 26851 2150
rect 26875 2148 26931 2150
rect 26955 2148 27011 2150
rect 26715 1114 26771 1116
rect 26795 1114 26851 1116
rect 26875 1114 26931 1116
rect 26955 1114 27011 1116
rect 26715 1062 26761 1114
rect 26761 1062 26771 1114
rect 26795 1062 26825 1114
rect 26825 1062 26837 1114
rect 26837 1062 26851 1114
rect 26875 1062 26889 1114
rect 26889 1062 26901 1114
rect 26901 1062 26931 1114
rect 26955 1062 26965 1114
rect 26965 1062 27011 1114
rect 26715 1060 26771 1062
rect 26795 1060 26851 1062
rect 26875 1060 26931 1062
rect 26955 1060 27011 1062
<< metal3 >>
rect 11247 48448 11567 48449
rect 11247 48384 11255 48448
rect 11319 48384 11335 48448
rect 11399 48384 11415 48448
rect 11479 48384 11495 48448
rect 11559 48384 11567 48448
rect 11247 48383 11567 48384
rect 21551 48448 21871 48449
rect 21551 48384 21559 48448
rect 21623 48384 21639 48448
rect 21703 48384 21719 48448
rect 21783 48384 21799 48448
rect 21863 48384 21871 48448
rect 21551 48383 21871 48384
rect 6096 47904 6416 47905
rect 6096 47840 6104 47904
rect 6168 47840 6184 47904
rect 6248 47840 6264 47904
rect 6328 47840 6344 47904
rect 6408 47840 6416 47904
rect 6096 47839 6416 47840
rect 16399 47904 16719 47905
rect 16399 47840 16407 47904
rect 16471 47840 16487 47904
rect 16551 47840 16567 47904
rect 16631 47840 16647 47904
rect 16711 47840 16719 47904
rect 16399 47839 16719 47840
rect 26703 47904 27023 47905
rect 26703 47840 26711 47904
rect 26775 47840 26791 47904
rect 26855 47840 26871 47904
rect 26935 47840 26951 47904
rect 27015 47840 27023 47904
rect 26703 47839 27023 47840
rect 11247 47360 11567 47361
rect 11247 47296 11255 47360
rect 11319 47296 11335 47360
rect 11399 47296 11415 47360
rect 11479 47296 11495 47360
rect 11559 47296 11567 47360
rect 11247 47295 11567 47296
rect 21551 47360 21871 47361
rect 21551 47296 21559 47360
rect 21623 47296 21639 47360
rect 21703 47296 21719 47360
rect 21783 47296 21799 47360
rect 21863 47296 21871 47360
rect 21551 47295 21871 47296
rect 6096 46816 6416 46817
rect 6096 46752 6104 46816
rect 6168 46752 6184 46816
rect 6248 46752 6264 46816
rect 6328 46752 6344 46816
rect 6408 46752 6416 46816
rect 6096 46751 6416 46752
rect 16399 46816 16719 46817
rect 16399 46752 16407 46816
rect 16471 46752 16487 46816
rect 16551 46752 16567 46816
rect 16631 46752 16647 46816
rect 16711 46752 16719 46816
rect 16399 46751 16719 46752
rect 26703 46816 27023 46817
rect 26703 46752 26711 46816
rect 26775 46752 26791 46816
rect 26855 46752 26871 46816
rect 26935 46752 26951 46816
rect 27015 46752 27023 46816
rect 26703 46751 27023 46752
rect 11247 46272 11567 46273
rect 11247 46208 11255 46272
rect 11319 46208 11335 46272
rect 11399 46208 11415 46272
rect 11479 46208 11495 46272
rect 11559 46208 11567 46272
rect 11247 46207 11567 46208
rect 21551 46272 21871 46273
rect 21551 46208 21559 46272
rect 21623 46208 21639 46272
rect 21703 46208 21719 46272
rect 21783 46208 21799 46272
rect 21863 46208 21871 46272
rect 21551 46207 21871 46208
rect 6096 45728 6416 45729
rect 6096 45664 6104 45728
rect 6168 45664 6184 45728
rect 6248 45664 6264 45728
rect 6328 45664 6344 45728
rect 6408 45664 6416 45728
rect 6096 45663 6416 45664
rect 16399 45728 16719 45729
rect 16399 45664 16407 45728
rect 16471 45664 16487 45728
rect 16551 45664 16567 45728
rect 16631 45664 16647 45728
rect 16711 45664 16719 45728
rect 16399 45663 16719 45664
rect 26703 45728 27023 45729
rect 26703 45664 26711 45728
rect 26775 45664 26791 45728
rect 26855 45664 26871 45728
rect 26935 45664 26951 45728
rect 27015 45664 27023 45728
rect 26703 45663 27023 45664
rect 11247 45184 11567 45185
rect 11247 45120 11255 45184
rect 11319 45120 11335 45184
rect 11399 45120 11415 45184
rect 11479 45120 11495 45184
rect 11559 45120 11567 45184
rect 11247 45119 11567 45120
rect 21551 45184 21871 45185
rect 21551 45120 21559 45184
rect 21623 45120 21639 45184
rect 21703 45120 21719 45184
rect 21783 45120 21799 45184
rect 21863 45120 21871 45184
rect 21551 45119 21871 45120
rect 6096 44640 6416 44641
rect 6096 44576 6104 44640
rect 6168 44576 6184 44640
rect 6248 44576 6264 44640
rect 6328 44576 6344 44640
rect 6408 44576 6416 44640
rect 6096 44575 6416 44576
rect 16399 44640 16719 44641
rect 16399 44576 16407 44640
rect 16471 44576 16487 44640
rect 16551 44576 16567 44640
rect 16631 44576 16647 44640
rect 16711 44576 16719 44640
rect 16399 44575 16719 44576
rect 26703 44640 27023 44641
rect 26703 44576 26711 44640
rect 26775 44576 26791 44640
rect 26855 44576 26871 44640
rect 26935 44576 26951 44640
rect 27015 44576 27023 44640
rect 26703 44575 27023 44576
rect 11247 44096 11567 44097
rect 11247 44032 11255 44096
rect 11319 44032 11335 44096
rect 11399 44032 11415 44096
rect 11479 44032 11495 44096
rect 11559 44032 11567 44096
rect 11247 44031 11567 44032
rect 21551 44096 21871 44097
rect 21551 44032 21559 44096
rect 21623 44032 21639 44096
rect 21703 44032 21719 44096
rect 21783 44032 21799 44096
rect 21863 44032 21871 44096
rect 21551 44031 21871 44032
rect 6096 43552 6416 43553
rect 6096 43488 6104 43552
rect 6168 43488 6184 43552
rect 6248 43488 6264 43552
rect 6328 43488 6344 43552
rect 6408 43488 6416 43552
rect 6096 43487 6416 43488
rect 16399 43552 16719 43553
rect 16399 43488 16407 43552
rect 16471 43488 16487 43552
rect 16551 43488 16567 43552
rect 16631 43488 16647 43552
rect 16711 43488 16719 43552
rect 16399 43487 16719 43488
rect 26703 43552 27023 43553
rect 26703 43488 26711 43552
rect 26775 43488 26791 43552
rect 26855 43488 26871 43552
rect 26935 43488 26951 43552
rect 27015 43488 27023 43552
rect 26703 43487 27023 43488
rect 11247 43008 11567 43009
rect 11247 42944 11255 43008
rect 11319 42944 11335 43008
rect 11399 42944 11415 43008
rect 11479 42944 11495 43008
rect 11559 42944 11567 43008
rect 11247 42943 11567 42944
rect 21551 43008 21871 43009
rect 21551 42944 21559 43008
rect 21623 42944 21639 43008
rect 21703 42944 21719 43008
rect 21783 42944 21799 43008
rect 21863 42944 21871 43008
rect 21551 42943 21871 42944
rect 6096 42464 6416 42465
rect 6096 42400 6104 42464
rect 6168 42400 6184 42464
rect 6248 42400 6264 42464
rect 6328 42400 6344 42464
rect 6408 42400 6416 42464
rect 6096 42399 6416 42400
rect 16399 42464 16719 42465
rect 16399 42400 16407 42464
rect 16471 42400 16487 42464
rect 16551 42400 16567 42464
rect 16631 42400 16647 42464
rect 16711 42400 16719 42464
rect 16399 42399 16719 42400
rect 26703 42464 27023 42465
rect 26703 42400 26711 42464
rect 26775 42400 26791 42464
rect 26855 42400 26871 42464
rect 26935 42400 26951 42464
rect 27015 42400 27023 42464
rect 26703 42399 27023 42400
rect 11247 41920 11567 41921
rect 11247 41856 11255 41920
rect 11319 41856 11335 41920
rect 11399 41856 11415 41920
rect 11479 41856 11495 41920
rect 11559 41856 11567 41920
rect 11247 41855 11567 41856
rect 21551 41920 21871 41921
rect 21551 41856 21559 41920
rect 21623 41856 21639 41920
rect 21703 41856 21719 41920
rect 21783 41856 21799 41920
rect 21863 41856 21871 41920
rect 21551 41855 21871 41856
rect 6096 41376 6416 41377
rect 6096 41312 6104 41376
rect 6168 41312 6184 41376
rect 6248 41312 6264 41376
rect 6328 41312 6344 41376
rect 6408 41312 6416 41376
rect 6096 41311 6416 41312
rect 16399 41376 16719 41377
rect 16399 41312 16407 41376
rect 16471 41312 16487 41376
rect 16551 41312 16567 41376
rect 16631 41312 16647 41376
rect 16711 41312 16719 41376
rect 16399 41311 16719 41312
rect 26703 41376 27023 41377
rect 26703 41312 26711 41376
rect 26775 41312 26791 41376
rect 26855 41312 26871 41376
rect 26935 41312 26951 41376
rect 27015 41312 27023 41376
rect 26703 41311 27023 41312
rect 11247 40832 11567 40833
rect 11247 40768 11255 40832
rect 11319 40768 11335 40832
rect 11399 40768 11415 40832
rect 11479 40768 11495 40832
rect 11559 40768 11567 40832
rect 11247 40767 11567 40768
rect 21551 40832 21871 40833
rect 21551 40768 21559 40832
rect 21623 40768 21639 40832
rect 21703 40768 21719 40832
rect 21783 40768 21799 40832
rect 21863 40768 21871 40832
rect 21551 40767 21871 40768
rect 6096 40288 6416 40289
rect 6096 40224 6104 40288
rect 6168 40224 6184 40288
rect 6248 40224 6264 40288
rect 6328 40224 6344 40288
rect 6408 40224 6416 40288
rect 6096 40223 6416 40224
rect 16399 40288 16719 40289
rect 16399 40224 16407 40288
rect 16471 40224 16487 40288
rect 16551 40224 16567 40288
rect 16631 40224 16647 40288
rect 16711 40224 16719 40288
rect 16399 40223 16719 40224
rect 26703 40288 27023 40289
rect 26703 40224 26711 40288
rect 26775 40224 26791 40288
rect 26855 40224 26871 40288
rect 26935 40224 26951 40288
rect 27015 40224 27023 40288
rect 26703 40223 27023 40224
rect 11247 39744 11567 39745
rect 11247 39680 11255 39744
rect 11319 39680 11335 39744
rect 11399 39680 11415 39744
rect 11479 39680 11495 39744
rect 11559 39680 11567 39744
rect 11247 39679 11567 39680
rect 21551 39744 21871 39745
rect 21551 39680 21559 39744
rect 21623 39680 21639 39744
rect 21703 39680 21719 39744
rect 21783 39680 21799 39744
rect 21863 39680 21871 39744
rect 21551 39679 21871 39680
rect 6096 39200 6416 39201
rect 6096 39136 6104 39200
rect 6168 39136 6184 39200
rect 6248 39136 6264 39200
rect 6328 39136 6344 39200
rect 6408 39136 6416 39200
rect 6096 39135 6416 39136
rect 16399 39200 16719 39201
rect 16399 39136 16407 39200
rect 16471 39136 16487 39200
rect 16551 39136 16567 39200
rect 16631 39136 16647 39200
rect 16711 39136 16719 39200
rect 16399 39135 16719 39136
rect 26703 39200 27023 39201
rect 26703 39136 26711 39200
rect 26775 39136 26791 39200
rect 26855 39136 26871 39200
rect 26935 39136 26951 39200
rect 27015 39136 27023 39200
rect 26703 39135 27023 39136
rect 11247 38656 11567 38657
rect 11247 38592 11255 38656
rect 11319 38592 11335 38656
rect 11399 38592 11415 38656
rect 11479 38592 11495 38656
rect 11559 38592 11567 38656
rect 11247 38591 11567 38592
rect 21551 38656 21871 38657
rect 21551 38592 21559 38656
rect 21623 38592 21639 38656
rect 21703 38592 21719 38656
rect 21783 38592 21799 38656
rect 21863 38592 21871 38656
rect 21551 38591 21871 38592
rect 6096 38112 6416 38113
rect 6096 38048 6104 38112
rect 6168 38048 6184 38112
rect 6248 38048 6264 38112
rect 6328 38048 6344 38112
rect 6408 38048 6416 38112
rect 6096 38047 6416 38048
rect 16399 38112 16719 38113
rect 16399 38048 16407 38112
rect 16471 38048 16487 38112
rect 16551 38048 16567 38112
rect 16631 38048 16647 38112
rect 16711 38048 16719 38112
rect 16399 38047 16719 38048
rect 26703 38112 27023 38113
rect 26703 38048 26711 38112
rect 26775 38048 26791 38112
rect 26855 38048 26871 38112
rect 26935 38048 26951 38112
rect 27015 38048 27023 38112
rect 26703 38047 27023 38048
rect 11247 37568 11567 37569
rect 11247 37504 11255 37568
rect 11319 37504 11335 37568
rect 11399 37504 11415 37568
rect 11479 37504 11495 37568
rect 11559 37504 11567 37568
rect 11247 37503 11567 37504
rect 21551 37568 21871 37569
rect 21551 37504 21559 37568
rect 21623 37504 21639 37568
rect 21703 37504 21719 37568
rect 21783 37504 21799 37568
rect 21863 37504 21871 37568
rect 21551 37503 21871 37504
rect 6096 37024 6416 37025
rect 6096 36960 6104 37024
rect 6168 36960 6184 37024
rect 6248 36960 6264 37024
rect 6328 36960 6344 37024
rect 6408 36960 6416 37024
rect 6096 36959 6416 36960
rect 16399 37024 16719 37025
rect 16399 36960 16407 37024
rect 16471 36960 16487 37024
rect 16551 36960 16567 37024
rect 16631 36960 16647 37024
rect 16711 36960 16719 37024
rect 16399 36959 16719 36960
rect 26703 37024 27023 37025
rect 26703 36960 26711 37024
rect 26775 36960 26791 37024
rect 26855 36960 26871 37024
rect 26935 36960 26951 37024
rect 27015 36960 27023 37024
rect 26703 36959 27023 36960
rect 11247 36480 11567 36481
rect 11247 36416 11255 36480
rect 11319 36416 11335 36480
rect 11399 36416 11415 36480
rect 11479 36416 11495 36480
rect 11559 36416 11567 36480
rect 11247 36415 11567 36416
rect 21551 36480 21871 36481
rect 21551 36416 21559 36480
rect 21623 36416 21639 36480
rect 21703 36416 21719 36480
rect 21783 36416 21799 36480
rect 21863 36416 21871 36480
rect 21551 36415 21871 36416
rect 6096 35936 6416 35937
rect 6096 35872 6104 35936
rect 6168 35872 6184 35936
rect 6248 35872 6264 35936
rect 6328 35872 6344 35936
rect 6408 35872 6416 35936
rect 6096 35871 6416 35872
rect 16399 35936 16719 35937
rect 16399 35872 16407 35936
rect 16471 35872 16487 35936
rect 16551 35872 16567 35936
rect 16631 35872 16647 35936
rect 16711 35872 16719 35936
rect 16399 35871 16719 35872
rect 26703 35936 27023 35937
rect 26703 35872 26711 35936
rect 26775 35872 26791 35936
rect 26855 35872 26871 35936
rect 26935 35872 26951 35936
rect 27015 35872 27023 35936
rect 26703 35871 27023 35872
rect 11247 35392 11567 35393
rect 11247 35328 11255 35392
rect 11319 35328 11335 35392
rect 11399 35328 11415 35392
rect 11479 35328 11495 35392
rect 11559 35328 11567 35392
rect 11247 35327 11567 35328
rect 21551 35392 21871 35393
rect 21551 35328 21559 35392
rect 21623 35328 21639 35392
rect 21703 35328 21719 35392
rect 21783 35328 21799 35392
rect 21863 35328 21871 35392
rect 21551 35327 21871 35328
rect 6096 34848 6416 34849
rect 6096 34784 6104 34848
rect 6168 34784 6184 34848
rect 6248 34784 6264 34848
rect 6328 34784 6344 34848
rect 6408 34784 6416 34848
rect 6096 34783 6416 34784
rect 16399 34848 16719 34849
rect 16399 34784 16407 34848
rect 16471 34784 16487 34848
rect 16551 34784 16567 34848
rect 16631 34784 16647 34848
rect 16711 34784 16719 34848
rect 16399 34783 16719 34784
rect 26703 34848 27023 34849
rect 26703 34784 26711 34848
rect 26775 34784 26791 34848
rect 26855 34784 26871 34848
rect 26935 34784 26951 34848
rect 27015 34784 27023 34848
rect 26703 34783 27023 34784
rect 11247 34304 11567 34305
rect 11247 34240 11255 34304
rect 11319 34240 11335 34304
rect 11399 34240 11415 34304
rect 11479 34240 11495 34304
rect 11559 34240 11567 34304
rect 11247 34239 11567 34240
rect 21551 34304 21871 34305
rect 21551 34240 21559 34304
rect 21623 34240 21639 34304
rect 21703 34240 21719 34304
rect 21783 34240 21799 34304
rect 21863 34240 21871 34304
rect 21551 34239 21871 34240
rect 6096 33760 6416 33761
rect 6096 33696 6104 33760
rect 6168 33696 6184 33760
rect 6248 33696 6264 33760
rect 6328 33696 6344 33760
rect 6408 33696 6416 33760
rect 6096 33695 6416 33696
rect 16399 33760 16719 33761
rect 16399 33696 16407 33760
rect 16471 33696 16487 33760
rect 16551 33696 16567 33760
rect 16631 33696 16647 33760
rect 16711 33696 16719 33760
rect 16399 33695 16719 33696
rect 26703 33760 27023 33761
rect 26703 33696 26711 33760
rect 26775 33696 26791 33760
rect 26855 33696 26871 33760
rect 26935 33696 26951 33760
rect 27015 33696 27023 33760
rect 26703 33695 27023 33696
rect 11247 33216 11567 33217
rect 11247 33152 11255 33216
rect 11319 33152 11335 33216
rect 11399 33152 11415 33216
rect 11479 33152 11495 33216
rect 11559 33152 11567 33216
rect 11247 33151 11567 33152
rect 21551 33216 21871 33217
rect 21551 33152 21559 33216
rect 21623 33152 21639 33216
rect 21703 33152 21719 33216
rect 21783 33152 21799 33216
rect 21863 33152 21871 33216
rect 21551 33151 21871 33152
rect 6096 32672 6416 32673
rect 6096 32608 6104 32672
rect 6168 32608 6184 32672
rect 6248 32608 6264 32672
rect 6328 32608 6344 32672
rect 6408 32608 6416 32672
rect 6096 32607 6416 32608
rect 16399 32672 16719 32673
rect 16399 32608 16407 32672
rect 16471 32608 16487 32672
rect 16551 32608 16567 32672
rect 16631 32608 16647 32672
rect 16711 32608 16719 32672
rect 16399 32607 16719 32608
rect 26703 32672 27023 32673
rect 26703 32608 26711 32672
rect 26775 32608 26791 32672
rect 26855 32608 26871 32672
rect 26935 32608 26951 32672
rect 27015 32608 27023 32672
rect 26703 32607 27023 32608
rect 11247 32128 11567 32129
rect 11247 32064 11255 32128
rect 11319 32064 11335 32128
rect 11399 32064 11415 32128
rect 11479 32064 11495 32128
rect 11559 32064 11567 32128
rect 11247 32063 11567 32064
rect 21551 32128 21871 32129
rect 21551 32064 21559 32128
rect 21623 32064 21639 32128
rect 21703 32064 21719 32128
rect 21783 32064 21799 32128
rect 21863 32064 21871 32128
rect 21551 32063 21871 32064
rect 6096 31584 6416 31585
rect 6096 31520 6104 31584
rect 6168 31520 6184 31584
rect 6248 31520 6264 31584
rect 6328 31520 6344 31584
rect 6408 31520 6416 31584
rect 6096 31519 6416 31520
rect 16399 31584 16719 31585
rect 16399 31520 16407 31584
rect 16471 31520 16487 31584
rect 16551 31520 16567 31584
rect 16631 31520 16647 31584
rect 16711 31520 16719 31584
rect 16399 31519 16719 31520
rect 26703 31584 27023 31585
rect 26703 31520 26711 31584
rect 26775 31520 26791 31584
rect 26855 31520 26871 31584
rect 26935 31520 26951 31584
rect 27015 31520 27023 31584
rect 26703 31519 27023 31520
rect 11247 31040 11567 31041
rect 11247 30976 11255 31040
rect 11319 30976 11335 31040
rect 11399 30976 11415 31040
rect 11479 30976 11495 31040
rect 11559 30976 11567 31040
rect 11247 30975 11567 30976
rect 21551 31040 21871 31041
rect 21551 30976 21559 31040
rect 21623 30976 21639 31040
rect 21703 30976 21719 31040
rect 21783 30976 21799 31040
rect 21863 30976 21871 31040
rect 21551 30975 21871 30976
rect 6096 30496 6416 30497
rect 6096 30432 6104 30496
rect 6168 30432 6184 30496
rect 6248 30432 6264 30496
rect 6328 30432 6344 30496
rect 6408 30432 6416 30496
rect 6096 30431 6416 30432
rect 16399 30496 16719 30497
rect 16399 30432 16407 30496
rect 16471 30432 16487 30496
rect 16551 30432 16567 30496
rect 16631 30432 16647 30496
rect 16711 30432 16719 30496
rect 16399 30431 16719 30432
rect 26703 30496 27023 30497
rect 26703 30432 26711 30496
rect 26775 30432 26791 30496
rect 26855 30432 26871 30496
rect 26935 30432 26951 30496
rect 27015 30432 27023 30496
rect 26703 30431 27023 30432
rect 11247 29952 11567 29953
rect 11247 29888 11255 29952
rect 11319 29888 11335 29952
rect 11399 29888 11415 29952
rect 11479 29888 11495 29952
rect 11559 29888 11567 29952
rect 11247 29887 11567 29888
rect 21551 29952 21871 29953
rect 21551 29888 21559 29952
rect 21623 29888 21639 29952
rect 21703 29888 21719 29952
rect 21783 29888 21799 29952
rect 21863 29888 21871 29952
rect 21551 29887 21871 29888
rect 6096 29408 6416 29409
rect 6096 29344 6104 29408
rect 6168 29344 6184 29408
rect 6248 29344 6264 29408
rect 6328 29344 6344 29408
rect 6408 29344 6416 29408
rect 6096 29343 6416 29344
rect 16399 29408 16719 29409
rect 16399 29344 16407 29408
rect 16471 29344 16487 29408
rect 16551 29344 16567 29408
rect 16631 29344 16647 29408
rect 16711 29344 16719 29408
rect 16399 29343 16719 29344
rect 26703 29408 27023 29409
rect 26703 29344 26711 29408
rect 26775 29344 26791 29408
rect 26855 29344 26871 29408
rect 26935 29344 26951 29408
rect 27015 29344 27023 29408
rect 26703 29343 27023 29344
rect 11247 28864 11567 28865
rect 11247 28800 11255 28864
rect 11319 28800 11335 28864
rect 11399 28800 11415 28864
rect 11479 28800 11495 28864
rect 11559 28800 11567 28864
rect 11247 28799 11567 28800
rect 21551 28864 21871 28865
rect 21551 28800 21559 28864
rect 21623 28800 21639 28864
rect 21703 28800 21719 28864
rect 21783 28800 21799 28864
rect 21863 28800 21871 28864
rect 21551 28799 21871 28800
rect 6096 28320 6416 28321
rect 6096 28256 6104 28320
rect 6168 28256 6184 28320
rect 6248 28256 6264 28320
rect 6328 28256 6344 28320
rect 6408 28256 6416 28320
rect 6096 28255 6416 28256
rect 16399 28320 16719 28321
rect 16399 28256 16407 28320
rect 16471 28256 16487 28320
rect 16551 28256 16567 28320
rect 16631 28256 16647 28320
rect 16711 28256 16719 28320
rect 16399 28255 16719 28256
rect 26703 28320 27023 28321
rect 26703 28256 26711 28320
rect 26775 28256 26791 28320
rect 26855 28256 26871 28320
rect 26935 28256 26951 28320
rect 27015 28256 27023 28320
rect 26703 28255 27023 28256
rect 11247 27776 11567 27777
rect 11247 27712 11255 27776
rect 11319 27712 11335 27776
rect 11399 27712 11415 27776
rect 11479 27712 11495 27776
rect 11559 27712 11567 27776
rect 11247 27711 11567 27712
rect 21551 27776 21871 27777
rect 21551 27712 21559 27776
rect 21623 27712 21639 27776
rect 21703 27712 21719 27776
rect 21783 27712 21799 27776
rect 21863 27712 21871 27776
rect 21551 27711 21871 27712
rect 6096 27232 6416 27233
rect 6096 27168 6104 27232
rect 6168 27168 6184 27232
rect 6248 27168 6264 27232
rect 6328 27168 6344 27232
rect 6408 27168 6416 27232
rect 6096 27167 6416 27168
rect 16399 27232 16719 27233
rect 16399 27168 16407 27232
rect 16471 27168 16487 27232
rect 16551 27168 16567 27232
rect 16631 27168 16647 27232
rect 16711 27168 16719 27232
rect 16399 27167 16719 27168
rect 26703 27232 27023 27233
rect 26703 27168 26711 27232
rect 26775 27168 26791 27232
rect 26855 27168 26871 27232
rect 26935 27168 26951 27232
rect 27015 27168 27023 27232
rect 26703 27167 27023 27168
rect 11247 26688 11567 26689
rect 11247 26624 11255 26688
rect 11319 26624 11335 26688
rect 11399 26624 11415 26688
rect 11479 26624 11495 26688
rect 11559 26624 11567 26688
rect 11247 26623 11567 26624
rect 21551 26688 21871 26689
rect 21551 26624 21559 26688
rect 21623 26624 21639 26688
rect 21703 26624 21719 26688
rect 21783 26624 21799 26688
rect 21863 26624 21871 26688
rect 21551 26623 21871 26624
rect 6096 26144 6416 26145
rect 6096 26080 6104 26144
rect 6168 26080 6184 26144
rect 6248 26080 6264 26144
rect 6328 26080 6344 26144
rect 6408 26080 6416 26144
rect 6096 26079 6416 26080
rect 16399 26144 16719 26145
rect 16399 26080 16407 26144
rect 16471 26080 16487 26144
rect 16551 26080 16567 26144
rect 16631 26080 16647 26144
rect 16711 26080 16719 26144
rect 16399 26079 16719 26080
rect 26703 26144 27023 26145
rect 26703 26080 26711 26144
rect 26775 26080 26791 26144
rect 26855 26080 26871 26144
rect 26935 26080 26951 26144
rect 27015 26080 27023 26144
rect 26703 26079 27023 26080
rect 11247 25600 11567 25601
rect 11247 25536 11255 25600
rect 11319 25536 11335 25600
rect 11399 25536 11415 25600
rect 11479 25536 11495 25600
rect 11559 25536 11567 25600
rect 11247 25535 11567 25536
rect 21551 25600 21871 25601
rect 21551 25536 21559 25600
rect 21623 25536 21639 25600
rect 21703 25536 21719 25600
rect 21783 25536 21799 25600
rect 21863 25536 21871 25600
rect 21551 25535 21871 25536
rect 6096 25056 6416 25057
rect 6096 24992 6104 25056
rect 6168 24992 6184 25056
rect 6248 24992 6264 25056
rect 6328 24992 6344 25056
rect 6408 24992 6416 25056
rect 6096 24991 6416 24992
rect 16399 25056 16719 25057
rect 16399 24992 16407 25056
rect 16471 24992 16487 25056
rect 16551 24992 16567 25056
rect 16631 24992 16647 25056
rect 16711 24992 16719 25056
rect 16399 24991 16719 24992
rect 26703 25056 27023 25057
rect 26703 24992 26711 25056
rect 26775 24992 26791 25056
rect 26855 24992 26871 25056
rect 26935 24992 26951 25056
rect 27015 24992 27023 25056
rect 26703 24991 27023 24992
rect 11247 24512 11567 24513
rect 11247 24448 11255 24512
rect 11319 24448 11335 24512
rect 11399 24448 11415 24512
rect 11479 24448 11495 24512
rect 11559 24448 11567 24512
rect 11247 24447 11567 24448
rect 21551 24512 21871 24513
rect 21551 24448 21559 24512
rect 21623 24448 21639 24512
rect 21703 24448 21719 24512
rect 21783 24448 21799 24512
rect 21863 24448 21871 24512
rect 21551 24447 21871 24448
rect 6096 23968 6416 23969
rect 6096 23904 6104 23968
rect 6168 23904 6184 23968
rect 6248 23904 6264 23968
rect 6328 23904 6344 23968
rect 6408 23904 6416 23968
rect 6096 23903 6416 23904
rect 16399 23968 16719 23969
rect 16399 23904 16407 23968
rect 16471 23904 16487 23968
rect 16551 23904 16567 23968
rect 16631 23904 16647 23968
rect 16711 23904 16719 23968
rect 16399 23903 16719 23904
rect 26703 23968 27023 23969
rect 26703 23904 26711 23968
rect 26775 23904 26791 23968
rect 26855 23904 26871 23968
rect 26935 23904 26951 23968
rect 27015 23904 27023 23968
rect 26703 23903 27023 23904
rect 11247 23424 11567 23425
rect 11247 23360 11255 23424
rect 11319 23360 11335 23424
rect 11399 23360 11415 23424
rect 11479 23360 11495 23424
rect 11559 23360 11567 23424
rect 11247 23359 11567 23360
rect 21551 23424 21871 23425
rect 21551 23360 21559 23424
rect 21623 23360 21639 23424
rect 21703 23360 21719 23424
rect 21783 23360 21799 23424
rect 21863 23360 21871 23424
rect 21551 23359 21871 23360
rect 6096 22880 6416 22881
rect 6096 22816 6104 22880
rect 6168 22816 6184 22880
rect 6248 22816 6264 22880
rect 6328 22816 6344 22880
rect 6408 22816 6416 22880
rect 6096 22815 6416 22816
rect 16399 22880 16719 22881
rect 16399 22816 16407 22880
rect 16471 22816 16487 22880
rect 16551 22816 16567 22880
rect 16631 22816 16647 22880
rect 16711 22816 16719 22880
rect 16399 22815 16719 22816
rect 26703 22880 27023 22881
rect 26703 22816 26711 22880
rect 26775 22816 26791 22880
rect 26855 22816 26871 22880
rect 26935 22816 26951 22880
rect 27015 22816 27023 22880
rect 26703 22815 27023 22816
rect 11247 22336 11567 22337
rect 11247 22272 11255 22336
rect 11319 22272 11335 22336
rect 11399 22272 11415 22336
rect 11479 22272 11495 22336
rect 11559 22272 11567 22336
rect 11247 22271 11567 22272
rect 21551 22336 21871 22337
rect 21551 22272 21559 22336
rect 21623 22272 21639 22336
rect 21703 22272 21719 22336
rect 21783 22272 21799 22336
rect 21863 22272 21871 22336
rect 21551 22271 21871 22272
rect 6096 21792 6416 21793
rect 6096 21728 6104 21792
rect 6168 21728 6184 21792
rect 6248 21728 6264 21792
rect 6328 21728 6344 21792
rect 6408 21728 6416 21792
rect 6096 21727 6416 21728
rect 16399 21792 16719 21793
rect 16399 21728 16407 21792
rect 16471 21728 16487 21792
rect 16551 21728 16567 21792
rect 16631 21728 16647 21792
rect 16711 21728 16719 21792
rect 16399 21727 16719 21728
rect 26703 21792 27023 21793
rect 26703 21728 26711 21792
rect 26775 21728 26791 21792
rect 26855 21728 26871 21792
rect 26935 21728 26951 21792
rect 27015 21728 27023 21792
rect 26703 21727 27023 21728
rect 11247 21248 11567 21249
rect 11247 21184 11255 21248
rect 11319 21184 11335 21248
rect 11399 21184 11415 21248
rect 11479 21184 11495 21248
rect 11559 21184 11567 21248
rect 11247 21183 11567 21184
rect 21551 21248 21871 21249
rect 21551 21184 21559 21248
rect 21623 21184 21639 21248
rect 21703 21184 21719 21248
rect 21783 21184 21799 21248
rect 21863 21184 21871 21248
rect 21551 21183 21871 21184
rect 6096 20704 6416 20705
rect 6096 20640 6104 20704
rect 6168 20640 6184 20704
rect 6248 20640 6264 20704
rect 6328 20640 6344 20704
rect 6408 20640 6416 20704
rect 6096 20639 6416 20640
rect 16399 20704 16719 20705
rect 16399 20640 16407 20704
rect 16471 20640 16487 20704
rect 16551 20640 16567 20704
rect 16631 20640 16647 20704
rect 16711 20640 16719 20704
rect 16399 20639 16719 20640
rect 26703 20704 27023 20705
rect 26703 20640 26711 20704
rect 26775 20640 26791 20704
rect 26855 20640 26871 20704
rect 26935 20640 26951 20704
rect 27015 20640 27023 20704
rect 26703 20639 27023 20640
rect 11247 20160 11567 20161
rect 11247 20096 11255 20160
rect 11319 20096 11335 20160
rect 11399 20096 11415 20160
rect 11479 20096 11495 20160
rect 11559 20096 11567 20160
rect 11247 20095 11567 20096
rect 21551 20160 21871 20161
rect 21551 20096 21559 20160
rect 21623 20096 21639 20160
rect 21703 20096 21719 20160
rect 21783 20096 21799 20160
rect 21863 20096 21871 20160
rect 21551 20095 21871 20096
rect 6096 19616 6416 19617
rect 6096 19552 6104 19616
rect 6168 19552 6184 19616
rect 6248 19552 6264 19616
rect 6328 19552 6344 19616
rect 6408 19552 6416 19616
rect 6096 19551 6416 19552
rect 16399 19616 16719 19617
rect 16399 19552 16407 19616
rect 16471 19552 16487 19616
rect 16551 19552 16567 19616
rect 16631 19552 16647 19616
rect 16711 19552 16719 19616
rect 16399 19551 16719 19552
rect 26703 19616 27023 19617
rect 26703 19552 26711 19616
rect 26775 19552 26791 19616
rect 26855 19552 26871 19616
rect 26935 19552 26951 19616
rect 27015 19552 27023 19616
rect 26703 19551 27023 19552
rect 11247 19072 11567 19073
rect 11247 19008 11255 19072
rect 11319 19008 11335 19072
rect 11399 19008 11415 19072
rect 11479 19008 11495 19072
rect 11559 19008 11567 19072
rect 11247 19007 11567 19008
rect 21551 19072 21871 19073
rect 21551 19008 21559 19072
rect 21623 19008 21639 19072
rect 21703 19008 21719 19072
rect 21783 19008 21799 19072
rect 21863 19008 21871 19072
rect 21551 19007 21871 19008
rect 6096 18528 6416 18529
rect 6096 18464 6104 18528
rect 6168 18464 6184 18528
rect 6248 18464 6264 18528
rect 6328 18464 6344 18528
rect 6408 18464 6416 18528
rect 6096 18463 6416 18464
rect 16399 18528 16719 18529
rect 16399 18464 16407 18528
rect 16471 18464 16487 18528
rect 16551 18464 16567 18528
rect 16631 18464 16647 18528
rect 16711 18464 16719 18528
rect 16399 18463 16719 18464
rect 26703 18528 27023 18529
rect 26703 18464 26711 18528
rect 26775 18464 26791 18528
rect 26855 18464 26871 18528
rect 26935 18464 26951 18528
rect 27015 18464 27023 18528
rect 26703 18463 27023 18464
rect 11247 17984 11567 17985
rect 11247 17920 11255 17984
rect 11319 17920 11335 17984
rect 11399 17920 11415 17984
rect 11479 17920 11495 17984
rect 11559 17920 11567 17984
rect 11247 17919 11567 17920
rect 21551 17984 21871 17985
rect 21551 17920 21559 17984
rect 21623 17920 21639 17984
rect 21703 17920 21719 17984
rect 21783 17920 21799 17984
rect 21863 17920 21871 17984
rect 21551 17919 21871 17920
rect 6096 17440 6416 17441
rect 6096 17376 6104 17440
rect 6168 17376 6184 17440
rect 6248 17376 6264 17440
rect 6328 17376 6344 17440
rect 6408 17376 6416 17440
rect 6096 17375 6416 17376
rect 16399 17440 16719 17441
rect 16399 17376 16407 17440
rect 16471 17376 16487 17440
rect 16551 17376 16567 17440
rect 16631 17376 16647 17440
rect 16711 17376 16719 17440
rect 16399 17375 16719 17376
rect 26703 17440 27023 17441
rect 26703 17376 26711 17440
rect 26775 17376 26791 17440
rect 26855 17376 26871 17440
rect 26935 17376 26951 17440
rect 27015 17376 27023 17440
rect 26703 17375 27023 17376
rect 11247 16896 11567 16897
rect 11247 16832 11255 16896
rect 11319 16832 11335 16896
rect 11399 16832 11415 16896
rect 11479 16832 11495 16896
rect 11559 16832 11567 16896
rect 11247 16831 11567 16832
rect 21551 16896 21871 16897
rect 21551 16832 21559 16896
rect 21623 16832 21639 16896
rect 21703 16832 21719 16896
rect 21783 16832 21799 16896
rect 21863 16832 21871 16896
rect 21551 16831 21871 16832
rect 6096 16352 6416 16353
rect 6096 16288 6104 16352
rect 6168 16288 6184 16352
rect 6248 16288 6264 16352
rect 6328 16288 6344 16352
rect 6408 16288 6416 16352
rect 6096 16287 6416 16288
rect 16399 16352 16719 16353
rect 16399 16288 16407 16352
rect 16471 16288 16487 16352
rect 16551 16288 16567 16352
rect 16631 16288 16647 16352
rect 16711 16288 16719 16352
rect 16399 16287 16719 16288
rect 26703 16352 27023 16353
rect 26703 16288 26711 16352
rect 26775 16288 26791 16352
rect 26855 16288 26871 16352
rect 26935 16288 26951 16352
rect 27015 16288 27023 16352
rect 26703 16287 27023 16288
rect 11247 15808 11567 15809
rect 11247 15744 11255 15808
rect 11319 15744 11335 15808
rect 11399 15744 11415 15808
rect 11479 15744 11495 15808
rect 11559 15744 11567 15808
rect 11247 15743 11567 15744
rect 21551 15808 21871 15809
rect 21551 15744 21559 15808
rect 21623 15744 21639 15808
rect 21703 15744 21719 15808
rect 21783 15744 21799 15808
rect 21863 15744 21871 15808
rect 21551 15743 21871 15744
rect 6096 15264 6416 15265
rect 6096 15200 6104 15264
rect 6168 15200 6184 15264
rect 6248 15200 6264 15264
rect 6328 15200 6344 15264
rect 6408 15200 6416 15264
rect 6096 15199 6416 15200
rect 16399 15264 16719 15265
rect 16399 15200 16407 15264
rect 16471 15200 16487 15264
rect 16551 15200 16567 15264
rect 16631 15200 16647 15264
rect 16711 15200 16719 15264
rect 16399 15199 16719 15200
rect 26703 15264 27023 15265
rect 26703 15200 26711 15264
rect 26775 15200 26791 15264
rect 26855 15200 26871 15264
rect 26935 15200 26951 15264
rect 27015 15200 27023 15264
rect 26703 15199 27023 15200
rect 11247 14720 11567 14721
rect 11247 14656 11255 14720
rect 11319 14656 11335 14720
rect 11399 14656 11415 14720
rect 11479 14656 11495 14720
rect 11559 14656 11567 14720
rect 11247 14655 11567 14656
rect 21551 14720 21871 14721
rect 21551 14656 21559 14720
rect 21623 14656 21639 14720
rect 21703 14656 21719 14720
rect 21783 14656 21799 14720
rect 21863 14656 21871 14720
rect 21551 14655 21871 14656
rect 6096 14176 6416 14177
rect 6096 14112 6104 14176
rect 6168 14112 6184 14176
rect 6248 14112 6264 14176
rect 6328 14112 6344 14176
rect 6408 14112 6416 14176
rect 6096 14111 6416 14112
rect 16399 14176 16719 14177
rect 16399 14112 16407 14176
rect 16471 14112 16487 14176
rect 16551 14112 16567 14176
rect 16631 14112 16647 14176
rect 16711 14112 16719 14176
rect 16399 14111 16719 14112
rect 26703 14176 27023 14177
rect 26703 14112 26711 14176
rect 26775 14112 26791 14176
rect 26855 14112 26871 14176
rect 26935 14112 26951 14176
rect 27015 14112 27023 14176
rect 26703 14111 27023 14112
rect 11247 13632 11567 13633
rect 11247 13568 11255 13632
rect 11319 13568 11335 13632
rect 11399 13568 11415 13632
rect 11479 13568 11495 13632
rect 11559 13568 11567 13632
rect 11247 13567 11567 13568
rect 21551 13632 21871 13633
rect 21551 13568 21559 13632
rect 21623 13568 21639 13632
rect 21703 13568 21719 13632
rect 21783 13568 21799 13632
rect 21863 13568 21871 13632
rect 21551 13567 21871 13568
rect 6096 13088 6416 13089
rect 6096 13024 6104 13088
rect 6168 13024 6184 13088
rect 6248 13024 6264 13088
rect 6328 13024 6344 13088
rect 6408 13024 6416 13088
rect 6096 13023 6416 13024
rect 16399 13088 16719 13089
rect 16399 13024 16407 13088
rect 16471 13024 16487 13088
rect 16551 13024 16567 13088
rect 16631 13024 16647 13088
rect 16711 13024 16719 13088
rect 16399 13023 16719 13024
rect 26703 13088 27023 13089
rect 26703 13024 26711 13088
rect 26775 13024 26791 13088
rect 26855 13024 26871 13088
rect 26935 13024 26951 13088
rect 27015 13024 27023 13088
rect 26703 13023 27023 13024
rect 11247 12544 11567 12545
rect 11247 12480 11255 12544
rect 11319 12480 11335 12544
rect 11399 12480 11415 12544
rect 11479 12480 11495 12544
rect 11559 12480 11567 12544
rect 11247 12479 11567 12480
rect 21551 12544 21871 12545
rect 21551 12480 21559 12544
rect 21623 12480 21639 12544
rect 21703 12480 21719 12544
rect 21783 12480 21799 12544
rect 21863 12480 21871 12544
rect 21551 12479 21871 12480
rect 6096 12000 6416 12001
rect 6096 11936 6104 12000
rect 6168 11936 6184 12000
rect 6248 11936 6264 12000
rect 6328 11936 6344 12000
rect 6408 11936 6416 12000
rect 6096 11935 6416 11936
rect 16399 12000 16719 12001
rect 16399 11936 16407 12000
rect 16471 11936 16487 12000
rect 16551 11936 16567 12000
rect 16631 11936 16647 12000
rect 16711 11936 16719 12000
rect 16399 11935 16719 11936
rect 26703 12000 27023 12001
rect 26703 11936 26711 12000
rect 26775 11936 26791 12000
rect 26855 11936 26871 12000
rect 26935 11936 26951 12000
rect 27015 11936 27023 12000
rect 26703 11935 27023 11936
rect 11247 11456 11567 11457
rect 11247 11392 11255 11456
rect 11319 11392 11335 11456
rect 11399 11392 11415 11456
rect 11479 11392 11495 11456
rect 11559 11392 11567 11456
rect 11247 11391 11567 11392
rect 21551 11456 21871 11457
rect 21551 11392 21559 11456
rect 21623 11392 21639 11456
rect 21703 11392 21719 11456
rect 21783 11392 21799 11456
rect 21863 11392 21871 11456
rect 21551 11391 21871 11392
rect 6096 10912 6416 10913
rect 6096 10848 6104 10912
rect 6168 10848 6184 10912
rect 6248 10848 6264 10912
rect 6328 10848 6344 10912
rect 6408 10848 6416 10912
rect 6096 10847 6416 10848
rect 16399 10912 16719 10913
rect 16399 10848 16407 10912
rect 16471 10848 16487 10912
rect 16551 10848 16567 10912
rect 16631 10848 16647 10912
rect 16711 10848 16719 10912
rect 16399 10847 16719 10848
rect 26703 10912 27023 10913
rect 26703 10848 26711 10912
rect 26775 10848 26791 10912
rect 26855 10848 26871 10912
rect 26935 10848 26951 10912
rect 27015 10848 27023 10912
rect 26703 10847 27023 10848
rect 11247 10368 11567 10369
rect 11247 10304 11255 10368
rect 11319 10304 11335 10368
rect 11399 10304 11415 10368
rect 11479 10304 11495 10368
rect 11559 10304 11567 10368
rect 11247 10303 11567 10304
rect 21551 10368 21871 10369
rect 21551 10304 21559 10368
rect 21623 10304 21639 10368
rect 21703 10304 21719 10368
rect 21783 10304 21799 10368
rect 21863 10304 21871 10368
rect 21551 10303 21871 10304
rect 6096 9824 6416 9825
rect 6096 9760 6104 9824
rect 6168 9760 6184 9824
rect 6248 9760 6264 9824
rect 6328 9760 6344 9824
rect 6408 9760 6416 9824
rect 6096 9759 6416 9760
rect 16399 9824 16719 9825
rect 16399 9760 16407 9824
rect 16471 9760 16487 9824
rect 16551 9760 16567 9824
rect 16631 9760 16647 9824
rect 16711 9760 16719 9824
rect 16399 9759 16719 9760
rect 26703 9824 27023 9825
rect 26703 9760 26711 9824
rect 26775 9760 26791 9824
rect 26855 9760 26871 9824
rect 26935 9760 26951 9824
rect 27015 9760 27023 9824
rect 26703 9759 27023 9760
rect 11247 9280 11567 9281
rect 11247 9216 11255 9280
rect 11319 9216 11335 9280
rect 11399 9216 11415 9280
rect 11479 9216 11495 9280
rect 11559 9216 11567 9280
rect 11247 9215 11567 9216
rect 21551 9280 21871 9281
rect 21551 9216 21559 9280
rect 21623 9216 21639 9280
rect 21703 9216 21719 9280
rect 21783 9216 21799 9280
rect 21863 9216 21871 9280
rect 21551 9215 21871 9216
rect 6096 8736 6416 8737
rect 6096 8672 6104 8736
rect 6168 8672 6184 8736
rect 6248 8672 6264 8736
rect 6328 8672 6344 8736
rect 6408 8672 6416 8736
rect 6096 8671 6416 8672
rect 16399 8736 16719 8737
rect 16399 8672 16407 8736
rect 16471 8672 16487 8736
rect 16551 8672 16567 8736
rect 16631 8672 16647 8736
rect 16711 8672 16719 8736
rect 16399 8671 16719 8672
rect 26703 8736 27023 8737
rect 26703 8672 26711 8736
rect 26775 8672 26791 8736
rect 26855 8672 26871 8736
rect 26935 8672 26951 8736
rect 27015 8672 27023 8736
rect 26703 8671 27023 8672
rect 11247 8192 11567 8193
rect 11247 8128 11255 8192
rect 11319 8128 11335 8192
rect 11399 8128 11415 8192
rect 11479 8128 11495 8192
rect 11559 8128 11567 8192
rect 11247 8127 11567 8128
rect 21551 8192 21871 8193
rect 21551 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21799 8192
rect 21863 8128 21871 8192
rect 21551 8127 21871 8128
rect 6096 7648 6416 7649
rect 6096 7584 6104 7648
rect 6168 7584 6184 7648
rect 6248 7584 6264 7648
rect 6328 7584 6344 7648
rect 6408 7584 6416 7648
rect 6096 7583 6416 7584
rect 16399 7648 16719 7649
rect 16399 7584 16407 7648
rect 16471 7584 16487 7648
rect 16551 7584 16567 7648
rect 16631 7584 16647 7648
rect 16711 7584 16719 7648
rect 16399 7583 16719 7584
rect 26703 7648 27023 7649
rect 26703 7584 26711 7648
rect 26775 7584 26791 7648
rect 26855 7584 26871 7648
rect 26935 7584 26951 7648
rect 27015 7584 27023 7648
rect 26703 7583 27023 7584
rect 11247 7104 11567 7105
rect 11247 7040 11255 7104
rect 11319 7040 11335 7104
rect 11399 7040 11415 7104
rect 11479 7040 11495 7104
rect 11559 7040 11567 7104
rect 11247 7039 11567 7040
rect 21551 7104 21871 7105
rect 21551 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21799 7104
rect 21863 7040 21871 7104
rect 21551 7039 21871 7040
rect 6096 6560 6416 6561
rect 6096 6496 6104 6560
rect 6168 6496 6184 6560
rect 6248 6496 6264 6560
rect 6328 6496 6344 6560
rect 6408 6496 6416 6560
rect 6096 6495 6416 6496
rect 16399 6560 16719 6561
rect 16399 6496 16407 6560
rect 16471 6496 16487 6560
rect 16551 6496 16567 6560
rect 16631 6496 16647 6560
rect 16711 6496 16719 6560
rect 16399 6495 16719 6496
rect 26703 6560 27023 6561
rect 26703 6496 26711 6560
rect 26775 6496 26791 6560
rect 26855 6496 26871 6560
rect 26935 6496 26951 6560
rect 27015 6496 27023 6560
rect 26703 6495 27023 6496
rect 11247 6016 11567 6017
rect 11247 5952 11255 6016
rect 11319 5952 11335 6016
rect 11399 5952 11415 6016
rect 11479 5952 11495 6016
rect 11559 5952 11567 6016
rect 11247 5951 11567 5952
rect 21551 6016 21871 6017
rect 21551 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21799 6016
rect 21863 5952 21871 6016
rect 21551 5951 21871 5952
rect 6096 5472 6416 5473
rect 6096 5408 6104 5472
rect 6168 5408 6184 5472
rect 6248 5408 6264 5472
rect 6328 5408 6344 5472
rect 6408 5408 6416 5472
rect 6096 5407 6416 5408
rect 16399 5472 16719 5473
rect 16399 5408 16407 5472
rect 16471 5408 16487 5472
rect 16551 5408 16567 5472
rect 16631 5408 16647 5472
rect 16711 5408 16719 5472
rect 16399 5407 16719 5408
rect 26703 5472 27023 5473
rect 26703 5408 26711 5472
rect 26775 5408 26791 5472
rect 26855 5408 26871 5472
rect 26935 5408 26951 5472
rect 27015 5408 27023 5472
rect 26703 5407 27023 5408
rect 11247 4928 11567 4929
rect 11247 4864 11255 4928
rect 11319 4864 11335 4928
rect 11399 4864 11415 4928
rect 11479 4864 11495 4928
rect 11559 4864 11567 4928
rect 11247 4863 11567 4864
rect 21551 4928 21871 4929
rect 21551 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21799 4928
rect 21863 4864 21871 4928
rect 21551 4863 21871 4864
rect 6096 4384 6416 4385
rect 6096 4320 6104 4384
rect 6168 4320 6184 4384
rect 6248 4320 6264 4384
rect 6328 4320 6344 4384
rect 6408 4320 6416 4384
rect 6096 4319 6416 4320
rect 16399 4384 16719 4385
rect 16399 4320 16407 4384
rect 16471 4320 16487 4384
rect 16551 4320 16567 4384
rect 16631 4320 16647 4384
rect 16711 4320 16719 4384
rect 16399 4319 16719 4320
rect 26703 4384 27023 4385
rect 26703 4320 26711 4384
rect 26775 4320 26791 4384
rect 26855 4320 26871 4384
rect 26935 4320 26951 4384
rect 27015 4320 27023 4384
rect 26703 4319 27023 4320
rect 11247 3840 11567 3841
rect 11247 3776 11255 3840
rect 11319 3776 11335 3840
rect 11399 3776 11415 3840
rect 11479 3776 11495 3840
rect 11559 3776 11567 3840
rect 11247 3775 11567 3776
rect 21551 3840 21871 3841
rect 21551 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21799 3840
rect 21863 3776 21871 3840
rect 21551 3775 21871 3776
rect 6096 3296 6416 3297
rect 6096 3232 6104 3296
rect 6168 3232 6184 3296
rect 6248 3232 6264 3296
rect 6328 3232 6344 3296
rect 6408 3232 6416 3296
rect 6096 3231 6416 3232
rect 16399 3296 16719 3297
rect 16399 3232 16407 3296
rect 16471 3232 16487 3296
rect 16551 3232 16567 3296
rect 16631 3232 16647 3296
rect 16711 3232 16719 3296
rect 16399 3231 16719 3232
rect 26703 3296 27023 3297
rect 26703 3232 26711 3296
rect 26775 3232 26791 3296
rect 26855 3232 26871 3296
rect 26935 3232 26951 3296
rect 27015 3232 27023 3296
rect 26703 3231 27023 3232
rect 11247 2752 11567 2753
rect 11247 2688 11255 2752
rect 11319 2688 11335 2752
rect 11399 2688 11415 2752
rect 11479 2688 11495 2752
rect 11559 2688 11567 2752
rect 11247 2687 11567 2688
rect 21551 2752 21871 2753
rect 21551 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21799 2752
rect 21863 2688 21871 2752
rect 21551 2687 21871 2688
rect 6096 2208 6416 2209
rect 6096 2144 6104 2208
rect 6168 2144 6184 2208
rect 6248 2144 6264 2208
rect 6328 2144 6344 2208
rect 6408 2144 6416 2208
rect 6096 2143 6416 2144
rect 16399 2208 16719 2209
rect 16399 2144 16407 2208
rect 16471 2144 16487 2208
rect 16551 2144 16567 2208
rect 16631 2144 16647 2208
rect 16711 2144 16719 2208
rect 16399 2143 16719 2144
rect 26703 2208 27023 2209
rect 26703 2144 26711 2208
rect 26775 2144 26791 2208
rect 26855 2144 26871 2208
rect 26935 2144 26951 2208
rect 27015 2144 27023 2208
rect 26703 2143 27023 2144
rect 11247 1664 11567 1665
rect 11247 1600 11255 1664
rect 11319 1600 11335 1664
rect 11399 1600 11415 1664
rect 11479 1600 11495 1664
rect 11559 1600 11567 1664
rect 11247 1599 11567 1600
rect 21551 1664 21871 1665
rect 21551 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21799 1664
rect 21863 1600 21871 1664
rect 21551 1599 21871 1600
rect 6096 1120 6416 1121
rect 6096 1056 6104 1120
rect 6168 1056 6184 1120
rect 6248 1056 6264 1120
rect 6328 1056 6344 1120
rect 6408 1056 6416 1120
rect 6096 1055 6416 1056
rect 16399 1120 16719 1121
rect 16399 1056 16407 1120
rect 16471 1056 16487 1120
rect 16551 1056 16567 1120
rect 16631 1056 16647 1120
rect 16711 1056 16719 1120
rect 16399 1055 16719 1056
rect 26703 1120 27023 1121
rect 26703 1056 26711 1120
rect 26775 1056 26791 1120
rect 26855 1056 26871 1120
rect 26935 1056 26951 1120
rect 27015 1056 27023 1120
rect 26703 1055 27023 1056
rect 11247 576 11567 577
rect 11247 512 11255 576
rect 11319 512 11335 576
rect 11399 512 11415 576
rect 11479 512 11495 576
rect 11559 512 11567 576
rect 11247 511 11567 512
rect 21551 576 21871 577
rect 21551 512 21559 576
rect 21623 512 21639 576
rect 21703 512 21719 576
rect 21783 512 21799 576
rect 21863 512 21871 576
rect 21551 511 21871 512
<< via3 >>
rect 11255 48444 11319 48448
rect 11255 48388 11259 48444
rect 11259 48388 11315 48444
rect 11315 48388 11319 48444
rect 11255 48384 11319 48388
rect 11335 48444 11399 48448
rect 11335 48388 11339 48444
rect 11339 48388 11395 48444
rect 11395 48388 11399 48444
rect 11335 48384 11399 48388
rect 11415 48444 11479 48448
rect 11415 48388 11419 48444
rect 11419 48388 11475 48444
rect 11475 48388 11479 48444
rect 11415 48384 11479 48388
rect 11495 48444 11559 48448
rect 11495 48388 11499 48444
rect 11499 48388 11555 48444
rect 11555 48388 11559 48444
rect 11495 48384 11559 48388
rect 21559 48444 21623 48448
rect 21559 48388 21563 48444
rect 21563 48388 21619 48444
rect 21619 48388 21623 48444
rect 21559 48384 21623 48388
rect 21639 48444 21703 48448
rect 21639 48388 21643 48444
rect 21643 48388 21699 48444
rect 21699 48388 21703 48444
rect 21639 48384 21703 48388
rect 21719 48444 21783 48448
rect 21719 48388 21723 48444
rect 21723 48388 21779 48444
rect 21779 48388 21783 48444
rect 21719 48384 21783 48388
rect 21799 48444 21863 48448
rect 21799 48388 21803 48444
rect 21803 48388 21859 48444
rect 21859 48388 21863 48444
rect 21799 48384 21863 48388
rect 6104 47900 6168 47904
rect 6104 47844 6108 47900
rect 6108 47844 6164 47900
rect 6164 47844 6168 47900
rect 6104 47840 6168 47844
rect 6184 47900 6248 47904
rect 6184 47844 6188 47900
rect 6188 47844 6244 47900
rect 6244 47844 6248 47900
rect 6184 47840 6248 47844
rect 6264 47900 6328 47904
rect 6264 47844 6268 47900
rect 6268 47844 6324 47900
rect 6324 47844 6328 47900
rect 6264 47840 6328 47844
rect 6344 47900 6408 47904
rect 6344 47844 6348 47900
rect 6348 47844 6404 47900
rect 6404 47844 6408 47900
rect 6344 47840 6408 47844
rect 16407 47900 16471 47904
rect 16407 47844 16411 47900
rect 16411 47844 16467 47900
rect 16467 47844 16471 47900
rect 16407 47840 16471 47844
rect 16487 47900 16551 47904
rect 16487 47844 16491 47900
rect 16491 47844 16547 47900
rect 16547 47844 16551 47900
rect 16487 47840 16551 47844
rect 16567 47900 16631 47904
rect 16567 47844 16571 47900
rect 16571 47844 16627 47900
rect 16627 47844 16631 47900
rect 16567 47840 16631 47844
rect 16647 47900 16711 47904
rect 16647 47844 16651 47900
rect 16651 47844 16707 47900
rect 16707 47844 16711 47900
rect 16647 47840 16711 47844
rect 26711 47900 26775 47904
rect 26711 47844 26715 47900
rect 26715 47844 26771 47900
rect 26771 47844 26775 47900
rect 26711 47840 26775 47844
rect 26791 47900 26855 47904
rect 26791 47844 26795 47900
rect 26795 47844 26851 47900
rect 26851 47844 26855 47900
rect 26791 47840 26855 47844
rect 26871 47900 26935 47904
rect 26871 47844 26875 47900
rect 26875 47844 26931 47900
rect 26931 47844 26935 47900
rect 26871 47840 26935 47844
rect 26951 47900 27015 47904
rect 26951 47844 26955 47900
rect 26955 47844 27011 47900
rect 27011 47844 27015 47900
rect 26951 47840 27015 47844
rect 11255 47356 11319 47360
rect 11255 47300 11259 47356
rect 11259 47300 11315 47356
rect 11315 47300 11319 47356
rect 11255 47296 11319 47300
rect 11335 47356 11399 47360
rect 11335 47300 11339 47356
rect 11339 47300 11395 47356
rect 11395 47300 11399 47356
rect 11335 47296 11399 47300
rect 11415 47356 11479 47360
rect 11415 47300 11419 47356
rect 11419 47300 11475 47356
rect 11475 47300 11479 47356
rect 11415 47296 11479 47300
rect 11495 47356 11559 47360
rect 11495 47300 11499 47356
rect 11499 47300 11555 47356
rect 11555 47300 11559 47356
rect 11495 47296 11559 47300
rect 21559 47356 21623 47360
rect 21559 47300 21563 47356
rect 21563 47300 21619 47356
rect 21619 47300 21623 47356
rect 21559 47296 21623 47300
rect 21639 47356 21703 47360
rect 21639 47300 21643 47356
rect 21643 47300 21699 47356
rect 21699 47300 21703 47356
rect 21639 47296 21703 47300
rect 21719 47356 21783 47360
rect 21719 47300 21723 47356
rect 21723 47300 21779 47356
rect 21779 47300 21783 47356
rect 21719 47296 21783 47300
rect 21799 47356 21863 47360
rect 21799 47300 21803 47356
rect 21803 47300 21859 47356
rect 21859 47300 21863 47356
rect 21799 47296 21863 47300
rect 6104 46812 6168 46816
rect 6104 46756 6108 46812
rect 6108 46756 6164 46812
rect 6164 46756 6168 46812
rect 6104 46752 6168 46756
rect 6184 46812 6248 46816
rect 6184 46756 6188 46812
rect 6188 46756 6244 46812
rect 6244 46756 6248 46812
rect 6184 46752 6248 46756
rect 6264 46812 6328 46816
rect 6264 46756 6268 46812
rect 6268 46756 6324 46812
rect 6324 46756 6328 46812
rect 6264 46752 6328 46756
rect 6344 46812 6408 46816
rect 6344 46756 6348 46812
rect 6348 46756 6404 46812
rect 6404 46756 6408 46812
rect 6344 46752 6408 46756
rect 16407 46812 16471 46816
rect 16407 46756 16411 46812
rect 16411 46756 16467 46812
rect 16467 46756 16471 46812
rect 16407 46752 16471 46756
rect 16487 46812 16551 46816
rect 16487 46756 16491 46812
rect 16491 46756 16547 46812
rect 16547 46756 16551 46812
rect 16487 46752 16551 46756
rect 16567 46812 16631 46816
rect 16567 46756 16571 46812
rect 16571 46756 16627 46812
rect 16627 46756 16631 46812
rect 16567 46752 16631 46756
rect 16647 46812 16711 46816
rect 16647 46756 16651 46812
rect 16651 46756 16707 46812
rect 16707 46756 16711 46812
rect 16647 46752 16711 46756
rect 26711 46812 26775 46816
rect 26711 46756 26715 46812
rect 26715 46756 26771 46812
rect 26771 46756 26775 46812
rect 26711 46752 26775 46756
rect 26791 46812 26855 46816
rect 26791 46756 26795 46812
rect 26795 46756 26851 46812
rect 26851 46756 26855 46812
rect 26791 46752 26855 46756
rect 26871 46812 26935 46816
rect 26871 46756 26875 46812
rect 26875 46756 26931 46812
rect 26931 46756 26935 46812
rect 26871 46752 26935 46756
rect 26951 46812 27015 46816
rect 26951 46756 26955 46812
rect 26955 46756 27011 46812
rect 27011 46756 27015 46812
rect 26951 46752 27015 46756
rect 11255 46268 11319 46272
rect 11255 46212 11259 46268
rect 11259 46212 11315 46268
rect 11315 46212 11319 46268
rect 11255 46208 11319 46212
rect 11335 46268 11399 46272
rect 11335 46212 11339 46268
rect 11339 46212 11395 46268
rect 11395 46212 11399 46268
rect 11335 46208 11399 46212
rect 11415 46268 11479 46272
rect 11415 46212 11419 46268
rect 11419 46212 11475 46268
rect 11475 46212 11479 46268
rect 11415 46208 11479 46212
rect 11495 46268 11559 46272
rect 11495 46212 11499 46268
rect 11499 46212 11555 46268
rect 11555 46212 11559 46268
rect 11495 46208 11559 46212
rect 21559 46268 21623 46272
rect 21559 46212 21563 46268
rect 21563 46212 21619 46268
rect 21619 46212 21623 46268
rect 21559 46208 21623 46212
rect 21639 46268 21703 46272
rect 21639 46212 21643 46268
rect 21643 46212 21699 46268
rect 21699 46212 21703 46268
rect 21639 46208 21703 46212
rect 21719 46268 21783 46272
rect 21719 46212 21723 46268
rect 21723 46212 21779 46268
rect 21779 46212 21783 46268
rect 21719 46208 21783 46212
rect 21799 46268 21863 46272
rect 21799 46212 21803 46268
rect 21803 46212 21859 46268
rect 21859 46212 21863 46268
rect 21799 46208 21863 46212
rect 6104 45724 6168 45728
rect 6104 45668 6108 45724
rect 6108 45668 6164 45724
rect 6164 45668 6168 45724
rect 6104 45664 6168 45668
rect 6184 45724 6248 45728
rect 6184 45668 6188 45724
rect 6188 45668 6244 45724
rect 6244 45668 6248 45724
rect 6184 45664 6248 45668
rect 6264 45724 6328 45728
rect 6264 45668 6268 45724
rect 6268 45668 6324 45724
rect 6324 45668 6328 45724
rect 6264 45664 6328 45668
rect 6344 45724 6408 45728
rect 6344 45668 6348 45724
rect 6348 45668 6404 45724
rect 6404 45668 6408 45724
rect 6344 45664 6408 45668
rect 16407 45724 16471 45728
rect 16407 45668 16411 45724
rect 16411 45668 16467 45724
rect 16467 45668 16471 45724
rect 16407 45664 16471 45668
rect 16487 45724 16551 45728
rect 16487 45668 16491 45724
rect 16491 45668 16547 45724
rect 16547 45668 16551 45724
rect 16487 45664 16551 45668
rect 16567 45724 16631 45728
rect 16567 45668 16571 45724
rect 16571 45668 16627 45724
rect 16627 45668 16631 45724
rect 16567 45664 16631 45668
rect 16647 45724 16711 45728
rect 16647 45668 16651 45724
rect 16651 45668 16707 45724
rect 16707 45668 16711 45724
rect 16647 45664 16711 45668
rect 26711 45724 26775 45728
rect 26711 45668 26715 45724
rect 26715 45668 26771 45724
rect 26771 45668 26775 45724
rect 26711 45664 26775 45668
rect 26791 45724 26855 45728
rect 26791 45668 26795 45724
rect 26795 45668 26851 45724
rect 26851 45668 26855 45724
rect 26791 45664 26855 45668
rect 26871 45724 26935 45728
rect 26871 45668 26875 45724
rect 26875 45668 26931 45724
rect 26931 45668 26935 45724
rect 26871 45664 26935 45668
rect 26951 45724 27015 45728
rect 26951 45668 26955 45724
rect 26955 45668 27011 45724
rect 27011 45668 27015 45724
rect 26951 45664 27015 45668
rect 11255 45180 11319 45184
rect 11255 45124 11259 45180
rect 11259 45124 11315 45180
rect 11315 45124 11319 45180
rect 11255 45120 11319 45124
rect 11335 45180 11399 45184
rect 11335 45124 11339 45180
rect 11339 45124 11395 45180
rect 11395 45124 11399 45180
rect 11335 45120 11399 45124
rect 11415 45180 11479 45184
rect 11415 45124 11419 45180
rect 11419 45124 11475 45180
rect 11475 45124 11479 45180
rect 11415 45120 11479 45124
rect 11495 45180 11559 45184
rect 11495 45124 11499 45180
rect 11499 45124 11555 45180
rect 11555 45124 11559 45180
rect 11495 45120 11559 45124
rect 21559 45180 21623 45184
rect 21559 45124 21563 45180
rect 21563 45124 21619 45180
rect 21619 45124 21623 45180
rect 21559 45120 21623 45124
rect 21639 45180 21703 45184
rect 21639 45124 21643 45180
rect 21643 45124 21699 45180
rect 21699 45124 21703 45180
rect 21639 45120 21703 45124
rect 21719 45180 21783 45184
rect 21719 45124 21723 45180
rect 21723 45124 21779 45180
rect 21779 45124 21783 45180
rect 21719 45120 21783 45124
rect 21799 45180 21863 45184
rect 21799 45124 21803 45180
rect 21803 45124 21859 45180
rect 21859 45124 21863 45180
rect 21799 45120 21863 45124
rect 6104 44636 6168 44640
rect 6104 44580 6108 44636
rect 6108 44580 6164 44636
rect 6164 44580 6168 44636
rect 6104 44576 6168 44580
rect 6184 44636 6248 44640
rect 6184 44580 6188 44636
rect 6188 44580 6244 44636
rect 6244 44580 6248 44636
rect 6184 44576 6248 44580
rect 6264 44636 6328 44640
rect 6264 44580 6268 44636
rect 6268 44580 6324 44636
rect 6324 44580 6328 44636
rect 6264 44576 6328 44580
rect 6344 44636 6408 44640
rect 6344 44580 6348 44636
rect 6348 44580 6404 44636
rect 6404 44580 6408 44636
rect 6344 44576 6408 44580
rect 16407 44636 16471 44640
rect 16407 44580 16411 44636
rect 16411 44580 16467 44636
rect 16467 44580 16471 44636
rect 16407 44576 16471 44580
rect 16487 44636 16551 44640
rect 16487 44580 16491 44636
rect 16491 44580 16547 44636
rect 16547 44580 16551 44636
rect 16487 44576 16551 44580
rect 16567 44636 16631 44640
rect 16567 44580 16571 44636
rect 16571 44580 16627 44636
rect 16627 44580 16631 44636
rect 16567 44576 16631 44580
rect 16647 44636 16711 44640
rect 16647 44580 16651 44636
rect 16651 44580 16707 44636
rect 16707 44580 16711 44636
rect 16647 44576 16711 44580
rect 26711 44636 26775 44640
rect 26711 44580 26715 44636
rect 26715 44580 26771 44636
rect 26771 44580 26775 44636
rect 26711 44576 26775 44580
rect 26791 44636 26855 44640
rect 26791 44580 26795 44636
rect 26795 44580 26851 44636
rect 26851 44580 26855 44636
rect 26791 44576 26855 44580
rect 26871 44636 26935 44640
rect 26871 44580 26875 44636
rect 26875 44580 26931 44636
rect 26931 44580 26935 44636
rect 26871 44576 26935 44580
rect 26951 44636 27015 44640
rect 26951 44580 26955 44636
rect 26955 44580 27011 44636
rect 27011 44580 27015 44636
rect 26951 44576 27015 44580
rect 11255 44092 11319 44096
rect 11255 44036 11259 44092
rect 11259 44036 11315 44092
rect 11315 44036 11319 44092
rect 11255 44032 11319 44036
rect 11335 44092 11399 44096
rect 11335 44036 11339 44092
rect 11339 44036 11395 44092
rect 11395 44036 11399 44092
rect 11335 44032 11399 44036
rect 11415 44092 11479 44096
rect 11415 44036 11419 44092
rect 11419 44036 11475 44092
rect 11475 44036 11479 44092
rect 11415 44032 11479 44036
rect 11495 44092 11559 44096
rect 11495 44036 11499 44092
rect 11499 44036 11555 44092
rect 11555 44036 11559 44092
rect 11495 44032 11559 44036
rect 21559 44092 21623 44096
rect 21559 44036 21563 44092
rect 21563 44036 21619 44092
rect 21619 44036 21623 44092
rect 21559 44032 21623 44036
rect 21639 44092 21703 44096
rect 21639 44036 21643 44092
rect 21643 44036 21699 44092
rect 21699 44036 21703 44092
rect 21639 44032 21703 44036
rect 21719 44092 21783 44096
rect 21719 44036 21723 44092
rect 21723 44036 21779 44092
rect 21779 44036 21783 44092
rect 21719 44032 21783 44036
rect 21799 44092 21863 44096
rect 21799 44036 21803 44092
rect 21803 44036 21859 44092
rect 21859 44036 21863 44092
rect 21799 44032 21863 44036
rect 6104 43548 6168 43552
rect 6104 43492 6108 43548
rect 6108 43492 6164 43548
rect 6164 43492 6168 43548
rect 6104 43488 6168 43492
rect 6184 43548 6248 43552
rect 6184 43492 6188 43548
rect 6188 43492 6244 43548
rect 6244 43492 6248 43548
rect 6184 43488 6248 43492
rect 6264 43548 6328 43552
rect 6264 43492 6268 43548
rect 6268 43492 6324 43548
rect 6324 43492 6328 43548
rect 6264 43488 6328 43492
rect 6344 43548 6408 43552
rect 6344 43492 6348 43548
rect 6348 43492 6404 43548
rect 6404 43492 6408 43548
rect 6344 43488 6408 43492
rect 16407 43548 16471 43552
rect 16407 43492 16411 43548
rect 16411 43492 16467 43548
rect 16467 43492 16471 43548
rect 16407 43488 16471 43492
rect 16487 43548 16551 43552
rect 16487 43492 16491 43548
rect 16491 43492 16547 43548
rect 16547 43492 16551 43548
rect 16487 43488 16551 43492
rect 16567 43548 16631 43552
rect 16567 43492 16571 43548
rect 16571 43492 16627 43548
rect 16627 43492 16631 43548
rect 16567 43488 16631 43492
rect 16647 43548 16711 43552
rect 16647 43492 16651 43548
rect 16651 43492 16707 43548
rect 16707 43492 16711 43548
rect 16647 43488 16711 43492
rect 26711 43548 26775 43552
rect 26711 43492 26715 43548
rect 26715 43492 26771 43548
rect 26771 43492 26775 43548
rect 26711 43488 26775 43492
rect 26791 43548 26855 43552
rect 26791 43492 26795 43548
rect 26795 43492 26851 43548
rect 26851 43492 26855 43548
rect 26791 43488 26855 43492
rect 26871 43548 26935 43552
rect 26871 43492 26875 43548
rect 26875 43492 26931 43548
rect 26931 43492 26935 43548
rect 26871 43488 26935 43492
rect 26951 43548 27015 43552
rect 26951 43492 26955 43548
rect 26955 43492 27011 43548
rect 27011 43492 27015 43548
rect 26951 43488 27015 43492
rect 11255 43004 11319 43008
rect 11255 42948 11259 43004
rect 11259 42948 11315 43004
rect 11315 42948 11319 43004
rect 11255 42944 11319 42948
rect 11335 43004 11399 43008
rect 11335 42948 11339 43004
rect 11339 42948 11395 43004
rect 11395 42948 11399 43004
rect 11335 42944 11399 42948
rect 11415 43004 11479 43008
rect 11415 42948 11419 43004
rect 11419 42948 11475 43004
rect 11475 42948 11479 43004
rect 11415 42944 11479 42948
rect 11495 43004 11559 43008
rect 11495 42948 11499 43004
rect 11499 42948 11555 43004
rect 11555 42948 11559 43004
rect 11495 42944 11559 42948
rect 21559 43004 21623 43008
rect 21559 42948 21563 43004
rect 21563 42948 21619 43004
rect 21619 42948 21623 43004
rect 21559 42944 21623 42948
rect 21639 43004 21703 43008
rect 21639 42948 21643 43004
rect 21643 42948 21699 43004
rect 21699 42948 21703 43004
rect 21639 42944 21703 42948
rect 21719 43004 21783 43008
rect 21719 42948 21723 43004
rect 21723 42948 21779 43004
rect 21779 42948 21783 43004
rect 21719 42944 21783 42948
rect 21799 43004 21863 43008
rect 21799 42948 21803 43004
rect 21803 42948 21859 43004
rect 21859 42948 21863 43004
rect 21799 42944 21863 42948
rect 6104 42460 6168 42464
rect 6104 42404 6108 42460
rect 6108 42404 6164 42460
rect 6164 42404 6168 42460
rect 6104 42400 6168 42404
rect 6184 42460 6248 42464
rect 6184 42404 6188 42460
rect 6188 42404 6244 42460
rect 6244 42404 6248 42460
rect 6184 42400 6248 42404
rect 6264 42460 6328 42464
rect 6264 42404 6268 42460
rect 6268 42404 6324 42460
rect 6324 42404 6328 42460
rect 6264 42400 6328 42404
rect 6344 42460 6408 42464
rect 6344 42404 6348 42460
rect 6348 42404 6404 42460
rect 6404 42404 6408 42460
rect 6344 42400 6408 42404
rect 16407 42460 16471 42464
rect 16407 42404 16411 42460
rect 16411 42404 16467 42460
rect 16467 42404 16471 42460
rect 16407 42400 16471 42404
rect 16487 42460 16551 42464
rect 16487 42404 16491 42460
rect 16491 42404 16547 42460
rect 16547 42404 16551 42460
rect 16487 42400 16551 42404
rect 16567 42460 16631 42464
rect 16567 42404 16571 42460
rect 16571 42404 16627 42460
rect 16627 42404 16631 42460
rect 16567 42400 16631 42404
rect 16647 42460 16711 42464
rect 16647 42404 16651 42460
rect 16651 42404 16707 42460
rect 16707 42404 16711 42460
rect 16647 42400 16711 42404
rect 26711 42460 26775 42464
rect 26711 42404 26715 42460
rect 26715 42404 26771 42460
rect 26771 42404 26775 42460
rect 26711 42400 26775 42404
rect 26791 42460 26855 42464
rect 26791 42404 26795 42460
rect 26795 42404 26851 42460
rect 26851 42404 26855 42460
rect 26791 42400 26855 42404
rect 26871 42460 26935 42464
rect 26871 42404 26875 42460
rect 26875 42404 26931 42460
rect 26931 42404 26935 42460
rect 26871 42400 26935 42404
rect 26951 42460 27015 42464
rect 26951 42404 26955 42460
rect 26955 42404 27011 42460
rect 27011 42404 27015 42460
rect 26951 42400 27015 42404
rect 11255 41916 11319 41920
rect 11255 41860 11259 41916
rect 11259 41860 11315 41916
rect 11315 41860 11319 41916
rect 11255 41856 11319 41860
rect 11335 41916 11399 41920
rect 11335 41860 11339 41916
rect 11339 41860 11395 41916
rect 11395 41860 11399 41916
rect 11335 41856 11399 41860
rect 11415 41916 11479 41920
rect 11415 41860 11419 41916
rect 11419 41860 11475 41916
rect 11475 41860 11479 41916
rect 11415 41856 11479 41860
rect 11495 41916 11559 41920
rect 11495 41860 11499 41916
rect 11499 41860 11555 41916
rect 11555 41860 11559 41916
rect 11495 41856 11559 41860
rect 21559 41916 21623 41920
rect 21559 41860 21563 41916
rect 21563 41860 21619 41916
rect 21619 41860 21623 41916
rect 21559 41856 21623 41860
rect 21639 41916 21703 41920
rect 21639 41860 21643 41916
rect 21643 41860 21699 41916
rect 21699 41860 21703 41916
rect 21639 41856 21703 41860
rect 21719 41916 21783 41920
rect 21719 41860 21723 41916
rect 21723 41860 21779 41916
rect 21779 41860 21783 41916
rect 21719 41856 21783 41860
rect 21799 41916 21863 41920
rect 21799 41860 21803 41916
rect 21803 41860 21859 41916
rect 21859 41860 21863 41916
rect 21799 41856 21863 41860
rect 6104 41372 6168 41376
rect 6104 41316 6108 41372
rect 6108 41316 6164 41372
rect 6164 41316 6168 41372
rect 6104 41312 6168 41316
rect 6184 41372 6248 41376
rect 6184 41316 6188 41372
rect 6188 41316 6244 41372
rect 6244 41316 6248 41372
rect 6184 41312 6248 41316
rect 6264 41372 6328 41376
rect 6264 41316 6268 41372
rect 6268 41316 6324 41372
rect 6324 41316 6328 41372
rect 6264 41312 6328 41316
rect 6344 41372 6408 41376
rect 6344 41316 6348 41372
rect 6348 41316 6404 41372
rect 6404 41316 6408 41372
rect 6344 41312 6408 41316
rect 16407 41372 16471 41376
rect 16407 41316 16411 41372
rect 16411 41316 16467 41372
rect 16467 41316 16471 41372
rect 16407 41312 16471 41316
rect 16487 41372 16551 41376
rect 16487 41316 16491 41372
rect 16491 41316 16547 41372
rect 16547 41316 16551 41372
rect 16487 41312 16551 41316
rect 16567 41372 16631 41376
rect 16567 41316 16571 41372
rect 16571 41316 16627 41372
rect 16627 41316 16631 41372
rect 16567 41312 16631 41316
rect 16647 41372 16711 41376
rect 16647 41316 16651 41372
rect 16651 41316 16707 41372
rect 16707 41316 16711 41372
rect 16647 41312 16711 41316
rect 26711 41372 26775 41376
rect 26711 41316 26715 41372
rect 26715 41316 26771 41372
rect 26771 41316 26775 41372
rect 26711 41312 26775 41316
rect 26791 41372 26855 41376
rect 26791 41316 26795 41372
rect 26795 41316 26851 41372
rect 26851 41316 26855 41372
rect 26791 41312 26855 41316
rect 26871 41372 26935 41376
rect 26871 41316 26875 41372
rect 26875 41316 26931 41372
rect 26931 41316 26935 41372
rect 26871 41312 26935 41316
rect 26951 41372 27015 41376
rect 26951 41316 26955 41372
rect 26955 41316 27011 41372
rect 27011 41316 27015 41372
rect 26951 41312 27015 41316
rect 11255 40828 11319 40832
rect 11255 40772 11259 40828
rect 11259 40772 11315 40828
rect 11315 40772 11319 40828
rect 11255 40768 11319 40772
rect 11335 40828 11399 40832
rect 11335 40772 11339 40828
rect 11339 40772 11395 40828
rect 11395 40772 11399 40828
rect 11335 40768 11399 40772
rect 11415 40828 11479 40832
rect 11415 40772 11419 40828
rect 11419 40772 11475 40828
rect 11475 40772 11479 40828
rect 11415 40768 11479 40772
rect 11495 40828 11559 40832
rect 11495 40772 11499 40828
rect 11499 40772 11555 40828
rect 11555 40772 11559 40828
rect 11495 40768 11559 40772
rect 21559 40828 21623 40832
rect 21559 40772 21563 40828
rect 21563 40772 21619 40828
rect 21619 40772 21623 40828
rect 21559 40768 21623 40772
rect 21639 40828 21703 40832
rect 21639 40772 21643 40828
rect 21643 40772 21699 40828
rect 21699 40772 21703 40828
rect 21639 40768 21703 40772
rect 21719 40828 21783 40832
rect 21719 40772 21723 40828
rect 21723 40772 21779 40828
rect 21779 40772 21783 40828
rect 21719 40768 21783 40772
rect 21799 40828 21863 40832
rect 21799 40772 21803 40828
rect 21803 40772 21859 40828
rect 21859 40772 21863 40828
rect 21799 40768 21863 40772
rect 6104 40284 6168 40288
rect 6104 40228 6108 40284
rect 6108 40228 6164 40284
rect 6164 40228 6168 40284
rect 6104 40224 6168 40228
rect 6184 40284 6248 40288
rect 6184 40228 6188 40284
rect 6188 40228 6244 40284
rect 6244 40228 6248 40284
rect 6184 40224 6248 40228
rect 6264 40284 6328 40288
rect 6264 40228 6268 40284
rect 6268 40228 6324 40284
rect 6324 40228 6328 40284
rect 6264 40224 6328 40228
rect 6344 40284 6408 40288
rect 6344 40228 6348 40284
rect 6348 40228 6404 40284
rect 6404 40228 6408 40284
rect 6344 40224 6408 40228
rect 16407 40284 16471 40288
rect 16407 40228 16411 40284
rect 16411 40228 16467 40284
rect 16467 40228 16471 40284
rect 16407 40224 16471 40228
rect 16487 40284 16551 40288
rect 16487 40228 16491 40284
rect 16491 40228 16547 40284
rect 16547 40228 16551 40284
rect 16487 40224 16551 40228
rect 16567 40284 16631 40288
rect 16567 40228 16571 40284
rect 16571 40228 16627 40284
rect 16627 40228 16631 40284
rect 16567 40224 16631 40228
rect 16647 40284 16711 40288
rect 16647 40228 16651 40284
rect 16651 40228 16707 40284
rect 16707 40228 16711 40284
rect 16647 40224 16711 40228
rect 26711 40284 26775 40288
rect 26711 40228 26715 40284
rect 26715 40228 26771 40284
rect 26771 40228 26775 40284
rect 26711 40224 26775 40228
rect 26791 40284 26855 40288
rect 26791 40228 26795 40284
rect 26795 40228 26851 40284
rect 26851 40228 26855 40284
rect 26791 40224 26855 40228
rect 26871 40284 26935 40288
rect 26871 40228 26875 40284
rect 26875 40228 26931 40284
rect 26931 40228 26935 40284
rect 26871 40224 26935 40228
rect 26951 40284 27015 40288
rect 26951 40228 26955 40284
rect 26955 40228 27011 40284
rect 27011 40228 27015 40284
rect 26951 40224 27015 40228
rect 11255 39740 11319 39744
rect 11255 39684 11259 39740
rect 11259 39684 11315 39740
rect 11315 39684 11319 39740
rect 11255 39680 11319 39684
rect 11335 39740 11399 39744
rect 11335 39684 11339 39740
rect 11339 39684 11395 39740
rect 11395 39684 11399 39740
rect 11335 39680 11399 39684
rect 11415 39740 11479 39744
rect 11415 39684 11419 39740
rect 11419 39684 11475 39740
rect 11475 39684 11479 39740
rect 11415 39680 11479 39684
rect 11495 39740 11559 39744
rect 11495 39684 11499 39740
rect 11499 39684 11555 39740
rect 11555 39684 11559 39740
rect 11495 39680 11559 39684
rect 21559 39740 21623 39744
rect 21559 39684 21563 39740
rect 21563 39684 21619 39740
rect 21619 39684 21623 39740
rect 21559 39680 21623 39684
rect 21639 39740 21703 39744
rect 21639 39684 21643 39740
rect 21643 39684 21699 39740
rect 21699 39684 21703 39740
rect 21639 39680 21703 39684
rect 21719 39740 21783 39744
rect 21719 39684 21723 39740
rect 21723 39684 21779 39740
rect 21779 39684 21783 39740
rect 21719 39680 21783 39684
rect 21799 39740 21863 39744
rect 21799 39684 21803 39740
rect 21803 39684 21859 39740
rect 21859 39684 21863 39740
rect 21799 39680 21863 39684
rect 6104 39196 6168 39200
rect 6104 39140 6108 39196
rect 6108 39140 6164 39196
rect 6164 39140 6168 39196
rect 6104 39136 6168 39140
rect 6184 39196 6248 39200
rect 6184 39140 6188 39196
rect 6188 39140 6244 39196
rect 6244 39140 6248 39196
rect 6184 39136 6248 39140
rect 6264 39196 6328 39200
rect 6264 39140 6268 39196
rect 6268 39140 6324 39196
rect 6324 39140 6328 39196
rect 6264 39136 6328 39140
rect 6344 39196 6408 39200
rect 6344 39140 6348 39196
rect 6348 39140 6404 39196
rect 6404 39140 6408 39196
rect 6344 39136 6408 39140
rect 16407 39196 16471 39200
rect 16407 39140 16411 39196
rect 16411 39140 16467 39196
rect 16467 39140 16471 39196
rect 16407 39136 16471 39140
rect 16487 39196 16551 39200
rect 16487 39140 16491 39196
rect 16491 39140 16547 39196
rect 16547 39140 16551 39196
rect 16487 39136 16551 39140
rect 16567 39196 16631 39200
rect 16567 39140 16571 39196
rect 16571 39140 16627 39196
rect 16627 39140 16631 39196
rect 16567 39136 16631 39140
rect 16647 39196 16711 39200
rect 16647 39140 16651 39196
rect 16651 39140 16707 39196
rect 16707 39140 16711 39196
rect 16647 39136 16711 39140
rect 26711 39196 26775 39200
rect 26711 39140 26715 39196
rect 26715 39140 26771 39196
rect 26771 39140 26775 39196
rect 26711 39136 26775 39140
rect 26791 39196 26855 39200
rect 26791 39140 26795 39196
rect 26795 39140 26851 39196
rect 26851 39140 26855 39196
rect 26791 39136 26855 39140
rect 26871 39196 26935 39200
rect 26871 39140 26875 39196
rect 26875 39140 26931 39196
rect 26931 39140 26935 39196
rect 26871 39136 26935 39140
rect 26951 39196 27015 39200
rect 26951 39140 26955 39196
rect 26955 39140 27011 39196
rect 27011 39140 27015 39196
rect 26951 39136 27015 39140
rect 11255 38652 11319 38656
rect 11255 38596 11259 38652
rect 11259 38596 11315 38652
rect 11315 38596 11319 38652
rect 11255 38592 11319 38596
rect 11335 38652 11399 38656
rect 11335 38596 11339 38652
rect 11339 38596 11395 38652
rect 11395 38596 11399 38652
rect 11335 38592 11399 38596
rect 11415 38652 11479 38656
rect 11415 38596 11419 38652
rect 11419 38596 11475 38652
rect 11475 38596 11479 38652
rect 11415 38592 11479 38596
rect 11495 38652 11559 38656
rect 11495 38596 11499 38652
rect 11499 38596 11555 38652
rect 11555 38596 11559 38652
rect 11495 38592 11559 38596
rect 21559 38652 21623 38656
rect 21559 38596 21563 38652
rect 21563 38596 21619 38652
rect 21619 38596 21623 38652
rect 21559 38592 21623 38596
rect 21639 38652 21703 38656
rect 21639 38596 21643 38652
rect 21643 38596 21699 38652
rect 21699 38596 21703 38652
rect 21639 38592 21703 38596
rect 21719 38652 21783 38656
rect 21719 38596 21723 38652
rect 21723 38596 21779 38652
rect 21779 38596 21783 38652
rect 21719 38592 21783 38596
rect 21799 38652 21863 38656
rect 21799 38596 21803 38652
rect 21803 38596 21859 38652
rect 21859 38596 21863 38652
rect 21799 38592 21863 38596
rect 6104 38108 6168 38112
rect 6104 38052 6108 38108
rect 6108 38052 6164 38108
rect 6164 38052 6168 38108
rect 6104 38048 6168 38052
rect 6184 38108 6248 38112
rect 6184 38052 6188 38108
rect 6188 38052 6244 38108
rect 6244 38052 6248 38108
rect 6184 38048 6248 38052
rect 6264 38108 6328 38112
rect 6264 38052 6268 38108
rect 6268 38052 6324 38108
rect 6324 38052 6328 38108
rect 6264 38048 6328 38052
rect 6344 38108 6408 38112
rect 6344 38052 6348 38108
rect 6348 38052 6404 38108
rect 6404 38052 6408 38108
rect 6344 38048 6408 38052
rect 16407 38108 16471 38112
rect 16407 38052 16411 38108
rect 16411 38052 16467 38108
rect 16467 38052 16471 38108
rect 16407 38048 16471 38052
rect 16487 38108 16551 38112
rect 16487 38052 16491 38108
rect 16491 38052 16547 38108
rect 16547 38052 16551 38108
rect 16487 38048 16551 38052
rect 16567 38108 16631 38112
rect 16567 38052 16571 38108
rect 16571 38052 16627 38108
rect 16627 38052 16631 38108
rect 16567 38048 16631 38052
rect 16647 38108 16711 38112
rect 16647 38052 16651 38108
rect 16651 38052 16707 38108
rect 16707 38052 16711 38108
rect 16647 38048 16711 38052
rect 26711 38108 26775 38112
rect 26711 38052 26715 38108
rect 26715 38052 26771 38108
rect 26771 38052 26775 38108
rect 26711 38048 26775 38052
rect 26791 38108 26855 38112
rect 26791 38052 26795 38108
rect 26795 38052 26851 38108
rect 26851 38052 26855 38108
rect 26791 38048 26855 38052
rect 26871 38108 26935 38112
rect 26871 38052 26875 38108
rect 26875 38052 26931 38108
rect 26931 38052 26935 38108
rect 26871 38048 26935 38052
rect 26951 38108 27015 38112
rect 26951 38052 26955 38108
rect 26955 38052 27011 38108
rect 27011 38052 27015 38108
rect 26951 38048 27015 38052
rect 11255 37564 11319 37568
rect 11255 37508 11259 37564
rect 11259 37508 11315 37564
rect 11315 37508 11319 37564
rect 11255 37504 11319 37508
rect 11335 37564 11399 37568
rect 11335 37508 11339 37564
rect 11339 37508 11395 37564
rect 11395 37508 11399 37564
rect 11335 37504 11399 37508
rect 11415 37564 11479 37568
rect 11415 37508 11419 37564
rect 11419 37508 11475 37564
rect 11475 37508 11479 37564
rect 11415 37504 11479 37508
rect 11495 37564 11559 37568
rect 11495 37508 11499 37564
rect 11499 37508 11555 37564
rect 11555 37508 11559 37564
rect 11495 37504 11559 37508
rect 21559 37564 21623 37568
rect 21559 37508 21563 37564
rect 21563 37508 21619 37564
rect 21619 37508 21623 37564
rect 21559 37504 21623 37508
rect 21639 37564 21703 37568
rect 21639 37508 21643 37564
rect 21643 37508 21699 37564
rect 21699 37508 21703 37564
rect 21639 37504 21703 37508
rect 21719 37564 21783 37568
rect 21719 37508 21723 37564
rect 21723 37508 21779 37564
rect 21779 37508 21783 37564
rect 21719 37504 21783 37508
rect 21799 37564 21863 37568
rect 21799 37508 21803 37564
rect 21803 37508 21859 37564
rect 21859 37508 21863 37564
rect 21799 37504 21863 37508
rect 6104 37020 6168 37024
rect 6104 36964 6108 37020
rect 6108 36964 6164 37020
rect 6164 36964 6168 37020
rect 6104 36960 6168 36964
rect 6184 37020 6248 37024
rect 6184 36964 6188 37020
rect 6188 36964 6244 37020
rect 6244 36964 6248 37020
rect 6184 36960 6248 36964
rect 6264 37020 6328 37024
rect 6264 36964 6268 37020
rect 6268 36964 6324 37020
rect 6324 36964 6328 37020
rect 6264 36960 6328 36964
rect 6344 37020 6408 37024
rect 6344 36964 6348 37020
rect 6348 36964 6404 37020
rect 6404 36964 6408 37020
rect 6344 36960 6408 36964
rect 16407 37020 16471 37024
rect 16407 36964 16411 37020
rect 16411 36964 16467 37020
rect 16467 36964 16471 37020
rect 16407 36960 16471 36964
rect 16487 37020 16551 37024
rect 16487 36964 16491 37020
rect 16491 36964 16547 37020
rect 16547 36964 16551 37020
rect 16487 36960 16551 36964
rect 16567 37020 16631 37024
rect 16567 36964 16571 37020
rect 16571 36964 16627 37020
rect 16627 36964 16631 37020
rect 16567 36960 16631 36964
rect 16647 37020 16711 37024
rect 16647 36964 16651 37020
rect 16651 36964 16707 37020
rect 16707 36964 16711 37020
rect 16647 36960 16711 36964
rect 26711 37020 26775 37024
rect 26711 36964 26715 37020
rect 26715 36964 26771 37020
rect 26771 36964 26775 37020
rect 26711 36960 26775 36964
rect 26791 37020 26855 37024
rect 26791 36964 26795 37020
rect 26795 36964 26851 37020
rect 26851 36964 26855 37020
rect 26791 36960 26855 36964
rect 26871 37020 26935 37024
rect 26871 36964 26875 37020
rect 26875 36964 26931 37020
rect 26931 36964 26935 37020
rect 26871 36960 26935 36964
rect 26951 37020 27015 37024
rect 26951 36964 26955 37020
rect 26955 36964 27011 37020
rect 27011 36964 27015 37020
rect 26951 36960 27015 36964
rect 11255 36476 11319 36480
rect 11255 36420 11259 36476
rect 11259 36420 11315 36476
rect 11315 36420 11319 36476
rect 11255 36416 11319 36420
rect 11335 36476 11399 36480
rect 11335 36420 11339 36476
rect 11339 36420 11395 36476
rect 11395 36420 11399 36476
rect 11335 36416 11399 36420
rect 11415 36476 11479 36480
rect 11415 36420 11419 36476
rect 11419 36420 11475 36476
rect 11475 36420 11479 36476
rect 11415 36416 11479 36420
rect 11495 36476 11559 36480
rect 11495 36420 11499 36476
rect 11499 36420 11555 36476
rect 11555 36420 11559 36476
rect 11495 36416 11559 36420
rect 21559 36476 21623 36480
rect 21559 36420 21563 36476
rect 21563 36420 21619 36476
rect 21619 36420 21623 36476
rect 21559 36416 21623 36420
rect 21639 36476 21703 36480
rect 21639 36420 21643 36476
rect 21643 36420 21699 36476
rect 21699 36420 21703 36476
rect 21639 36416 21703 36420
rect 21719 36476 21783 36480
rect 21719 36420 21723 36476
rect 21723 36420 21779 36476
rect 21779 36420 21783 36476
rect 21719 36416 21783 36420
rect 21799 36476 21863 36480
rect 21799 36420 21803 36476
rect 21803 36420 21859 36476
rect 21859 36420 21863 36476
rect 21799 36416 21863 36420
rect 6104 35932 6168 35936
rect 6104 35876 6108 35932
rect 6108 35876 6164 35932
rect 6164 35876 6168 35932
rect 6104 35872 6168 35876
rect 6184 35932 6248 35936
rect 6184 35876 6188 35932
rect 6188 35876 6244 35932
rect 6244 35876 6248 35932
rect 6184 35872 6248 35876
rect 6264 35932 6328 35936
rect 6264 35876 6268 35932
rect 6268 35876 6324 35932
rect 6324 35876 6328 35932
rect 6264 35872 6328 35876
rect 6344 35932 6408 35936
rect 6344 35876 6348 35932
rect 6348 35876 6404 35932
rect 6404 35876 6408 35932
rect 6344 35872 6408 35876
rect 16407 35932 16471 35936
rect 16407 35876 16411 35932
rect 16411 35876 16467 35932
rect 16467 35876 16471 35932
rect 16407 35872 16471 35876
rect 16487 35932 16551 35936
rect 16487 35876 16491 35932
rect 16491 35876 16547 35932
rect 16547 35876 16551 35932
rect 16487 35872 16551 35876
rect 16567 35932 16631 35936
rect 16567 35876 16571 35932
rect 16571 35876 16627 35932
rect 16627 35876 16631 35932
rect 16567 35872 16631 35876
rect 16647 35932 16711 35936
rect 16647 35876 16651 35932
rect 16651 35876 16707 35932
rect 16707 35876 16711 35932
rect 16647 35872 16711 35876
rect 26711 35932 26775 35936
rect 26711 35876 26715 35932
rect 26715 35876 26771 35932
rect 26771 35876 26775 35932
rect 26711 35872 26775 35876
rect 26791 35932 26855 35936
rect 26791 35876 26795 35932
rect 26795 35876 26851 35932
rect 26851 35876 26855 35932
rect 26791 35872 26855 35876
rect 26871 35932 26935 35936
rect 26871 35876 26875 35932
rect 26875 35876 26931 35932
rect 26931 35876 26935 35932
rect 26871 35872 26935 35876
rect 26951 35932 27015 35936
rect 26951 35876 26955 35932
rect 26955 35876 27011 35932
rect 27011 35876 27015 35932
rect 26951 35872 27015 35876
rect 11255 35388 11319 35392
rect 11255 35332 11259 35388
rect 11259 35332 11315 35388
rect 11315 35332 11319 35388
rect 11255 35328 11319 35332
rect 11335 35388 11399 35392
rect 11335 35332 11339 35388
rect 11339 35332 11395 35388
rect 11395 35332 11399 35388
rect 11335 35328 11399 35332
rect 11415 35388 11479 35392
rect 11415 35332 11419 35388
rect 11419 35332 11475 35388
rect 11475 35332 11479 35388
rect 11415 35328 11479 35332
rect 11495 35388 11559 35392
rect 11495 35332 11499 35388
rect 11499 35332 11555 35388
rect 11555 35332 11559 35388
rect 11495 35328 11559 35332
rect 21559 35388 21623 35392
rect 21559 35332 21563 35388
rect 21563 35332 21619 35388
rect 21619 35332 21623 35388
rect 21559 35328 21623 35332
rect 21639 35388 21703 35392
rect 21639 35332 21643 35388
rect 21643 35332 21699 35388
rect 21699 35332 21703 35388
rect 21639 35328 21703 35332
rect 21719 35388 21783 35392
rect 21719 35332 21723 35388
rect 21723 35332 21779 35388
rect 21779 35332 21783 35388
rect 21719 35328 21783 35332
rect 21799 35388 21863 35392
rect 21799 35332 21803 35388
rect 21803 35332 21859 35388
rect 21859 35332 21863 35388
rect 21799 35328 21863 35332
rect 6104 34844 6168 34848
rect 6104 34788 6108 34844
rect 6108 34788 6164 34844
rect 6164 34788 6168 34844
rect 6104 34784 6168 34788
rect 6184 34844 6248 34848
rect 6184 34788 6188 34844
rect 6188 34788 6244 34844
rect 6244 34788 6248 34844
rect 6184 34784 6248 34788
rect 6264 34844 6328 34848
rect 6264 34788 6268 34844
rect 6268 34788 6324 34844
rect 6324 34788 6328 34844
rect 6264 34784 6328 34788
rect 6344 34844 6408 34848
rect 6344 34788 6348 34844
rect 6348 34788 6404 34844
rect 6404 34788 6408 34844
rect 6344 34784 6408 34788
rect 16407 34844 16471 34848
rect 16407 34788 16411 34844
rect 16411 34788 16467 34844
rect 16467 34788 16471 34844
rect 16407 34784 16471 34788
rect 16487 34844 16551 34848
rect 16487 34788 16491 34844
rect 16491 34788 16547 34844
rect 16547 34788 16551 34844
rect 16487 34784 16551 34788
rect 16567 34844 16631 34848
rect 16567 34788 16571 34844
rect 16571 34788 16627 34844
rect 16627 34788 16631 34844
rect 16567 34784 16631 34788
rect 16647 34844 16711 34848
rect 16647 34788 16651 34844
rect 16651 34788 16707 34844
rect 16707 34788 16711 34844
rect 16647 34784 16711 34788
rect 26711 34844 26775 34848
rect 26711 34788 26715 34844
rect 26715 34788 26771 34844
rect 26771 34788 26775 34844
rect 26711 34784 26775 34788
rect 26791 34844 26855 34848
rect 26791 34788 26795 34844
rect 26795 34788 26851 34844
rect 26851 34788 26855 34844
rect 26791 34784 26855 34788
rect 26871 34844 26935 34848
rect 26871 34788 26875 34844
rect 26875 34788 26931 34844
rect 26931 34788 26935 34844
rect 26871 34784 26935 34788
rect 26951 34844 27015 34848
rect 26951 34788 26955 34844
rect 26955 34788 27011 34844
rect 27011 34788 27015 34844
rect 26951 34784 27015 34788
rect 11255 34300 11319 34304
rect 11255 34244 11259 34300
rect 11259 34244 11315 34300
rect 11315 34244 11319 34300
rect 11255 34240 11319 34244
rect 11335 34300 11399 34304
rect 11335 34244 11339 34300
rect 11339 34244 11395 34300
rect 11395 34244 11399 34300
rect 11335 34240 11399 34244
rect 11415 34300 11479 34304
rect 11415 34244 11419 34300
rect 11419 34244 11475 34300
rect 11475 34244 11479 34300
rect 11415 34240 11479 34244
rect 11495 34300 11559 34304
rect 11495 34244 11499 34300
rect 11499 34244 11555 34300
rect 11555 34244 11559 34300
rect 11495 34240 11559 34244
rect 21559 34300 21623 34304
rect 21559 34244 21563 34300
rect 21563 34244 21619 34300
rect 21619 34244 21623 34300
rect 21559 34240 21623 34244
rect 21639 34300 21703 34304
rect 21639 34244 21643 34300
rect 21643 34244 21699 34300
rect 21699 34244 21703 34300
rect 21639 34240 21703 34244
rect 21719 34300 21783 34304
rect 21719 34244 21723 34300
rect 21723 34244 21779 34300
rect 21779 34244 21783 34300
rect 21719 34240 21783 34244
rect 21799 34300 21863 34304
rect 21799 34244 21803 34300
rect 21803 34244 21859 34300
rect 21859 34244 21863 34300
rect 21799 34240 21863 34244
rect 6104 33756 6168 33760
rect 6104 33700 6108 33756
rect 6108 33700 6164 33756
rect 6164 33700 6168 33756
rect 6104 33696 6168 33700
rect 6184 33756 6248 33760
rect 6184 33700 6188 33756
rect 6188 33700 6244 33756
rect 6244 33700 6248 33756
rect 6184 33696 6248 33700
rect 6264 33756 6328 33760
rect 6264 33700 6268 33756
rect 6268 33700 6324 33756
rect 6324 33700 6328 33756
rect 6264 33696 6328 33700
rect 6344 33756 6408 33760
rect 6344 33700 6348 33756
rect 6348 33700 6404 33756
rect 6404 33700 6408 33756
rect 6344 33696 6408 33700
rect 16407 33756 16471 33760
rect 16407 33700 16411 33756
rect 16411 33700 16467 33756
rect 16467 33700 16471 33756
rect 16407 33696 16471 33700
rect 16487 33756 16551 33760
rect 16487 33700 16491 33756
rect 16491 33700 16547 33756
rect 16547 33700 16551 33756
rect 16487 33696 16551 33700
rect 16567 33756 16631 33760
rect 16567 33700 16571 33756
rect 16571 33700 16627 33756
rect 16627 33700 16631 33756
rect 16567 33696 16631 33700
rect 16647 33756 16711 33760
rect 16647 33700 16651 33756
rect 16651 33700 16707 33756
rect 16707 33700 16711 33756
rect 16647 33696 16711 33700
rect 26711 33756 26775 33760
rect 26711 33700 26715 33756
rect 26715 33700 26771 33756
rect 26771 33700 26775 33756
rect 26711 33696 26775 33700
rect 26791 33756 26855 33760
rect 26791 33700 26795 33756
rect 26795 33700 26851 33756
rect 26851 33700 26855 33756
rect 26791 33696 26855 33700
rect 26871 33756 26935 33760
rect 26871 33700 26875 33756
rect 26875 33700 26931 33756
rect 26931 33700 26935 33756
rect 26871 33696 26935 33700
rect 26951 33756 27015 33760
rect 26951 33700 26955 33756
rect 26955 33700 27011 33756
rect 27011 33700 27015 33756
rect 26951 33696 27015 33700
rect 11255 33212 11319 33216
rect 11255 33156 11259 33212
rect 11259 33156 11315 33212
rect 11315 33156 11319 33212
rect 11255 33152 11319 33156
rect 11335 33212 11399 33216
rect 11335 33156 11339 33212
rect 11339 33156 11395 33212
rect 11395 33156 11399 33212
rect 11335 33152 11399 33156
rect 11415 33212 11479 33216
rect 11415 33156 11419 33212
rect 11419 33156 11475 33212
rect 11475 33156 11479 33212
rect 11415 33152 11479 33156
rect 11495 33212 11559 33216
rect 11495 33156 11499 33212
rect 11499 33156 11555 33212
rect 11555 33156 11559 33212
rect 11495 33152 11559 33156
rect 21559 33212 21623 33216
rect 21559 33156 21563 33212
rect 21563 33156 21619 33212
rect 21619 33156 21623 33212
rect 21559 33152 21623 33156
rect 21639 33212 21703 33216
rect 21639 33156 21643 33212
rect 21643 33156 21699 33212
rect 21699 33156 21703 33212
rect 21639 33152 21703 33156
rect 21719 33212 21783 33216
rect 21719 33156 21723 33212
rect 21723 33156 21779 33212
rect 21779 33156 21783 33212
rect 21719 33152 21783 33156
rect 21799 33212 21863 33216
rect 21799 33156 21803 33212
rect 21803 33156 21859 33212
rect 21859 33156 21863 33212
rect 21799 33152 21863 33156
rect 6104 32668 6168 32672
rect 6104 32612 6108 32668
rect 6108 32612 6164 32668
rect 6164 32612 6168 32668
rect 6104 32608 6168 32612
rect 6184 32668 6248 32672
rect 6184 32612 6188 32668
rect 6188 32612 6244 32668
rect 6244 32612 6248 32668
rect 6184 32608 6248 32612
rect 6264 32668 6328 32672
rect 6264 32612 6268 32668
rect 6268 32612 6324 32668
rect 6324 32612 6328 32668
rect 6264 32608 6328 32612
rect 6344 32668 6408 32672
rect 6344 32612 6348 32668
rect 6348 32612 6404 32668
rect 6404 32612 6408 32668
rect 6344 32608 6408 32612
rect 16407 32668 16471 32672
rect 16407 32612 16411 32668
rect 16411 32612 16467 32668
rect 16467 32612 16471 32668
rect 16407 32608 16471 32612
rect 16487 32668 16551 32672
rect 16487 32612 16491 32668
rect 16491 32612 16547 32668
rect 16547 32612 16551 32668
rect 16487 32608 16551 32612
rect 16567 32668 16631 32672
rect 16567 32612 16571 32668
rect 16571 32612 16627 32668
rect 16627 32612 16631 32668
rect 16567 32608 16631 32612
rect 16647 32668 16711 32672
rect 16647 32612 16651 32668
rect 16651 32612 16707 32668
rect 16707 32612 16711 32668
rect 16647 32608 16711 32612
rect 26711 32668 26775 32672
rect 26711 32612 26715 32668
rect 26715 32612 26771 32668
rect 26771 32612 26775 32668
rect 26711 32608 26775 32612
rect 26791 32668 26855 32672
rect 26791 32612 26795 32668
rect 26795 32612 26851 32668
rect 26851 32612 26855 32668
rect 26791 32608 26855 32612
rect 26871 32668 26935 32672
rect 26871 32612 26875 32668
rect 26875 32612 26931 32668
rect 26931 32612 26935 32668
rect 26871 32608 26935 32612
rect 26951 32668 27015 32672
rect 26951 32612 26955 32668
rect 26955 32612 27011 32668
rect 27011 32612 27015 32668
rect 26951 32608 27015 32612
rect 11255 32124 11319 32128
rect 11255 32068 11259 32124
rect 11259 32068 11315 32124
rect 11315 32068 11319 32124
rect 11255 32064 11319 32068
rect 11335 32124 11399 32128
rect 11335 32068 11339 32124
rect 11339 32068 11395 32124
rect 11395 32068 11399 32124
rect 11335 32064 11399 32068
rect 11415 32124 11479 32128
rect 11415 32068 11419 32124
rect 11419 32068 11475 32124
rect 11475 32068 11479 32124
rect 11415 32064 11479 32068
rect 11495 32124 11559 32128
rect 11495 32068 11499 32124
rect 11499 32068 11555 32124
rect 11555 32068 11559 32124
rect 11495 32064 11559 32068
rect 21559 32124 21623 32128
rect 21559 32068 21563 32124
rect 21563 32068 21619 32124
rect 21619 32068 21623 32124
rect 21559 32064 21623 32068
rect 21639 32124 21703 32128
rect 21639 32068 21643 32124
rect 21643 32068 21699 32124
rect 21699 32068 21703 32124
rect 21639 32064 21703 32068
rect 21719 32124 21783 32128
rect 21719 32068 21723 32124
rect 21723 32068 21779 32124
rect 21779 32068 21783 32124
rect 21719 32064 21783 32068
rect 21799 32124 21863 32128
rect 21799 32068 21803 32124
rect 21803 32068 21859 32124
rect 21859 32068 21863 32124
rect 21799 32064 21863 32068
rect 6104 31580 6168 31584
rect 6104 31524 6108 31580
rect 6108 31524 6164 31580
rect 6164 31524 6168 31580
rect 6104 31520 6168 31524
rect 6184 31580 6248 31584
rect 6184 31524 6188 31580
rect 6188 31524 6244 31580
rect 6244 31524 6248 31580
rect 6184 31520 6248 31524
rect 6264 31580 6328 31584
rect 6264 31524 6268 31580
rect 6268 31524 6324 31580
rect 6324 31524 6328 31580
rect 6264 31520 6328 31524
rect 6344 31580 6408 31584
rect 6344 31524 6348 31580
rect 6348 31524 6404 31580
rect 6404 31524 6408 31580
rect 6344 31520 6408 31524
rect 16407 31580 16471 31584
rect 16407 31524 16411 31580
rect 16411 31524 16467 31580
rect 16467 31524 16471 31580
rect 16407 31520 16471 31524
rect 16487 31580 16551 31584
rect 16487 31524 16491 31580
rect 16491 31524 16547 31580
rect 16547 31524 16551 31580
rect 16487 31520 16551 31524
rect 16567 31580 16631 31584
rect 16567 31524 16571 31580
rect 16571 31524 16627 31580
rect 16627 31524 16631 31580
rect 16567 31520 16631 31524
rect 16647 31580 16711 31584
rect 16647 31524 16651 31580
rect 16651 31524 16707 31580
rect 16707 31524 16711 31580
rect 16647 31520 16711 31524
rect 26711 31580 26775 31584
rect 26711 31524 26715 31580
rect 26715 31524 26771 31580
rect 26771 31524 26775 31580
rect 26711 31520 26775 31524
rect 26791 31580 26855 31584
rect 26791 31524 26795 31580
rect 26795 31524 26851 31580
rect 26851 31524 26855 31580
rect 26791 31520 26855 31524
rect 26871 31580 26935 31584
rect 26871 31524 26875 31580
rect 26875 31524 26931 31580
rect 26931 31524 26935 31580
rect 26871 31520 26935 31524
rect 26951 31580 27015 31584
rect 26951 31524 26955 31580
rect 26955 31524 27011 31580
rect 27011 31524 27015 31580
rect 26951 31520 27015 31524
rect 11255 31036 11319 31040
rect 11255 30980 11259 31036
rect 11259 30980 11315 31036
rect 11315 30980 11319 31036
rect 11255 30976 11319 30980
rect 11335 31036 11399 31040
rect 11335 30980 11339 31036
rect 11339 30980 11395 31036
rect 11395 30980 11399 31036
rect 11335 30976 11399 30980
rect 11415 31036 11479 31040
rect 11415 30980 11419 31036
rect 11419 30980 11475 31036
rect 11475 30980 11479 31036
rect 11415 30976 11479 30980
rect 11495 31036 11559 31040
rect 11495 30980 11499 31036
rect 11499 30980 11555 31036
rect 11555 30980 11559 31036
rect 11495 30976 11559 30980
rect 21559 31036 21623 31040
rect 21559 30980 21563 31036
rect 21563 30980 21619 31036
rect 21619 30980 21623 31036
rect 21559 30976 21623 30980
rect 21639 31036 21703 31040
rect 21639 30980 21643 31036
rect 21643 30980 21699 31036
rect 21699 30980 21703 31036
rect 21639 30976 21703 30980
rect 21719 31036 21783 31040
rect 21719 30980 21723 31036
rect 21723 30980 21779 31036
rect 21779 30980 21783 31036
rect 21719 30976 21783 30980
rect 21799 31036 21863 31040
rect 21799 30980 21803 31036
rect 21803 30980 21859 31036
rect 21859 30980 21863 31036
rect 21799 30976 21863 30980
rect 6104 30492 6168 30496
rect 6104 30436 6108 30492
rect 6108 30436 6164 30492
rect 6164 30436 6168 30492
rect 6104 30432 6168 30436
rect 6184 30492 6248 30496
rect 6184 30436 6188 30492
rect 6188 30436 6244 30492
rect 6244 30436 6248 30492
rect 6184 30432 6248 30436
rect 6264 30492 6328 30496
rect 6264 30436 6268 30492
rect 6268 30436 6324 30492
rect 6324 30436 6328 30492
rect 6264 30432 6328 30436
rect 6344 30492 6408 30496
rect 6344 30436 6348 30492
rect 6348 30436 6404 30492
rect 6404 30436 6408 30492
rect 6344 30432 6408 30436
rect 16407 30492 16471 30496
rect 16407 30436 16411 30492
rect 16411 30436 16467 30492
rect 16467 30436 16471 30492
rect 16407 30432 16471 30436
rect 16487 30492 16551 30496
rect 16487 30436 16491 30492
rect 16491 30436 16547 30492
rect 16547 30436 16551 30492
rect 16487 30432 16551 30436
rect 16567 30492 16631 30496
rect 16567 30436 16571 30492
rect 16571 30436 16627 30492
rect 16627 30436 16631 30492
rect 16567 30432 16631 30436
rect 16647 30492 16711 30496
rect 16647 30436 16651 30492
rect 16651 30436 16707 30492
rect 16707 30436 16711 30492
rect 16647 30432 16711 30436
rect 26711 30492 26775 30496
rect 26711 30436 26715 30492
rect 26715 30436 26771 30492
rect 26771 30436 26775 30492
rect 26711 30432 26775 30436
rect 26791 30492 26855 30496
rect 26791 30436 26795 30492
rect 26795 30436 26851 30492
rect 26851 30436 26855 30492
rect 26791 30432 26855 30436
rect 26871 30492 26935 30496
rect 26871 30436 26875 30492
rect 26875 30436 26931 30492
rect 26931 30436 26935 30492
rect 26871 30432 26935 30436
rect 26951 30492 27015 30496
rect 26951 30436 26955 30492
rect 26955 30436 27011 30492
rect 27011 30436 27015 30492
rect 26951 30432 27015 30436
rect 11255 29948 11319 29952
rect 11255 29892 11259 29948
rect 11259 29892 11315 29948
rect 11315 29892 11319 29948
rect 11255 29888 11319 29892
rect 11335 29948 11399 29952
rect 11335 29892 11339 29948
rect 11339 29892 11395 29948
rect 11395 29892 11399 29948
rect 11335 29888 11399 29892
rect 11415 29948 11479 29952
rect 11415 29892 11419 29948
rect 11419 29892 11475 29948
rect 11475 29892 11479 29948
rect 11415 29888 11479 29892
rect 11495 29948 11559 29952
rect 11495 29892 11499 29948
rect 11499 29892 11555 29948
rect 11555 29892 11559 29948
rect 11495 29888 11559 29892
rect 21559 29948 21623 29952
rect 21559 29892 21563 29948
rect 21563 29892 21619 29948
rect 21619 29892 21623 29948
rect 21559 29888 21623 29892
rect 21639 29948 21703 29952
rect 21639 29892 21643 29948
rect 21643 29892 21699 29948
rect 21699 29892 21703 29948
rect 21639 29888 21703 29892
rect 21719 29948 21783 29952
rect 21719 29892 21723 29948
rect 21723 29892 21779 29948
rect 21779 29892 21783 29948
rect 21719 29888 21783 29892
rect 21799 29948 21863 29952
rect 21799 29892 21803 29948
rect 21803 29892 21859 29948
rect 21859 29892 21863 29948
rect 21799 29888 21863 29892
rect 6104 29404 6168 29408
rect 6104 29348 6108 29404
rect 6108 29348 6164 29404
rect 6164 29348 6168 29404
rect 6104 29344 6168 29348
rect 6184 29404 6248 29408
rect 6184 29348 6188 29404
rect 6188 29348 6244 29404
rect 6244 29348 6248 29404
rect 6184 29344 6248 29348
rect 6264 29404 6328 29408
rect 6264 29348 6268 29404
rect 6268 29348 6324 29404
rect 6324 29348 6328 29404
rect 6264 29344 6328 29348
rect 6344 29404 6408 29408
rect 6344 29348 6348 29404
rect 6348 29348 6404 29404
rect 6404 29348 6408 29404
rect 6344 29344 6408 29348
rect 16407 29404 16471 29408
rect 16407 29348 16411 29404
rect 16411 29348 16467 29404
rect 16467 29348 16471 29404
rect 16407 29344 16471 29348
rect 16487 29404 16551 29408
rect 16487 29348 16491 29404
rect 16491 29348 16547 29404
rect 16547 29348 16551 29404
rect 16487 29344 16551 29348
rect 16567 29404 16631 29408
rect 16567 29348 16571 29404
rect 16571 29348 16627 29404
rect 16627 29348 16631 29404
rect 16567 29344 16631 29348
rect 16647 29404 16711 29408
rect 16647 29348 16651 29404
rect 16651 29348 16707 29404
rect 16707 29348 16711 29404
rect 16647 29344 16711 29348
rect 26711 29404 26775 29408
rect 26711 29348 26715 29404
rect 26715 29348 26771 29404
rect 26771 29348 26775 29404
rect 26711 29344 26775 29348
rect 26791 29404 26855 29408
rect 26791 29348 26795 29404
rect 26795 29348 26851 29404
rect 26851 29348 26855 29404
rect 26791 29344 26855 29348
rect 26871 29404 26935 29408
rect 26871 29348 26875 29404
rect 26875 29348 26931 29404
rect 26931 29348 26935 29404
rect 26871 29344 26935 29348
rect 26951 29404 27015 29408
rect 26951 29348 26955 29404
rect 26955 29348 27011 29404
rect 27011 29348 27015 29404
rect 26951 29344 27015 29348
rect 11255 28860 11319 28864
rect 11255 28804 11259 28860
rect 11259 28804 11315 28860
rect 11315 28804 11319 28860
rect 11255 28800 11319 28804
rect 11335 28860 11399 28864
rect 11335 28804 11339 28860
rect 11339 28804 11395 28860
rect 11395 28804 11399 28860
rect 11335 28800 11399 28804
rect 11415 28860 11479 28864
rect 11415 28804 11419 28860
rect 11419 28804 11475 28860
rect 11475 28804 11479 28860
rect 11415 28800 11479 28804
rect 11495 28860 11559 28864
rect 11495 28804 11499 28860
rect 11499 28804 11555 28860
rect 11555 28804 11559 28860
rect 11495 28800 11559 28804
rect 21559 28860 21623 28864
rect 21559 28804 21563 28860
rect 21563 28804 21619 28860
rect 21619 28804 21623 28860
rect 21559 28800 21623 28804
rect 21639 28860 21703 28864
rect 21639 28804 21643 28860
rect 21643 28804 21699 28860
rect 21699 28804 21703 28860
rect 21639 28800 21703 28804
rect 21719 28860 21783 28864
rect 21719 28804 21723 28860
rect 21723 28804 21779 28860
rect 21779 28804 21783 28860
rect 21719 28800 21783 28804
rect 21799 28860 21863 28864
rect 21799 28804 21803 28860
rect 21803 28804 21859 28860
rect 21859 28804 21863 28860
rect 21799 28800 21863 28804
rect 6104 28316 6168 28320
rect 6104 28260 6108 28316
rect 6108 28260 6164 28316
rect 6164 28260 6168 28316
rect 6104 28256 6168 28260
rect 6184 28316 6248 28320
rect 6184 28260 6188 28316
rect 6188 28260 6244 28316
rect 6244 28260 6248 28316
rect 6184 28256 6248 28260
rect 6264 28316 6328 28320
rect 6264 28260 6268 28316
rect 6268 28260 6324 28316
rect 6324 28260 6328 28316
rect 6264 28256 6328 28260
rect 6344 28316 6408 28320
rect 6344 28260 6348 28316
rect 6348 28260 6404 28316
rect 6404 28260 6408 28316
rect 6344 28256 6408 28260
rect 16407 28316 16471 28320
rect 16407 28260 16411 28316
rect 16411 28260 16467 28316
rect 16467 28260 16471 28316
rect 16407 28256 16471 28260
rect 16487 28316 16551 28320
rect 16487 28260 16491 28316
rect 16491 28260 16547 28316
rect 16547 28260 16551 28316
rect 16487 28256 16551 28260
rect 16567 28316 16631 28320
rect 16567 28260 16571 28316
rect 16571 28260 16627 28316
rect 16627 28260 16631 28316
rect 16567 28256 16631 28260
rect 16647 28316 16711 28320
rect 16647 28260 16651 28316
rect 16651 28260 16707 28316
rect 16707 28260 16711 28316
rect 16647 28256 16711 28260
rect 26711 28316 26775 28320
rect 26711 28260 26715 28316
rect 26715 28260 26771 28316
rect 26771 28260 26775 28316
rect 26711 28256 26775 28260
rect 26791 28316 26855 28320
rect 26791 28260 26795 28316
rect 26795 28260 26851 28316
rect 26851 28260 26855 28316
rect 26791 28256 26855 28260
rect 26871 28316 26935 28320
rect 26871 28260 26875 28316
rect 26875 28260 26931 28316
rect 26931 28260 26935 28316
rect 26871 28256 26935 28260
rect 26951 28316 27015 28320
rect 26951 28260 26955 28316
rect 26955 28260 27011 28316
rect 27011 28260 27015 28316
rect 26951 28256 27015 28260
rect 11255 27772 11319 27776
rect 11255 27716 11259 27772
rect 11259 27716 11315 27772
rect 11315 27716 11319 27772
rect 11255 27712 11319 27716
rect 11335 27772 11399 27776
rect 11335 27716 11339 27772
rect 11339 27716 11395 27772
rect 11395 27716 11399 27772
rect 11335 27712 11399 27716
rect 11415 27772 11479 27776
rect 11415 27716 11419 27772
rect 11419 27716 11475 27772
rect 11475 27716 11479 27772
rect 11415 27712 11479 27716
rect 11495 27772 11559 27776
rect 11495 27716 11499 27772
rect 11499 27716 11555 27772
rect 11555 27716 11559 27772
rect 11495 27712 11559 27716
rect 21559 27772 21623 27776
rect 21559 27716 21563 27772
rect 21563 27716 21619 27772
rect 21619 27716 21623 27772
rect 21559 27712 21623 27716
rect 21639 27772 21703 27776
rect 21639 27716 21643 27772
rect 21643 27716 21699 27772
rect 21699 27716 21703 27772
rect 21639 27712 21703 27716
rect 21719 27772 21783 27776
rect 21719 27716 21723 27772
rect 21723 27716 21779 27772
rect 21779 27716 21783 27772
rect 21719 27712 21783 27716
rect 21799 27772 21863 27776
rect 21799 27716 21803 27772
rect 21803 27716 21859 27772
rect 21859 27716 21863 27772
rect 21799 27712 21863 27716
rect 6104 27228 6168 27232
rect 6104 27172 6108 27228
rect 6108 27172 6164 27228
rect 6164 27172 6168 27228
rect 6104 27168 6168 27172
rect 6184 27228 6248 27232
rect 6184 27172 6188 27228
rect 6188 27172 6244 27228
rect 6244 27172 6248 27228
rect 6184 27168 6248 27172
rect 6264 27228 6328 27232
rect 6264 27172 6268 27228
rect 6268 27172 6324 27228
rect 6324 27172 6328 27228
rect 6264 27168 6328 27172
rect 6344 27228 6408 27232
rect 6344 27172 6348 27228
rect 6348 27172 6404 27228
rect 6404 27172 6408 27228
rect 6344 27168 6408 27172
rect 16407 27228 16471 27232
rect 16407 27172 16411 27228
rect 16411 27172 16467 27228
rect 16467 27172 16471 27228
rect 16407 27168 16471 27172
rect 16487 27228 16551 27232
rect 16487 27172 16491 27228
rect 16491 27172 16547 27228
rect 16547 27172 16551 27228
rect 16487 27168 16551 27172
rect 16567 27228 16631 27232
rect 16567 27172 16571 27228
rect 16571 27172 16627 27228
rect 16627 27172 16631 27228
rect 16567 27168 16631 27172
rect 16647 27228 16711 27232
rect 16647 27172 16651 27228
rect 16651 27172 16707 27228
rect 16707 27172 16711 27228
rect 16647 27168 16711 27172
rect 26711 27228 26775 27232
rect 26711 27172 26715 27228
rect 26715 27172 26771 27228
rect 26771 27172 26775 27228
rect 26711 27168 26775 27172
rect 26791 27228 26855 27232
rect 26791 27172 26795 27228
rect 26795 27172 26851 27228
rect 26851 27172 26855 27228
rect 26791 27168 26855 27172
rect 26871 27228 26935 27232
rect 26871 27172 26875 27228
rect 26875 27172 26931 27228
rect 26931 27172 26935 27228
rect 26871 27168 26935 27172
rect 26951 27228 27015 27232
rect 26951 27172 26955 27228
rect 26955 27172 27011 27228
rect 27011 27172 27015 27228
rect 26951 27168 27015 27172
rect 11255 26684 11319 26688
rect 11255 26628 11259 26684
rect 11259 26628 11315 26684
rect 11315 26628 11319 26684
rect 11255 26624 11319 26628
rect 11335 26684 11399 26688
rect 11335 26628 11339 26684
rect 11339 26628 11395 26684
rect 11395 26628 11399 26684
rect 11335 26624 11399 26628
rect 11415 26684 11479 26688
rect 11415 26628 11419 26684
rect 11419 26628 11475 26684
rect 11475 26628 11479 26684
rect 11415 26624 11479 26628
rect 11495 26684 11559 26688
rect 11495 26628 11499 26684
rect 11499 26628 11555 26684
rect 11555 26628 11559 26684
rect 11495 26624 11559 26628
rect 21559 26684 21623 26688
rect 21559 26628 21563 26684
rect 21563 26628 21619 26684
rect 21619 26628 21623 26684
rect 21559 26624 21623 26628
rect 21639 26684 21703 26688
rect 21639 26628 21643 26684
rect 21643 26628 21699 26684
rect 21699 26628 21703 26684
rect 21639 26624 21703 26628
rect 21719 26684 21783 26688
rect 21719 26628 21723 26684
rect 21723 26628 21779 26684
rect 21779 26628 21783 26684
rect 21719 26624 21783 26628
rect 21799 26684 21863 26688
rect 21799 26628 21803 26684
rect 21803 26628 21859 26684
rect 21859 26628 21863 26684
rect 21799 26624 21863 26628
rect 6104 26140 6168 26144
rect 6104 26084 6108 26140
rect 6108 26084 6164 26140
rect 6164 26084 6168 26140
rect 6104 26080 6168 26084
rect 6184 26140 6248 26144
rect 6184 26084 6188 26140
rect 6188 26084 6244 26140
rect 6244 26084 6248 26140
rect 6184 26080 6248 26084
rect 6264 26140 6328 26144
rect 6264 26084 6268 26140
rect 6268 26084 6324 26140
rect 6324 26084 6328 26140
rect 6264 26080 6328 26084
rect 6344 26140 6408 26144
rect 6344 26084 6348 26140
rect 6348 26084 6404 26140
rect 6404 26084 6408 26140
rect 6344 26080 6408 26084
rect 16407 26140 16471 26144
rect 16407 26084 16411 26140
rect 16411 26084 16467 26140
rect 16467 26084 16471 26140
rect 16407 26080 16471 26084
rect 16487 26140 16551 26144
rect 16487 26084 16491 26140
rect 16491 26084 16547 26140
rect 16547 26084 16551 26140
rect 16487 26080 16551 26084
rect 16567 26140 16631 26144
rect 16567 26084 16571 26140
rect 16571 26084 16627 26140
rect 16627 26084 16631 26140
rect 16567 26080 16631 26084
rect 16647 26140 16711 26144
rect 16647 26084 16651 26140
rect 16651 26084 16707 26140
rect 16707 26084 16711 26140
rect 16647 26080 16711 26084
rect 26711 26140 26775 26144
rect 26711 26084 26715 26140
rect 26715 26084 26771 26140
rect 26771 26084 26775 26140
rect 26711 26080 26775 26084
rect 26791 26140 26855 26144
rect 26791 26084 26795 26140
rect 26795 26084 26851 26140
rect 26851 26084 26855 26140
rect 26791 26080 26855 26084
rect 26871 26140 26935 26144
rect 26871 26084 26875 26140
rect 26875 26084 26931 26140
rect 26931 26084 26935 26140
rect 26871 26080 26935 26084
rect 26951 26140 27015 26144
rect 26951 26084 26955 26140
rect 26955 26084 27011 26140
rect 27011 26084 27015 26140
rect 26951 26080 27015 26084
rect 11255 25596 11319 25600
rect 11255 25540 11259 25596
rect 11259 25540 11315 25596
rect 11315 25540 11319 25596
rect 11255 25536 11319 25540
rect 11335 25596 11399 25600
rect 11335 25540 11339 25596
rect 11339 25540 11395 25596
rect 11395 25540 11399 25596
rect 11335 25536 11399 25540
rect 11415 25596 11479 25600
rect 11415 25540 11419 25596
rect 11419 25540 11475 25596
rect 11475 25540 11479 25596
rect 11415 25536 11479 25540
rect 11495 25596 11559 25600
rect 11495 25540 11499 25596
rect 11499 25540 11555 25596
rect 11555 25540 11559 25596
rect 11495 25536 11559 25540
rect 21559 25596 21623 25600
rect 21559 25540 21563 25596
rect 21563 25540 21619 25596
rect 21619 25540 21623 25596
rect 21559 25536 21623 25540
rect 21639 25596 21703 25600
rect 21639 25540 21643 25596
rect 21643 25540 21699 25596
rect 21699 25540 21703 25596
rect 21639 25536 21703 25540
rect 21719 25596 21783 25600
rect 21719 25540 21723 25596
rect 21723 25540 21779 25596
rect 21779 25540 21783 25596
rect 21719 25536 21783 25540
rect 21799 25596 21863 25600
rect 21799 25540 21803 25596
rect 21803 25540 21859 25596
rect 21859 25540 21863 25596
rect 21799 25536 21863 25540
rect 6104 25052 6168 25056
rect 6104 24996 6108 25052
rect 6108 24996 6164 25052
rect 6164 24996 6168 25052
rect 6104 24992 6168 24996
rect 6184 25052 6248 25056
rect 6184 24996 6188 25052
rect 6188 24996 6244 25052
rect 6244 24996 6248 25052
rect 6184 24992 6248 24996
rect 6264 25052 6328 25056
rect 6264 24996 6268 25052
rect 6268 24996 6324 25052
rect 6324 24996 6328 25052
rect 6264 24992 6328 24996
rect 6344 25052 6408 25056
rect 6344 24996 6348 25052
rect 6348 24996 6404 25052
rect 6404 24996 6408 25052
rect 6344 24992 6408 24996
rect 16407 25052 16471 25056
rect 16407 24996 16411 25052
rect 16411 24996 16467 25052
rect 16467 24996 16471 25052
rect 16407 24992 16471 24996
rect 16487 25052 16551 25056
rect 16487 24996 16491 25052
rect 16491 24996 16547 25052
rect 16547 24996 16551 25052
rect 16487 24992 16551 24996
rect 16567 25052 16631 25056
rect 16567 24996 16571 25052
rect 16571 24996 16627 25052
rect 16627 24996 16631 25052
rect 16567 24992 16631 24996
rect 16647 25052 16711 25056
rect 16647 24996 16651 25052
rect 16651 24996 16707 25052
rect 16707 24996 16711 25052
rect 16647 24992 16711 24996
rect 26711 25052 26775 25056
rect 26711 24996 26715 25052
rect 26715 24996 26771 25052
rect 26771 24996 26775 25052
rect 26711 24992 26775 24996
rect 26791 25052 26855 25056
rect 26791 24996 26795 25052
rect 26795 24996 26851 25052
rect 26851 24996 26855 25052
rect 26791 24992 26855 24996
rect 26871 25052 26935 25056
rect 26871 24996 26875 25052
rect 26875 24996 26931 25052
rect 26931 24996 26935 25052
rect 26871 24992 26935 24996
rect 26951 25052 27015 25056
rect 26951 24996 26955 25052
rect 26955 24996 27011 25052
rect 27011 24996 27015 25052
rect 26951 24992 27015 24996
rect 11255 24508 11319 24512
rect 11255 24452 11259 24508
rect 11259 24452 11315 24508
rect 11315 24452 11319 24508
rect 11255 24448 11319 24452
rect 11335 24508 11399 24512
rect 11335 24452 11339 24508
rect 11339 24452 11395 24508
rect 11395 24452 11399 24508
rect 11335 24448 11399 24452
rect 11415 24508 11479 24512
rect 11415 24452 11419 24508
rect 11419 24452 11475 24508
rect 11475 24452 11479 24508
rect 11415 24448 11479 24452
rect 11495 24508 11559 24512
rect 11495 24452 11499 24508
rect 11499 24452 11555 24508
rect 11555 24452 11559 24508
rect 11495 24448 11559 24452
rect 21559 24508 21623 24512
rect 21559 24452 21563 24508
rect 21563 24452 21619 24508
rect 21619 24452 21623 24508
rect 21559 24448 21623 24452
rect 21639 24508 21703 24512
rect 21639 24452 21643 24508
rect 21643 24452 21699 24508
rect 21699 24452 21703 24508
rect 21639 24448 21703 24452
rect 21719 24508 21783 24512
rect 21719 24452 21723 24508
rect 21723 24452 21779 24508
rect 21779 24452 21783 24508
rect 21719 24448 21783 24452
rect 21799 24508 21863 24512
rect 21799 24452 21803 24508
rect 21803 24452 21859 24508
rect 21859 24452 21863 24508
rect 21799 24448 21863 24452
rect 6104 23964 6168 23968
rect 6104 23908 6108 23964
rect 6108 23908 6164 23964
rect 6164 23908 6168 23964
rect 6104 23904 6168 23908
rect 6184 23964 6248 23968
rect 6184 23908 6188 23964
rect 6188 23908 6244 23964
rect 6244 23908 6248 23964
rect 6184 23904 6248 23908
rect 6264 23964 6328 23968
rect 6264 23908 6268 23964
rect 6268 23908 6324 23964
rect 6324 23908 6328 23964
rect 6264 23904 6328 23908
rect 6344 23964 6408 23968
rect 6344 23908 6348 23964
rect 6348 23908 6404 23964
rect 6404 23908 6408 23964
rect 6344 23904 6408 23908
rect 16407 23964 16471 23968
rect 16407 23908 16411 23964
rect 16411 23908 16467 23964
rect 16467 23908 16471 23964
rect 16407 23904 16471 23908
rect 16487 23964 16551 23968
rect 16487 23908 16491 23964
rect 16491 23908 16547 23964
rect 16547 23908 16551 23964
rect 16487 23904 16551 23908
rect 16567 23964 16631 23968
rect 16567 23908 16571 23964
rect 16571 23908 16627 23964
rect 16627 23908 16631 23964
rect 16567 23904 16631 23908
rect 16647 23964 16711 23968
rect 16647 23908 16651 23964
rect 16651 23908 16707 23964
rect 16707 23908 16711 23964
rect 16647 23904 16711 23908
rect 26711 23964 26775 23968
rect 26711 23908 26715 23964
rect 26715 23908 26771 23964
rect 26771 23908 26775 23964
rect 26711 23904 26775 23908
rect 26791 23964 26855 23968
rect 26791 23908 26795 23964
rect 26795 23908 26851 23964
rect 26851 23908 26855 23964
rect 26791 23904 26855 23908
rect 26871 23964 26935 23968
rect 26871 23908 26875 23964
rect 26875 23908 26931 23964
rect 26931 23908 26935 23964
rect 26871 23904 26935 23908
rect 26951 23964 27015 23968
rect 26951 23908 26955 23964
rect 26955 23908 27011 23964
rect 27011 23908 27015 23964
rect 26951 23904 27015 23908
rect 11255 23420 11319 23424
rect 11255 23364 11259 23420
rect 11259 23364 11315 23420
rect 11315 23364 11319 23420
rect 11255 23360 11319 23364
rect 11335 23420 11399 23424
rect 11335 23364 11339 23420
rect 11339 23364 11395 23420
rect 11395 23364 11399 23420
rect 11335 23360 11399 23364
rect 11415 23420 11479 23424
rect 11415 23364 11419 23420
rect 11419 23364 11475 23420
rect 11475 23364 11479 23420
rect 11415 23360 11479 23364
rect 11495 23420 11559 23424
rect 11495 23364 11499 23420
rect 11499 23364 11555 23420
rect 11555 23364 11559 23420
rect 11495 23360 11559 23364
rect 21559 23420 21623 23424
rect 21559 23364 21563 23420
rect 21563 23364 21619 23420
rect 21619 23364 21623 23420
rect 21559 23360 21623 23364
rect 21639 23420 21703 23424
rect 21639 23364 21643 23420
rect 21643 23364 21699 23420
rect 21699 23364 21703 23420
rect 21639 23360 21703 23364
rect 21719 23420 21783 23424
rect 21719 23364 21723 23420
rect 21723 23364 21779 23420
rect 21779 23364 21783 23420
rect 21719 23360 21783 23364
rect 21799 23420 21863 23424
rect 21799 23364 21803 23420
rect 21803 23364 21859 23420
rect 21859 23364 21863 23420
rect 21799 23360 21863 23364
rect 6104 22876 6168 22880
rect 6104 22820 6108 22876
rect 6108 22820 6164 22876
rect 6164 22820 6168 22876
rect 6104 22816 6168 22820
rect 6184 22876 6248 22880
rect 6184 22820 6188 22876
rect 6188 22820 6244 22876
rect 6244 22820 6248 22876
rect 6184 22816 6248 22820
rect 6264 22876 6328 22880
rect 6264 22820 6268 22876
rect 6268 22820 6324 22876
rect 6324 22820 6328 22876
rect 6264 22816 6328 22820
rect 6344 22876 6408 22880
rect 6344 22820 6348 22876
rect 6348 22820 6404 22876
rect 6404 22820 6408 22876
rect 6344 22816 6408 22820
rect 16407 22876 16471 22880
rect 16407 22820 16411 22876
rect 16411 22820 16467 22876
rect 16467 22820 16471 22876
rect 16407 22816 16471 22820
rect 16487 22876 16551 22880
rect 16487 22820 16491 22876
rect 16491 22820 16547 22876
rect 16547 22820 16551 22876
rect 16487 22816 16551 22820
rect 16567 22876 16631 22880
rect 16567 22820 16571 22876
rect 16571 22820 16627 22876
rect 16627 22820 16631 22876
rect 16567 22816 16631 22820
rect 16647 22876 16711 22880
rect 16647 22820 16651 22876
rect 16651 22820 16707 22876
rect 16707 22820 16711 22876
rect 16647 22816 16711 22820
rect 26711 22876 26775 22880
rect 26711 22820 26715 22876
rect 26715 22820 26771 22876
rect 26771 22820 26775 22876
rect 26711 22816 26775 22820
rect 26791 22876 26855 22880
rect 26791 22820 26795 22876
rect 26795 22820 26851 22876
rect 26851 22820 26855 22876
rect 26791 22816 26855 22820
rect 26871 22876 26935 22880
rect 26871 22820 26875 22876
rect 26875 22820 26931 22876
rect 26931 22820 26935 22876
rect 26871 22816 26935 22820
rect 26951 22876 27015 22880
rect 26951 22820 26955 22876
rect 26955 22820 27011 22876
rect 27011 22820 27015 22876
rect 26951 22816 27015 22820
rect 11255 22332 11319 22336
rect 11255 22276 11259 22332
rect 11259 22276 11315 22332
rect 11315 22276 11319 22332
rect 11255 22272 11319 22276
rect 11335 22332 11399 22336
rect 11335 22276 11339 22332
rect 11339 22276 11395 22332
rect 11395 22276 11399 22332
rect 11335 22272 11399 22276
rect 11415 22332 11479 22336
rect 11415 22276 11419 22332
rect 11419 22276 11475 22332
rect 11475 22276 11479 22332
rect 11415 22272 11479 22276
rect 11495 22332 11559 22336
rect 11495 22276 11499 22332
rect 11499 22276 11555 22332
rect 11555 22276 11559 22332
rect 11495 22272 11559 22276
rect 21559 22332 21623 22336
rect 21559 22276 21563 22332
rect 21563 22276 21619 22332
rect 21619 22276 21623 22332
rect 21559 22272 21623 22276
rect 21639 22332 21703 22336
rect 21639 22276 21643 22332
rect 21643 22276 21699 22332
rect 21699 22276 21703 22332
rect 21639 22272 21703 22276
rect 21719 22332 21783 22336
rect 21719 22276 21723 22332
rect 21723 22276 21779 22332
rect 21779 22276 21783 22332
rect 21719 22272 21783 22276
rect 21799 22332 21863 22336
rect 21799 22276 21803 22332
rect 21803 22276 21859 22332
rect 21859 22276 21863 22332
rect 21799 22272 21863 22276
rect 6104 21788 6168 21792
rect 6104 21732 6108 21788
rect 6108 21732 6164 21788
rect 6164 21732 6168 21788
rect 6104 21728 6168 21732
rect 6184 21788 6248 21792
rect 6184 21732 6188 21788
rect 6188 21732 6244 21788
rect 6244 21732 6248 21788
rect 6184 21728 6248 21732
rect 6264 21788 6328 21792
rect 6264 21732 6268 21788
rect 6268 21732 6324 21788
rect 6324 21732 6328 21788
rect 6264 21728 6328 21732
rect 6344 21788 6408 21792
rect 6344 21732 6348 21788
rect 6348 21732 6404 21788
rect 6404 21732 6408 21788
rect 6344 21728 6408 21732
rect 16407 21788 16471 21792
rect 16407 21732 16411 21788
rect 16411 21732 16467 21788
rect 16467 21732 16471 21788
rect 16407 21728 16471 21732
rect 16487 21788 16551 21792
rect 16487 21732 16491 21788
rect 16491 21732 16547 21788
rect 16547 21732 16551 21788
rect 16487 21728 16551 21732
rect 16567 21788 16631 21792
rect 16567 21732 16571 21788
rect 16571 21732 16627 21788
rect 16627 21732 16631 21788
rect 16567 21728 16631 21732
rect 16647 21788 16711 21792
rect 16647 21732 16651 21788
rect 16651 21732 16707 21788
rect 16707 21732 16711 21788
rect 16647 21728 16711 21732
rect 26711 21788 26775 21792
rect 26711 21732 26715 21788
rect 26715 21732 26771 21788
rect 26771 21732 26775 21788
rect 26711 21728 26775 21732
rect 26791 21788 26855 21792
rect 26791 21732 26795 21788
rect 26795 21732 26851 21788
rect 26851 21732 26855 21788
rect 26791 21728 26855 21732
rect 26871 21788 26935 21792
rect 26871 21732 26875 21788
rect 26875 21732 26931 21788
rect 26931 21732 26935 21788
rect 26871 21728 26935 21732
rect 26951 21788 27015 21792
rect 26951 21732 26955 21788
rect 26955 21732 27011 21788
rect 27011 21732 27015 21788
rect 26951 21728 27015 21732
rect 11255 21244 11319 21248
rect 11255 21188 11259 21244
rect 11259 21188 11315 21244
rect 11315 21188 11319 21244
rect 11255 21184 11319 21188
rect 11335 21244 11399 21248
rect 11335 21188 11339 21244
rect 11339 21188 11395 21244
rect 11395 21188 11399 21244
rect 11335 21184 11399 21188
rect 11415 21244 11479 21248
rect 11415 21188 11419 21244
rect 11419 21188 11475 21244
rect 11475 21188 11479 21244
rect 11415 21184 11479 21188
rect 11495 21244 11559 21248
rect 11495 21188 11499 21244
rect 11499 21188 11555 21244
rect 11555 21188 11559 21244
rect 11495 21184 11559 21188
rect 21559 21244 21623 21248
rect 21559 21188 21563 21244
rect 21563 21188 21619 21244
rect 21619 21188 21623 21244
rect 21559 21184 21623 21188
rect 21639 21244 21703 21248
rect 21639 21188 21643 21244
rect 21643 21188 21699 21244
rect 21699 21188 21703 21244
rect 21639 21184 21703 21188
rect 21719 21244 21783 21248
rect 21719 21188 21723 21244
rect 21723 21188 21779 21244
rect 21779 21188 21783 21244
rect 21719 21184 21783 21188
rect 21799 21244 21863 21248
rect 21799 21188 21803 21244
rect 21803 21188 21859 21244
rect 21859 21188 21863 21244
rect 21799 21184 21863 21188
rect 6104 20700 6168 20704
rect 6104 20644 6108 20700
rect 6108 20644 6164 20700
rect 6164 20644 6168 20700
rect 6104 20640 6168 20644
rect 6184 20700 6248 20704
rect 6184 20644 6188 20700
rect 6188 20644 6244 20700
rect 6244 20644 6248 20700
rect 6184 20640 6248 20644
rect 6264 20700 6328 20704
rect 6264 20644 6268 20700
rect 6268 20644 6324 20700
rect 6324 20644 6328 20700
rect 6264 20640 6328 20644
rect 6344 20700 6408 20704
rect 6344 20644 6348 20700
rect 6348 20644 6404 20700
rect 6404 20644 6408 20700
rect 6344 20640 6408 20644
rect 16407 20700 16471 20704
rect 16407 20644 16411 20700
rect 16411 20644 16467 20700
rect 16467 20644 16471 20700
rect 16407 20640 16471 20644
rect 16487 20700 16551 20704
rect 16487 20644 16491 20700
rect 16491 20644 16547 20700
rect 16547 20644 16551 20700
rect 16487 20640 16551 20644
rect 16567 20700 16631 20704
rect 16567 20644 16571 20700
rect 16571 20644 16627 20700
rect 16627 20644 16631 20700
rect 16567 20640 16631 20644
rect 16647 20700 16711 20704
rect 16647 20644 16651 20700
rect 16651 20644 16707 20700
rect 16707 20644 16711 20700
rect 16647 20640 16711 20644
rect 26711 20700 26775 20704
rect 26711 20644 26715 20700
rect 26715 20644 26771 20700
rect 26771 20644 26775 20700
rect 26711 20640 26775 20644
rect 26791 20700 26855 20704
rect 26791 20644 26795 20700
rect 26795 20644 26851 20700
rect 26851 20644 26855 20700
rect 26791 20640 26855 20644
rect 26871 20700 26935 20704
rect 26871 20644 26875 20700
rect 26875 20644 26931 20700
rect 26931 20644 26935 20700
rect 26871 20640 26935 20644
rect 26951 20700 27015 20704
rect 26951 20644 26955 20700
rect 26955 20644 27011 20700
rect 27011 20644 27015 20700
rect 26951 20640 27015 20644
rect 11255 20156 11319 20160
rect 11255 20100 11259 20156
rect 11259 20100 11315 20156
rect 11315 20100 11319 20156
rect 11255 20096 11319 20100
rect 11335 20156 11399 20160
rect 11335 20100 11339 20156
rect 11339 20100 11395 20156
rect 11395 20100 11399 20156
rect 11335 20096 11399 20100
rect 11415 20156 11479 20160
rect 11415 20100 11419 20156
rect 11419 20100 11475 20156
rect 11475 20100 11479 20156
rect 11415 20096 11479 20100
rect 11495 20156 11559 20160
rect 11495 20100 11499 20156
rect 11499 20100 11555 20156
rect 11555 20100 11559 20156
rect 11495 20096 11559 20100
rect 21559 20156 21623 20160
rect 21559 20100 21563 20156
rect 21563 20100 21619 20156
rect 21619 20100 21623 20156
rect 21559 20096 21623 20100
rect 21639 20156 21703 20160
rect 21639 20100 21643 20156
rect 21643 20100 21699 20156
rect 21699 20100 21703 20156
rect 21639 20096 21703 20100
rect 21719 20156 21783 20160
rect 21719 20100 21723 20156
rect 21723 20100 21779 20156
rect 21779 20100 21783 20156
rect 21719 20096 21783 20100
rect 21799 20156 21863 20160
rect 21799 20100 21803 20156
rect 21803 20100 21859 20156
rect 21859 20100 21863 20156
rect 21799 20096 21863 20100
rect 6104 19612 6168 19616
rect 6104 19556 6108 19612
rect 6108 19556 6164 19612
rect 6164 19556 6168 19612
rect 6104 19552 6168 19556
rect 6184 19612 6248 19616
rect 6184 19556 6188 19612
rect 6188 19556 6244 19612
rect 6244 19556 6248 19612
rect 6184 19552 6248 19556
rect 6264 19612 6328 19616
rect 6264 19556 6268 19612
rect 6268 19556 6324 19612
rect 6324 19556 6328 19612
rect 6264 19552 6328 19556
rect 6344 19612 6408 19616
rect 6344 19556 6348 19612
rect 6348 19556 6404 19612
rect 6404 19556 6408 19612
rect 6344 19552 6408 19556
rect 16407 19612 16471 19616
rect 16407 19556 16411 19612
rect 16411 19556 16467 19612
rect 16467 19556 16471 19612
rect 16407 19552 16471 19556
rect 16487 19612 16551 19616
rect 16487 19556 16491 19612
rect 16491 19556 16547 19612
rect 16547 19556 16551 19612
rect 16487 19552 16551 19556
rect 16567 19612 16631 19616
rect 16567 19556 16571 19612
rect 16571 19556 16627 19612
rect 16627 19556 16631 19612
rect 16567 19552 16631 19556
rect 16647 19612 16711 19616
rect 16647 19556 16651 19612
rect 16651 19556 16707 19612
rect 16707 19556 16711 19612
rect 16647 19552 16711 19556
rect 26711 19612 26775 19616
rect 26711 19556 26715 19612
rect 26715 19556 26771 19612
rect 26771 19556 26775 19612
rect 26711 19552 26775 19556
rect 26791 19612 26855 19616
rect 26791 19556 26795 19612
rect 26795 19556 26851 19612
rect 26851 19556 26855 19612
rect 26791 19552 26855 19556
rect 26871 19612 26935 19616
rect 26871 19556 26875 19612
rect 26875 19556 26931 19612
rect 26931 19556 26935 19612
rect 26871 19552 26935 19556
rect 26951 19612 27015 19616
rect 26951 19556 26955 19612
rect 26955 19556 27011 19612
rect 27011 19556 27015 19612
rect 26951 19552 27015 19556
rect 11255 19068 11319 19072
rect 11255 19012 11259 19068
rect 11259 19012 11315 19068
rect 11315 19012 11319 19068
rect 11255 19008 11319 19012
rect 11335 19068 11399 19072
rect 11335 19012 11339 19068
rect 11339 19012 11395 19068
rect 11395 19012 11399 19068
rect 11335 19008 11399 19012
rect 11415 19068 11479 19072
rect 11415 19012 11419 19068
rect 11419 19012 11475 19068
rect 11475 19012 11479 19068
rect 11415 19008 11479 19012
rect 11495 19068 11559 19072
rect 11495 19012 11499 19068
rect 11499 19012 11555 19068
rect 11555 19012 11559 19068
rect 11495 19008 11559 19012
rect 21559 19068 21623 19072
rect 21559 19012 21563 19068
rect 21563 19012 21619 19068
rect 21619 19012 21623 19068
rect 21559 19008 21623 19012
rect 21639 19068 21703 19072
rect 21639 19012 21643 19068
rect 21643 19012 21699 19068
rect 21699 19012 21703 19068
rect 21639 19008 21703 19012
rect 21719 19068 21783 19072
rect 21719 19012 21723 19068
rect 21723 19012 21779 19068
rect 21779 19012 21783 19068
rect 21719 19008 21783 19012
rect 21799 19068 21863 19072
rect 21799 19012 21803 19068
rect 21803 19012 21859 19068
rect 21859 19012 21863 19068
rect 21799 19008 21863 19012
rect 6104 18524 6168 18528
rect 6104 18468 6108 18524
rect 6108 18468 6164 18524
rect 6164 18468 6168 18524
rect 6104 18464 6168 18468
rect 6184 18524 6248 18528
rect 6184 18468 6188 18524
rect 6188 18468 6244 18524
rect 6244 18468 6248 18524
rect 6184 18464 6248 18468
rect 6264 18524 6328 18528
rect 6264 18468 6268 18524
rect 6268 18468 6324 18524
rect 6324 18468 6328 18524
rect 6264 18464 6328 18468
rect 6344 18524 6408 18528
rect 6344 18468 6348 18524
rect 6348 18468 6404 18524
rect 6404 18468 6408 18524
rect 6344 18464 6408 18468
rect 16407 18524 16471 18528
rect 16407 18468 16411 18524
rect 16411 18468 16467 18524
rect 16467 18468 16471 18524
rect 16407 18464 16471 18468
rect 16487 18524 16551 18528
rect 16487 18468 16491 18524
rect 16491 18468 16547 18524
rect 16547 18468 16551 18524
rect 16487 18464 16551 18468
rect 16567 18524 16631 18528
rect 16567 18468 16571 18524
rect 16571 18468 16627 18524
rect 16627 18468 16631 18524
rect 16567 18464 16631 18468
rect 16647 18524 16711 18528
rect 16647 18468 16651 18524
rect 16651 18468 16707 18524
rect 16707 18468 16711 18524
rect 16647 18464 16711 18468
rect 26711 18524 26775 18528
rect 26711 18468 26715 18524
rect 26715 18468 26771 18524
rect 26771 18468 26775 18524
rect 26711 18464 26775 18468
rect 26791 18524 26855 18528
rect 26791 18468 26795 18524
rect 26795 18468 26851 18524
rect 26851 18468 26855 18524
rect 26791 18464 26855 18468
rect 26871 18524 26935 18528
rect 26871 18468 26875 18524
rect 26875 18468 26931 18524
rect 26931 18468 26935 18524
rect 26871 18464 26935 18468
rect 26951 18524 27015 18528
rect 26951 18468 26955 18524
rect 26955 18468 27011 18524
rect 27011 18468 27015 18524
rect 26951 18464 27015 18468
rect 11255 17980 11319 17984
rect 11255 17924 11259 17980
rect 11259 17924 11315 17980
rect 11315 17924 11319 17980
rect 11255 17920 11319 17924
rect 11335 17980 11399 17984
rect 11335 17924 11339 17980
rect 11339 17924 11395 17980
rect 11395 17924 11399 17980
rect 11335 17920 11399 17924
rect 11415 17980 11479 17984
rect 11415 17924 11419 17980
rect 11419 17924 11475 17980
rect 11475 17924 11479 17980
rect 11415 17920 11479 17924
rect 11495 17980 11559 17984
rect 11495 17924 11499 17980
rect 11499 17924 11555 17980
rect 11555 17924 11559 17980
rect 11495 17920 11559 17924
rect 21559 17980 21623 17984
rect 21559 17924 21563 17980
rect 21563 17924 21619 17980
rect 21619 17924 21623 17980
rect 21559 17920 21623 17924
rect 21639 17980 21703 17984
rect 21639 17924 21643 17980
rect 21643 17924 21699 17980
rect 21699 17924 21703 17980
rect 21639 17920 21703 17924
rect 21719 17980 21783 17984
rect 21719 17924 21723 17980
rect 21723 17924 21779 17980
rect 21779 17924 21783 17980
rect 21719 17920 21783 17924
rect 21799 17980 21863 17984
rect 21799 17924 21803 17980
rect 21803 17924 21859 17980
rect 21859 17924 21863 17980
rect 21799 17920 21863 17924
rect 6104 17436 6168 17440
rect 6104 17380 6108 17436
rect 6108 17380 6164 17436
rect 6164 17380 6168 17436
rect 6104 17376 6168 17380
rect 6184 17436 6248 17440
rect 6184 17380 6188 17436
rect 6188 17380 6244 17436
rect 6244 17380 6248 17436
rect 6184 17376 6248 17380
rect 6264 17436 6328 17440
rect 6264 17380 6268 17436
rect 6268 17380 6324 17436
rect 6324 17380 6328 17436
rect 6264 17376 6328 17380
rect 6344 17436 6408 17440
rect 6344 17380 6348 17436
rect 6348 17380 6404 17436
rect 6404 17380 6408 17436
rect 6344 17376 6408 17380
rect 16407 17436 16471 17440
rect 16407 17380 16411 17436
rect 16411 17380 16467 17436
rect 16467 17380 16471 17436
rect 16407 17376 16471 17380
rect 16487 17436 16551 17440
rect 16487 17380 16491 17436
rect 16491 17380 16547 17436
rect 16547 17380 16551 17436
rect 16487 17376 16551 17380
rect 16567 17436 16631 17440
rect 16567 17380 16571 17436
rect 16571 17380 16627 17436
rect 16627 17380 16631 17436
rect 16567 17376 16631 17380
rect 16647 17436 16711 17440
rect 16647 17380 16651 17436
rect 16651 17380 16707 17436
rect 16707 17380 16711 17436
rect 16647 17376 16711 17380
rect 26711 17436 26775 17440
rect 26711 17380 26715 17436
rect 26715 17380 26771 17436
rect 26771 17380 26775 17436
rect 26711 17376 26775 17380
rect 26791 17436 26855 17440
rect 26791 17380 26795 17436
rect 26795 17380 26851 17436
rect 26851 17380 26855 17436
rect 26791 17376 26855 17380
rect 26871 17436 26935 17440
rect 26871 17380 26875 17436
rect 26875 17380 26931 17436
rect 26931 17380 26935 17436
rect 26871 17376 26935 17380
rect 26951 17436 27015 17440
rect 26951 17380 26955 17436
rect 26955 17380 27011 17436
rect 27011 17380 27015 17436
rect 26951 17376 27015 17380
rect 11255 16892 11319 16896
rect 11255 16836 11259 16892
rect 11259 16836 11315 16892
rect 11315 16836 11319 16892
rect 11255 16832 11319 16836
rect 11335 16892 11399 16896
rect 11335 16836 11339 16892
rect 11339 16836 11395 16892
rect 11395 16836 11399 16892
rect 11335 16832 11399 16836
rect 11415 16892 11479 16896
rect 11415 16836 11419 16892
rect 11419 16836 11475 16892
rect 11475 16836 11479 16892
rect 11415 16832 11479 16836
rect 11495 16892 11559 16896
rect 11495 16836 11499 16892
rect 11499 16836 11555 16892
rect 11555 16836 11559 16892
rect 11495 16832 11559 16836
rect 21559 16892 21623 16896
rect 21559 16836 21563 16892
rect 21563 16836 21619 16892
rect 21619 16836 21623 16892
rect 21559 16832 21623 16836
rect 21639 16892 21703 16896
rect 21639 16836 21643 16892
rect 21643 16836 21699 16892
rect 21699 16836 21703 16892
rect 21639 16832 21703 16836
rect 21719 16892 21783 16896
rect 21719 16836 21723 16892
rect 21723 16836 21779 16892
rect 21779 16836 21783 16892
rect 21719 16832 21783 16836
rect 21799 16892 21863 16896
rect 21799 16836 21803 16892
rect 21803 16836 21859 16892
rect 21859 16836 21863 16892
rect 21799 16832 21863 16836
rect 6104 16348 6168 16352
rect 6104 16292 6108 16348
rect 6108 16292 6164 16348
rect 6164 16292 6168 16348
rect 6104 16288 6168 16292
rect 6184 16348 6248 16352
rect 6184 16292 6188 16348
rect 6188 16292 6244 16348
rect 6244 16292 6248 16348
rect 6184 16288 6248 16292
rect 6264 16348 6328 16352
rect 6264 16292 6268 16348
rect 6268 16292 6324 16348
rect 6324 16292 6328 16348
rect 6264 16288 6328 16292
rect 6344 16348 6408 16352
rect 6344 16292 6348 16348
rect 6348 16292 6404 16348
rect 6404 16292 6408 16348
rect 6344 16288 6408 16292
rect 16407 16348 16471 16352
rect 16407 16292 16411 16348
rect 16411 16292 16467 16348
rect 16467 16292 16471 16348
rect 16407 16288 16471 16292
rect 16487 16348 16551 16352
rect 16487 16292 16491 16348
rect 16491 16292 16547 16348
rect 16547 16292 16551 16348
rect 16487 16288 16551 16292
rect 16567 16348 16631 16352
rect 16567 16292 16571 16348
rect 16571 16292 16627 16348
rect 16627 16292 16631 16348
rect 16567 16288 16631 16292
rect 16647 16348 16711 16352
rect 16647 16292 16651 16348
rect 16651 16292 16707 16348
rect 16707 16292 16711 16348
rect 16647 16288 16711 16292
rect 26711 16348 26775 16352
rect 26711 16292 26715 16348
rect 26715 16292 26771 16348
rect 26771 16292 26775 16348
rect 26711 16288 26775 16292
rect 26791 16348 26855 16352
rect 26791 16292 26795 16348
rect 26795 16292 26851 16348
rect 26851 16292 26855 16348
rect 26791 16288 26855 16292
rect 26871 16348 26935 16352
rect 26871 16292 26875 16348
rect 26875 16292 26931 16348
rect 26931 16292 26935 16348
rect 26871 16288 26935 16292
rect 26951 16348 27015 16352
rect 26951 16292 26955 16348
rect 26955 16292 27011 16348
rect 27011 16292 27015 16348
rect 26951 16288 27015 16292
rect 11255 15804 11319 15808
rect 11255 15748 11259 15804
rect 11259 15748 11315 15804
rect 11315 15748 11319 15804
rect 11255 15744 11319 15748
rect 11335 15804 11399 15808
rect 11335 15748 11339 15804
rect 11339 15748 11395 15804
rect 11395 15748 11399 15804
rect 11335 15744 11399 15748
rect 11415 15804 11479 15808
rect 11415 15748 11419 15804
rect 11419 15748 11475 15804
rect 11475 15748 11479 15804
rect 11415 15744 11479 15748
rect 11495 15804 11559 15808
rect 11495 15748 11499 15804
rect 11499 15748 11555 15804
rect 11555 15748 11559 15804
rect 11495 15744 11559 15748
rect 21559 15804 21623 15808
rect 21559 15748 21563 15804
rect 21563 15748 21619 15804
rect 21619 15748 21623 15804
rect 21559 15744 21623 15748
rect 21639 15804 21703 15808
rect 21639 15748 21643 15804
rect 21643 15748 21699 15804
rect 21699 15748 21703 15804
rect 21639 15744 21703 15748
rect 21719 15804 21783 15808
rect 21719 15748 21723 15804
rect 21723 15748 21779 15804
rect 21779 15748 21783 15804
rect 21719 15744 21783 15748
rect 21799 15804 21863 15808
rect 21799 15748 21803 15804
rect 21803 15748 21859 15804
rect 21859 15748 21863 15804
rect 21799 15744 21863 15748
rect 6104 15260 6168 15264
rect 6104 15204 6108 15260
rect 6108 15204 6164 15260
rect 6164 15204 6168 15260
rect 6104 15200 6168 15204
rect 6184 15260 6248 15264
rect 6184 15204 6188 15260
rect 6188 15204 6244 15260
rect 6244 15204 6248 15260
rect 6184 15200 6248 15204
rect 6264 15260 6328 15264
rect 6264 15204 6268 15260
rect 6268 15204 6324 15260
rect 6324 15204 6328 15260
rect 6264 15200 6328 15204
rect 6344 15260 6408 15264
rect 6344 15204 6348 15260
rect 6348 15204 6404 15260
rect 6404 15204 6408 15260
rect 6344 15200 6408 15204
rect 16407 15260 16471 15264
rect 16407 15204 16411 15260
rect 16411 15204 16467 15260
rect 16467 15204 16471 15260
rect 16407 15200 16471 15204
rect 16487 15260 16551 15264
rect 16487 15204 16491 15260
rect 16491 15204 16547 15260
rect 16547 15204 16551 15260
rect 16487 15200 16551 15204
rect 16567 15260 16631 15264
rect 16567 15204 16571 15260
rect 16571 15204 16627 15260
rect 16627 15204 16631 15260
rect 16567 15200 16631 15204
rect 16647 15260 16711 15264
rect 16647 15204 16651 15260
rect 16651 15204 16707 15260
rect 16707 15204 16711 15260
rect 16647 15200 16711 15204
rect 26711 15260 26775 15264
rect 26711 15204 26715 15260
rect 26715 15204 26771 15260
rect 26771 15204 26775 15260
rect 26711 15200 26775 15204
rect 26791 15260 26855 15264
rect 26791 15204 26795 15260
rect 26795 15204 26851 15260
rect 26851 15204 26855 15260
rect 26791 15200 26855 15204
rect 26871 15260 26935 15264
rect 26871 15204 26875 15260
rect 26875 15204 26931 15260
rect 26931 15204 26935 15260
rect 26871 15200 26935 15204
rect 26951 15260 27015 15264
rect 26951 15204 26955 15260
rect 26955 15204 27011 15260
rect 27011 15204 27015 15260
rect 26951 15200 27015 15204
rect 11255 14716 11319 14720
rect 11255 14660 11259 14716
rect 11259 14660 11315 14716
rect 11315 14660 11319 14716
rect 11255 14656 11319 14660
rect 11335 14716 11399 14720
rect 11335 14660 11339 14716
rect 11339 14660 11395 14716
rect 11395 14660 11399 14716
rect 11335 14656 11399 14660
rect 11415 14716 11479 14720
rect 11415 14660 11419 14716
rect 11419 14660 11475 14716
rect 11475 14660 11479 14716
rect 11415 14656 11479 14660
rect 11495 14716 11559 14720
rect 11495 14660 11499 14716
rect 11499 14660 11555 14716
rect 11555 14660 11559 14716
rect 11495 14656 11559 14660
rect 21559 14716 21623 14720
rect 21559 14660 21563 14716
rect 21563 14660 21619 14716
rect 21619 14660 21623 14716
rect 21559 14656 21623 14660
rect 21639 14716 21703 14720
rect 21639 14660 21643 14716
rect 21643 14660 21699 14716
rect 21699 14660 21703 14716
rect 21639 14656 21703 14660
rect 21719 14716 21783 14720
rect 21719 14660 21723 14716
rect 21723 14660 21779 14716
rect 21779 14660 21783 14716
rect 21719 14656 21783 14660
rect 21799 14716 21863 14720
rect 21799 14660 21803 14716
rect 21803 14660 21859 14716
rect 21859 14660 21863 14716
rect 21799 14656 21863 14660
rect 6104 14172 6168 14176
rect 6104 14116 6108 14172
rect 6108 14116 6164 14172
rect 6164 14116 6168 14172
rect 6104 14112 6168 14116
rect 6184 14172 6248 14176
rect 6184 14116 6188 14172
rect 6188 14116 6244 14172
rect 6244 14116 6248 14172
rect 6184 14112 6248 14116
rect 6264 14172 6328 14176
rect 6264 14116 6268 14172
rect 6268 14116 6324 14172
rect 6324 14116 6328 14172
rect 6264 14112 6328 14116
rect 6344 14172 6408 14176
rect 6344 14116 6348 14172
rect 6348 14116 6404 14172
rect 6404 14116 6408 14172
rect 6344 14112 6408 14116
rect 16407 14172 16471 14176
rect 16407 14116 16411 14172
rect 16411 14116 16467 14172
rect 16467 14116 16471 14172
rect 16407 14112 16471 14116
rect 16487 14172 16551 14176
rect 16487 14116 16491 14172
rect 16491 14116 16547 14172
rect 16547 14116 16551 14172
rect 16487 14112 16551 14116
rect 16567 14172 16631 14176
rect 16567 14116 16571 14172
rect 16571 14116 16627 14172
rect 16627 14116 16631 14172
rect 16567 14112 16631 14116
rect 16647 14172 16711 14176
rect 16647 14116 16651 14172
rect 16651 14116 16707 14172
rect 16707 14116 16711 14172
rect 16647 14112 16711 14116
rect 26711 14172 26775 14176
rect 26711 14116 26715 14172
rect 26715 14116 26771 14172
rect 26771 14116 26775 14172
rect 26711 14112 26775 14116
rect 26791 14172 26855 14176
rect 26791 14116 26795 14172
rect 26795 14116 26851 14172
rect 26851 14116 26855 14172
rect 26791 14112 26855 14116
rect 26871 14172 26935 14176
rect 26871 14116 26875 14172
rect 26875 14116 26931 14172
rect 26931 14116 26935 14172
rect 26871 14112 26935 14116
rect 26951 14172 27015 14176
rect 26951 14116 26955 14172
rect 26955 14116 27011 14172
rect 27011 14116 27015 14172
rect 26951 14112 27015 14116
rect 11255 13628 11319 13632
rect 11255 13572 11259 13628
rect 11259 13572 11315 13628
rect 11315 13572 11319 13628
rect 11255 13568 11319 13572
rect 11335 13628 11399 13632
rect 11335 13572 11339 13628
rect 11339 13572 11395 13628
rect 11395 13572 11399 13628
rect 11335 13568 11399 13572
rect 11415 13628 11479 13632
rect 11415 13572 11419 13628
rect 11419 13572 11475 13628
rect 11475 13572 11479 13628
rect 11415 13568 11479 13572
rect 11495 13628 11559 13632
rect 11495 13572 11499 13628
rect 11499 13572 11555 13628
rect 11555 13572 11559 13628
rect 11495 13568 11559 13572
rect 21559 13628 21623 13632
rect 21559 13572 21563 13628
rect 21563 13572 21619 13628
rect 21619 13572 21623 13628
rect 21559 13568 21623 13572
rect 21639 13628 21703 13632
rect 21639 13572 21643 13628
rect 21643 13572 21699 13628
rect 21699 13572 21703 13628
rect 21639 13568 21703 13572
rect 21719 13628 21783 13632
rect 21719 13572 21723 13628
rect 21723 13572 21779 13628
rect 21779 13572 21783 13628
rect 21719 13568 21783 13572
rect 21799 13628 21863 13632
rect 21799 13572 21803 13628
rect 21803 13572 21859 13628
rect 21859 13572 21863 13628
rect 21799 13568 21863 13572
rect 6104 13084 6168 13088
rect 6104 13028 6108 13084
rect 6108 13028 6164 13084
rect 6164 13028 6168 13084
rect 6104 13024 6168 13028
rect 6184 13084 6248 13088
rect 6184 13028 6188 13084
rect 6188 13028 6244 13084
rect 6244 13028 6248 13084
rect 6184 13024 6248 13028
rect 6264 13084 6328 13088
rect 6264 13028 6268 13084
rect 6268 13028 6324 13084
rect 6324 13028 6328 13084
rect 6264 13024 6328 13028
rect 6344 13084 6408 13088
rect 6344 13028 6348 13084
rect 6348 13028 6404 13084
rect 6404 13028 6408 13084
rect 6344 13024 6408 13028
rect 16407 13084 16471 13088
rect 16407 13028 16411 13084
rect 16411 13028 16467 13084
rect 16467 13028 16471 13084
rect 16407 13024 16471 13028
rect 16487 13084 16551 13088
rect 16487 13028 16491 13084
rect 16491 13028 16547 13084
rect 16547 13028 16551 13084
rect 16487 13024 16551 13028
rect 16567 13084 16631 13088
rect 16567 13028 16571 13084
rect 16571 13028 16627 13084
rect 16627 13028 16631 13084
rect 16567 13024 16631 13028
rect 16647 13084 16711 13088
rect 16647 13028 16651 13084
rect 16651 13028 16707 13084
rect 16707 13028 16711 13084
rect 16647 13024 16711 13028
rect 26711 13084 26775 13088
rect 26711 13028 26715 13084
rect 26715 13028 26771 13084
rect 26771 13028 26775 13084
rect 26711 13024 26775 13028
rect 26791 13084 26855 13088
rect 26791 13028 26795 13084
rect 26795 13028 26851 13084
rect 26851 13028 26855 13084
rect 26791 13024 26855 13028
rect 26871 13084 26935 13088
rect 26871 13028 26875 13084
rect 26875 13028 26931 13084
rect 26931 13028 26935 13084
rect 26871 13024 26935 13028
rect 26951 13084 27015 13088
rect 26951 13028 26955 13084
rect 26955 13028 27011 13084
rect 27011 13028 27015 13084
rect 26951 13024 27015 13028
rect 11255 12540 11319 12544
rect 11255 12484 11259 12540
rect 11259 12484 11315 12540
rect 11315 12484 11319 12540
rect 11255 12480 11319 12484
rect 11335 12540 11399 12544
rect 11335 12484 11339 12540
rect 11339 12484 11395 12540
rect 11395 12484 11399 12540
rect 11335 12480 11399 12484
rect 11415 12540 11479 12544
rect 11415 12484 11419 12540
rect 11419 12484 11475 12540
rect 11475 12484 11479 12540
rect 11415 12480 11479 12484
rect 11495 12540 11559 12544
rect 11495 12484 11499 12540
rect 11499 12484 11555 12540
rect 11555 12484 11559 12540
rect 11495 12480 11559 12484
rect 21559 12540 21623 12544
rect 21559 12484 21563 12540
rect 21563 12484 21619 12540
rect 21619 12484 21623 12540
rect 21559 12480 21623 12484
rect 21639 12540 21703 12544
rect 21639 12484 21643 12540
rect 21643 12484 21699 12540
rect 21699 12484 21703 12540
rect 21639 12480 21703 12484
rect 21719 12540 21783 12544
rect 21719 12484 21723 12540
rect 21723 12484 21779 12540
rect 21779 12484 21783 12540
rect 21719 12480 21783 12484
rect 21799 12540 21863 12544
rect 21799 12484 21803 12540
rect 21803 12484 21859 12540
rect 21859 12484 21863 12540
rect 21799 12480 21863 12484
rect 6104 11996 6168 12000
rect 6104 11940 6108 11996
rect 6108 11940 6164 11996
rect 6164 11940 6168 11996
rect 6104 11936 6168 11940
rect 6184 11996 6248 12000
rect 6184 11940 6188 11996
rect 6188 11940 6244 11996
rect 6244 11940 6248 11996
rect 6184 11936 6248 11940
rect 6264 11996 6328 12000
rect 6264 11940 6268 11996
rect 6268 11940 6324 11996
rect 6324 11940 6328 11996
rect 6264 11936 6328 11940
rect 6344 11996 6408 12000
rect 6344 11940 6348 11996
rect 6348 11940 6404 11996
rect 6404 11940 6408 11996
rect 6344 11936 6408 11940
rect 16407 11996 16471 12000
rect 16407 11940 16411 11996
rect 16411 11940 16467 11996
rect 16467 11940 16471 11996
rect 16407 11936 16471 11940
rect 16487 11996 16551 12000
rect 16487 11940 16491 11996
rect 16491 11940 16547 11996
rect 16547 11940 16551 11996
rect 16487 11936 16551 11940
rect 16567 11996 16631 12000
rect 16567 11940 16571 11996
rect 16571 11940 16627 11996
rect 16627 11940 16631 11996
rect 16567 11936 16631 11940
rect 16647 11996 16711 12000
rect 16647 11940 16651 11996
rect 16651 11940 16707 11996
rect 16707 11940 16711 11996
rect 16647 11936 16711 11940
rect 26711 11996 26775 12000
rect 26711 11940 26715 11996
rect 26715 11940 26771 11996
rect 26771 11940 26775 11996
rect 26711 11936 26775 11940
rect 26791 11996 26855 12000
rect 26791 11940 26795 11996
rect 26795 11940 26851 11996
rect 26851 11940 26855 11996
rect 26791 11936 26855 11940
rect 26871 11996 26935 12000
rect 26871 11940 26875 11996
rect 26875 11940 26931 11996
rect 26931 11940 26935 11996
rect 26871 11936 26935 11940
rect 26951 11996 27015 12000
rect 26951 11940 26955 11996
rect 26955 11940 27011 11996
rect 27011 11940 27015 11996
rect 26951 11936 27015 11940
rect 11255 11452 11319 11456
rect 11255 11396 11259 11452
rect 11259 11396 11315 11452
rect 11315 11396 11319 11452
rect 11255 11392 11319 11396
rect 11335 11452 11399 11456
rect 11335 11396 11339 11452
rect 11339 11396 11395 11452
rect 11395 11396 11399 11452
rect 11335 11392 11399 11396
rect 11415 11452 11479 11456
rect 11415 11396 11419 11452
rect 11419 11396 11475 11452
rect 11475 11396 11479 11452
rect 11415 11392 11479 11396
rect 11495 11452 11559 11456
rect 11495 11396 11499 11452
rect 11499 11396 11555 11452
rect 11555 11396 11559 11452
rect 11495 11392 11559 11396
rect 21559 11452 21623 11456
rect 21559 11396 21563 11452
rect 21563 11396 21619 11452
rect 21619 11396 21623 11452
rect 21559 11392 21623 11396
rect 21639 11452 21703 11456
rect 21639 11396 21643 11452
rect 21643 11396 21699 11452
rect 21699 11396 21703 11452
rect 21639 11392 21703 11396
rect 21719 11452 21783 11456
rect 21719 11396 21723 11452
rect 21723 11396 21779 11452
rect 21779 11396 21783 11452
rect 21719 11392 21783 11396
rect 21799 11452 21863 11456
rect 21799 11396 21803 11452
rect 21803 11396 21859 11452
rect 21859 11396 21863 11452
rect 21799 11392 21863 11396
rect 6104 10908 6168 10912
rect 6104 10852 6108 10908
rect 6108 10852 6164 10908
rect 6164 10852 6168 10908
rect 6104 10848 6168 10852
rect 6184 10908 6248 10912
rect 6184 10852 6188 10908
rect 6188 10852 6244 10908
rect 6244 10852 6248 10908
rect 6184 10848 6248 10852
rect 6264 10908 6328 10912
rect 6264 10852 6268 10908
rect 6268 10852 6324 10908
rect 6324 10852 6328 10908
rect 6264 10848 6328 10852
rect 6344 10908 6408 10912
rect 6344 10852 6348 10908
rect 6348 10852 6404 10908
rect 6404 10852 6408 10908
rect 6344 10848 6408 10852
rect 16407 10908 16471 10912
rect 16407 10852 16411 10908
rect 16411 10852 16467 10908
rect 16467 10852 16471 10908
rect 16407 10848 16471 10852
rect 16487 10908 16551 10912
rect 16487 10852 16491 10908
rect 16491 10852 16547 10908
rect 16547 10852 16551 10908
rect 16487 10848 16551 10852
rect 16567 10908 16631 10912
rect 16567 10852 16571 10908
rect 16571 10852 16627 10908
rect 16627 10852 16631 10908
rect 16567 10848 16631 10852
rect 16647 10908 16711 10912
rect 16647 10852 16651 10908
rect 16651 10852 16707 10908
rect 16707 10852 16711 10908
rect 16647 10848 16711 10852
rect 26711 10908 26775 10912
rect 26711 10852 26715 10908
rect 26715 10852 26771 10908
rect 26771 10852 26775 10908
rect 26711 10848 26775 10852
rect 26791 10908 26855 10912
rect 26791 10852 26795 10908
rect 26795 10852 26851 10908
rect 26851 10852 26855 10908
rect 26791 10848 26855 10852
rect 26871 10908 26935 10912
rect 26871 10852 26875 10908
rect 26875 10852 26931 10908
rect 26931 10852 26935 10908
rect 26871 10848 26935 10852
rect 26951 10908 27015 10912
rect 26951 10852 26955 10908
rect 26955 10852 27011 10908
rect 27011 10852 27015 10908
rect 26951 10848 27015 10852
rect 11255 10364 11319 10368
rect 11255 10308 11259 10364
rect 11259 10308 11315 10364
rect 11315 10308 11319 10364
rect 11255 10304 11319 10308
rect 11335 10364 11399 10368
rect 11335 10308 11339 10364
rect 11339 10308 11395 10364
rect 11395 10308 11399 10364
rect 11335 10304 11399 10308
rect 11415 10364 11479 10368
rect 11415 10308 11419 10364
rect 11419 10308 11475 10364
rect 11475 10308 11479 10364
rect 11415 10304 11479 10308
rect 11495 10364 11559 10368
rect 11495 10308 11499 10364
rect 11499 10308 11555 10364
rect 11555 10308 11559 10364
rect 11495 10304 11559 10308
rect 21559 10364 21623 10368
rect 21559 10308 21563 10364
rect 21563 10308 21619 10364
rect 21619 10308 21623 10364
rect 21559 10304 21623 10308
rect 21639 10364 21703 10368
rect 21639 10308 21643 10364
rect 21643 10308 21699 10364
rect 21699 10308 21703 10364
rect 21639 10304 21703 10308
rect 21719 10364 21783 10368
rect 21719 10308 21723 10364
rect 21723 10308 21779 10364
rect 21779 10308 21783 10364
rect 21719 10304 21783 10308
rect 21799 10364 21863 10368
rect 21799 10308 21803 10364
rect 21803 10308 21859 10364
rect 21859 10308 21863 10364
rect 21799 10304 21863 10308
rect 6104 9820 6168 9824
rect 6104 9764 6108 9820
rect 6108 9764 6164 9820
rect 6164 9764 6168 9820
rect 6104 9760 6168 9764
rect 6184 9820 6248 9824
rect 6184 9764 6188 9820
rect 6188 9764 6244 9820
rect 6244 9764 6248 9820
rect 6184 9760 6248 9764
rect 6264 9820 6328 9824
rect 6264 9764 6268 9820
rect 6268 9764 6324 9820
rect 6324 9764 6328 9820
rect 6264 9760 6328 9764
rect 6344 9820 6408 9824
rect 6344 9764 6348 9820
rect 6348 9764 6404 9820
rect 6404 9764 6408 9820
rect 6344 9760 6408 9764
rect 16407 9820 16471 9824
rect 16407 9764 16411 9820
rect 16411 9764 16467 9820
rect 16467 9764 16471 9820
rect 16407 9760 16471 9764
rect 16487 9820 16551 9824
rect 16487 9764 16491 9820
rect 16491 9764 16547 9820
rect 16547 9764 16551 9820
rect 16487 9760 16551 9764
rect 16567 9820 16631 9824
rect 16567 9764 16571 9820
rect 16571 9764 16627 9820
rect 16627 9764 16631 9820
rect 16567 9760 16631 9764
rect 16647 9820 16711 9824
rect 16647 9764 16651 9820
rect 16651 9764 16707 9820
rect 16707 9764 16711 9820
rect 16647 9760 16711 9764
rect 26711 9820 26775 9824
rect 26711 9764 26715 9820
rect 26715 9764 26771 9820
rect 26771 9764 26775 9820
rect 26711 9760 26775 9764
rect 26791 9820 26855 9824
rect 26791 9764 26795 9820
rect 26795 9764 26851 9820
rect 26851 9764 26855 9820
rect 26791 9760 26855 9764
rect 26871 9820 26935 9824
rect 26871 9764 26875 9820
rect 26875 9764 26931 9820
rect 26931 9764 26935 9820
rect 26871 9760 26935 9764
rect 26951 9820 27015 9824
rect 26951 9764 26955 9820
rect 26955 9764 27011 9820
rect 27011 9764 27015 9820
rect 26951 9760 27015 9764
rect 11255 9276 11319 9280
rect 11255 9220 11259 9276
rect 11259 9220 11315 9276
rect 11315 9220 11319 9276
rect 11255 9216 11319 9220
rect 11335 9276 11399 9280
rect 11335 9220 11339 9276
rect 11339 9220 11395 9276
rect 11395 9220 11399 9276
rect 11335 9216 11399 9220
rect 11415 9276 11479 9280
rect 11415 9220 11419 9276
rect 11419 9220 11475 9276
rect 11475 9220 11479 9276
rect 11415 9216 11479 9220
rect 11495 9276 11559 9280
rect 11495 9220 11499 9276
rect 11499 9220 11555 9276
rect 11555 9220 11559 9276
rect 11495 9216 11559 9220
rect 21559 9276 21623 9280
rect 21559 9220 21563 9276
rect 21563 9220 21619 9276
rect 21619 9220 21623 9276
rect 21559 9216 21623 9220
rect 21639 9276 21703 9280
rect 21639 9220 21643 9276
rect 21643 9220 21699 9276
rect 21699 9220 21703 9276
rect 21639 9216 21703 9220
rect 21719 9276 21783 9280
rect 21719 9220 21723 9276
rect 21723 9220 21779 9276
rect 21779 9220 21783 9276
rect 21719 9216 21783 9220
rect 21799 9276 21863 9280
rect 21799 9220 21803 9276
rect 21803 9220 21859 9276
rect 21859 9220 21863 9276
rect 21799 9216 21863 9220
rect 6104 8732 6168 8736
rect 6104 8676 6108 8732
rect 6108 8676 6164 8732
rect 6164 8676 6168 8732
rect 6104 8672 6168 8676
rect 6184 8732 6248 8736
rect 6184 8676 6188 8732
rect 6188 8676 6244 8732
rect 6244 8676 6248 8732
rect 6184 8672 6248 8676
rect 6264 8732 6328 8736
rect 6264 8676 6268 8732
rect 6268 8676 6324 8732
rect 6324 8676 6328 8732
rect 6264 8672 6328 8676
rect 6344 8732 6408 8736
rect 6344 8676 6348 8732
rect 6348 8676 6404 8732
rect 6404 8676 6408 8732
rect 6344 8672 6408 8676
rect 16407 8732 16471 8736
rect 16407 8676 16411 8732
rect 16411 8676 16467 8732
rect 16467 8676 16471 8732
rect 16407 8672 16471 8676
rect 16487 8732 16551 8736
rect 16487 8676 16491 8732
rect 16491 8676 16547 8732
rect 16547 8676 16551 8732
rect 16487 8672 16551 8676
rect 16567 8732 16631 8736
rect 16567 8676 16571 8732
rect 16571 8676 16627 8732
rect 16627 8676 16631 8732
rect 16567 8672 16631 8676
rect 16647 8732 16711 8736
rect 16647 8676 16651 8732
rect 16651 8676 16707 8732
rect 16707 8676 16711 8732
rect 16647 8672 16711 8676
rect 26711 8732 26775 8736
rect 26711 8676 26715 8732
rect 26715 8676 26771 8732
rect 26771 8676 26775 8732
rect 26711 8672 26775 8676
rect 26791 8732 26855 8736
rect 26791 8676 26795 8732
rect 26795 8676 26851 8732
rect 26851 8676 26855 8732
rect 26791 8672 26855 8676
rect 26871 8732 26935 8736
rect 26871 8676 26875 8732
rect 26875 8676 26931 8732
rect 26931 8676 26935 8732
rect 26871 8672 26935 8676
rect 26951 8732 27015 8736
rect 26951 8676 26955 8732
rect 26955 8676 27011 8732
rect 27011 8676 27015 8732
rect 26951 8672 27015 8676
rect 11255 8188 11319 8192
rect 11255 8132 11259 8188
rect 11259 8132 11315 8188
rect 11315 8132 11319 8188
rect 11255 8128 11319 8132
rect 11335 8188 11399 8192
rect 11335 8132 11339 8188
rect 11339 8132 11395 8188
rect 11395 8132 11399 8188
rect 11335 8128 11399 8132
rect 11415 8188 11479 8192
rect 11415 8132 11419 8188
rect 11419 8132 11475 8188
rect 11475 8132 11479 8188
rect 11415 8128 11479 8132
rect 11495 8188 11559 8192
rect 11495 8132 11499 8188
rect 11499 8132 11555 8188
rect 11555 8132 11559 8188
rect 11495 8128 11559 8132
rect 21559 8188 21623 8192
rect 21559 8132 21563 8188
rect 21563 8132 21619 8188
rect 21619 8132 21623 8188
rect 21559 8128 21623 8132
rect 21639 8188 21703 8192
rect 21639 8132 21643 8188
rect 21643 8132 21699 8188
rect 21699 8132 21703 8188
rect 21639 8128 21703 8132
rect 21719 8188 21783 8192
rect 21719 8132 21723 8188
rect 21723 8132 21779 8188
rect 21779 8132 21783 8188
rect 21719 8128 21783 8132
rect 21799 8188 21863 8192
rect 21799 8132 21803 8188
rect 21803 8132 21859 8188
rect 21859 8132 21863 8188
rect 21799 8128 21863 8132
rect 6104 7644 6168 7648
rect 6104 7588 6108 7644
rect 6108 7588 6164 7644
rect 6164 7588 6168 7644
rect 6104 7584 6168 7588
rect 6184 7644 6248 7648
rect 6184 7588 6188 7644
rect 6188 7588 6244 7644
rect 6244 7588 6248 7644
rect 6184 7584 6248 7588
rect 6264 7644 6328 7648
rect 6264 7588 6268 7644
rect 6268 7588 6324 7644
rect 6324 7588 6328 7644
rect 6264 7584 6328 7588
rect 6344 7644 6408 7648
rect 6344 7588 6348 7644
rect 6348 7588 6404 7644
rect 6404 7588 6408 7644
rect 6344 7584 6408 7588
rect 16407 7644 16471 7648
rect 16407 7588 16411 7644
rect 16411 7588 16467 7644
rect 16467 7588 16471 7644
rect 16407 7584 16471 7588
rect 16487 7644 16551 7648
rect 16487 7588 16491 7644
rect 16491 7588 16547 7644
rect 16547 7588 16551 7644
rect 16487 7584 16551 7588
rect 16567 7644 16631 7648
rect 16567 7588 16571 7644
rect 16571 7588 16627 7644
rect 16627 7588 16631 7644
rect 16567 7584 16631 7588
rect 16647 7644 16711 7648
rect 16647 7588 16651 7644
rect 16651 7588 16707 7644
rect 16707 7588 16711 7644
rect 16647 7584 16711 7588
rect 26711 7644 26775 7648
rect 26711 7588 26715 7644
rect 26715 7588 26771 7644
rect 26771 7588 26775 7644
rect 26711 7584 26775 7588
rect 26791 7644 26855 7648
rect 26791 7588 26795 7644
rect 26795 7588 26851 7644
rect 26851 7588 26855 7644
rect 26791 7584 26855 7588
rect 26871 7644 26935 7648
rect 26871 7588 26875 7644
rect 26875 7588 26931 7644
rect 26931 7588 26935 7644
rect 26871 7584 26935 7588
rect 26951 7644 27015 7648
rect 26951 7588 26955 7644
rect 26955 7588 27011 7644
rect 27011 7588 27015 7644
rect 26951 7584 27015 7588
rect 11255 7100 11319 7104
rect 11255 7044 11259 7100
rect 11259 7044 11315 7100
rect 11315 7044 11319 7100
rect 11255 7040 11319 7044
rect 11335 7100 11399 7104
rect 11335 7044 11339 7100
rect 11339 7044 11395 7100
rect 11395 7044 11399 7100
rect 11335 7040 11399 7044
rect 11415 7100 11479 7104
rect 11415 7044 11419 7100
rect 11419 7044 11475 7100
rect 11475 7044 11479 7100
rect 11415 7040 11479 7044
rect 11495 7100 11559 7104
rect 11495 7044 11499 7100
rect 11499 7044 11555 7100
rect 11555 7044 11559 7100
rect 11495 7040 11559 7044
rect 21559 7100 21623 7104
rect 21559 7044 21563 7100
rect 21563 7044 21619 7100
rect 21619 7044 21623 7100
rect 21559 7040 21623 7044
rect 21639 7100 21703 7104
rect 21639 7044 21643 7100
rect 21643 7044 21699 7100
rect 21699 7044 21703 7100
rect 21639 7040 21703 7044
rect 21719 7100 21783 7104
rect 21719 7044 21723 7100
rect 21723 7044 21779 7100
rect 21779 7044 21783 7100
rect 21719 7040 21783 7044
rect 21799 7100 21863 7104
rect 21799 7044 21803 7100
rect 21803 7044 21859 7100
rect 21859 7044 21863 7100
rect 21799 7040 21863 7044
rect 6104 6556 6168 6560
rect 6104 6500 6108 6556
rect 6108 6500 6164 6556
rect 6164 6500 6168 6556
rect 6104 6496 6168 6500
rect 6184 6556 6248 6560
rect 6184 6500 6188 6556
rect 6188 6500 6244 6556
rect 6244 6500 6248 6556
rect 6184 6496 6248 6500
rect 6264 6556 6328 6560
rect 6264 6500 6268 6556
rect 6268 6500 6324 6556
rect 6324 6500 6328 6556
rect 6264 6496 6328 6500
rect 6344 6556 6408 6560
rect 6344 6500 6348 6556
rect 6348 6500 6404 6556
rect 6404 6500 6408 6556
rect 6344 6496 6408 6500
rect 16407 6556 16471 6560
rect 16407 6500 16411 6556
rect 16411 6500 16467 6556
rect 16467 6500 16471 6556
rect 16407 6496 16471 6500
rect 16487 6556 16551 6560
rect 16487 6500 16491 6556
rect 16491 6500 16547 6556
rect 16547 6500 16551 6556
rect 16487 6496 16551 6500
rect 16567 6556 16631 6560
rect 16567 6500 16571 6556
rect 16571 6500 16627 6556
rect 16627 6500 16631 6556
rect 16567 6496 16631 6500
rect 16647 6556 16711 6560
rect 16647 6500 16651 6556
rect 16651 6500 16707 6556
rect 16707 6500 16711 6556
rect 16647 6496 16711 6500
rect 26711 6556 26775 6560
rect 26711 6500 26715 6556
rect 26715 6500 26771 6556
rect 26771 6500 26775 6556
rect 26711 6496 26775 6500
rect 26791 6556 26855 6560
rect 26791 6500 26795 6556
rect 26795 6500 26851 6556
rect 26851 6500 26855 6556
rect 26791 6496 26855 6500
rect 26871 6556 26935 6560
rect 26871 6500 26875 6556
rect 26875 6500 26931 6556
rect 26931 6500 26935 6556
rect 26871 6496 26935 6500
rect 26951 6556 27015 6560
rect 26951 6500 26955 6556
rect 26955 6500 27011 6556
rect 27011 6500 27015 6556
rect 26951 6496 27015 6500
rect 11255 6012 11319 6016
rect 11255 5956 11259 6012
rect 11259 5956 11315 6012
rect 11315 5956 11319 6012
rect 11255 5952 11319 5956
rect 11335 6012 11399 6016
rect 11335 5956 11339 6012
rect 11339 5956 11395 6012
rect 11395 5956 11399 6012
rect 11335 5952 11399 5956
rect 11415 6012 11479 6016
rect 11415 5956 11419 6012
rect 11419 5956 11475 6012
rect 11475 5956 11479 6012
rect 11415 5952 11479 5956
rect 11495 6012 11559 6016
rect 11495 5956 11499 6012
rect 11499 5956 11555 6012
rect 11555 5956 11559 6012
rect 11495 5952 11559 5956
rect 21559 6012 21623 6016
rect 21559 5956 21563 6012
rect 21563 5956 21619 6012
rect 21619 5956 21623 6012
rect 21559 5952 21623 5956
rect 21639 6012 21703 6016
rect 21639 5956 21643 6012
rect 21643 5956 21699 6012
rect 21699 5956 21703 6012
rect 21639 5952 21703 5956
rect 21719 6012 21783 6016
rect 21719 5956 21723 6012
rect 21723 5956 21779 6012
rect 21779 5956 21783 6012
rect 21719 5952 21783 5956
rect 21799 6012 21863 6016
rect 21799 5956 21803 6012
rect 21803 5956 21859 6012
rect 21859 5956 21863 6012
rect 21799 5952 21863 5956
rect 6104 5468 6168 5472
rect 6104 5412 6108 5468
rect 6108 5412 6164 5468
rect 6164 5412 6168 5468
rect 6104 5408 6168 5412
rect 6184 5468 6248 5472
rect 6184 5412 6188 5468
rect 6188 5412 6244 5468
rect 6244 5412 6248 5468
rect 6184 5408 6248 5412
rect 6264 5468 6328 5472
rect 6264 5412 6268 5468
rect 6268 5412 6324 5468
rect 6324 5412 6328 5468
rect 6264 5408 6328 5412
rect 6344 5468 6408 5472
rect 6344 5412 6348 5468
rect 6348 5412 6404 5468
rect 6404 5412 6408 5468
rect 6344 5408 6408 5412
rect 16407 5468 16471 5472
rect 16407 5412 16411 5468
rect 16411 5412 16467 5468
rect 16467 5412 16471 5468
rect 16407 5408 16471 5412
rect 16487 5468 16551 5472
rect 16487 5412 16491 5468
rect 16491 5412 16547 5468
rect 16547 5412 16551 5468
rect 16487 5408 16551 5412
rect 16567 5468 16631 5472
rect 16567 5412 16571 5468
rect 16571 5412 16627 5468
rect 16627 5412 16631 5468
rect 16567 5408 16631 5412
rect 16647 5468 16711 5472
rect 16647 5412 16651 5468
rect 16651 5412 16707 5468
rect 16707 5412 16711 5468
rect 16647 5408 16711 5412
rect 26711 5468 26775 5472
rect 26711 5412 26715 5468
rect 26715 5412 26771 5468
rect 26771 5412 26775 5468
rect 26711 5408 26775 5412
rect 26791 5468 26855 5472
rect 26791 5412 26795 5468
rect 26795 5412 26851 5468
rect 26851 5412 26855 5468
rect 26791 5408 26855 5412
rect 26871 5468 26935 5472
rect 26871 5412 26875 5468
rect 26875 5412 26931 5468
rect 26931 5412 26935 5468
rect 26871 5408 26935 5412
rect 26951 5468 27015 5472
rect 26951 5412 26955 5468
rect 26955 5412 27011 5468
rect 27011 5412 27015 5468
rect 26951 5408 27015 5412
rect 11255 4924 11319 4928
rect 11255 4868 11259 4924
rect 11259 4868 11315 4924
rect 11315 4868 11319 4924
rect 11255 4864 11319 4868
rect 11335 4924 11399 4928
rect 11335 4868 11339 4924
rect 11339 4868 11395 4924
rect 11395 4868 11399 4924
rect 11335 4864 11399 4868
rect 11415 4924 11479 4928
rect 11415 4868 11419 4924
rect 11419 4868 11475 4924
rect 11475 4868 11479 4924
rect 11415 4864 11479 4868
rect 11495 4924 11559 4928
rect 11495 4868 11499 4924
rect 11499 4868 11555 4924
rect 11555 4868 11559 4924
rect 11495 4864 11559 4868
rect 21559 4924 21623 4928
rect 21559 4868 21563 4924
rect 21563 4868 21619 4924
rect 21619 4868 21623 4924
rect 21559 4864 21623 4868
rect 21639 4924 21703 4928
rect 21639 4868 21643 4924
rect 21643 4868 21699 4924
rect 21699 4868 21703 4924
rect 21639 4864 21703 4868
rect 21719 4924 21783 4928
rect 21719 4868 21723 4924
rect 21723 4868 21779 4924
rect 21779 4868 21783 4924
rect 21719 4864 21783 4868
rect 21799 4924 21863 4928
rect 21799 4868 21803 4924
rect 21803 4868 21859 4924
rect 21859 4868 21863 4924
rect 21799 4864 21863 4868
rect 6104 4380 6168 4384
rect 6104 4324 6108 4380
rect 6108 4324 6164 4380
rect 6164 4324 6168 4380
rect 6104 4320 6168 4324
rect 6184 4380 6248 4384
rect 6184 4324 6188 4380
rect 6188 4324 6244 4380
rect 6244 4324 6248 4380
rect 6184 4320 6248 4324
rect 6264 4380 6328 4384
rect 6264 4324 6268 4380
rect 6268 4324 6324 4380
rect 6324 4324 6328 4380
rect 6264 4320 6328 4324
rect 6344 4380 6408 4384
rect 6344 4324 6348 4380
rect 6348 4324 6404 4380
rect 6404 4324 6408 4380
rect 6344 4320 6408 4324
rect 16407 4380 16471 4384
rect 16407 4324 16411 4380
rect 16411 4324 16467 4380
rect 16467 4324 16471 4380
rect 16407 4320 16471 4324
rect 16487 4380 16551 4384
rect 16487 4324 16491 4380
rect 16491 4324 16547 4380
rect 16547 4324 16551 4380
rect 16487 4320 16551 4324
rect 16567 4380 16631 4384
rect 16567 4324 16571 4380
rect 16571 4324 16627 4380
rect 16627 4324 16631 4380
rect 16567 4320 16631 4324
rect 16647 4380 16711 4384
rect 16647 4324 16651 4380
rect 16651 4324 16707 4380
rect 16707 4324 16711 4380
rect 16647 4320 16711 4324
rect 26711 4380 26775 4384
rect 26711 4324 26715 4380
rect 26715 4324 26771 4380
rect 26771 4324 26775 4380
rect 26711 4320 26775 4324
rect 26791 4380 26855 4384
rect 26791 4324 26795 4380
rect 26795 4324 26851 4380
rect 26851 4324 26855 4380
rect 26791 4320 26855 4324
rect 26871 4380 26935 4384
rect 26871 4324 26875 4380
rect 26875 4324 26931 4380
rect 26931 4324 26935 4380
rect 26871 4320 26935 4324
rect 26951 4380 27015 4384
rect 26951 4324 26955 4380
rect 26955 4324 27011 4380
rect 27011 4324 27015 4380
rect 26951 4320 27015 4324
rect 11255 3836 11319 3840
rect 11255 3780 11259 3836
rect 11259 3780 11315 3836
rect 11315 3780 11319 3836
rect 11255 3776 11319 3780
rect 11335 3836 11399 3840
rect 11335 3780 11339 3836
rect 11339 3780 11395 3836
rect 11395 3780 11399 3836
rect 11335 3776 11399 3780
rect 11415 3836 11479 3840
rect 11415 3780 11419 3836
rect 11419 3780 11475 3836
rect 11475 3780 11479 3836
rect 11415 3776 11479 3780
rect 11495 3836 11559 3840
rect 11495 3780 11499 3836
rect 11499 3780 11555 3836
rect 11555 3780 11559 3836
rect 11495 3776 11559 3780
rect 21559 3836 21623 3840
rect 21559 3780 21563 3836
rect 21563 3780 21619 3836
rect 21619 3780 21623 3836
rect 21559 3776 21623 3780
rect 21639 3836 21703 3840
rect 21639 3780 21643 3836
rect 21643 3780 21699 3836
rect 21699 3780 21703 3836
rect 21639 3776 21703 3780
rect 21719 3836 21783 3840
rect 21719 3780 21723 3836
rect 21723 3780 21779 3836
rect 21779 3780 21783 3836
rect 21719 3776 21783 3780
rect 21799 3836 21863 3840
rect 21799 3780 21803 3836
rect 21803 3780 21859 3836
rect 21859 3780 21863 3836
rect 21799 3776 21863 3780
rect 6104 3292 6168 3296
rect 6104 3236 6108 3292
rect 6108 3236 6164 3292
rect 6164 3236 6168 3292
rect 6104 3232 6168 3236
rect 6184 3292 6248 3296
rect 6184 3236 6188 3292
rect 6188 3236 6244 3292
rect 6244 3236 6248 3292
rect 6184 3232 6248 3236
rect 6264 3292 6328 3296
rect 6264 3236 6268 3292
rect 6268 3236 6324 3292
rect 6324 3236 6328 3292
rect 6264 3232 6328 3236
rect 6344 3292 6408 3296
rect 6344 3236 6348 3292
rect 6348 3236 6404 3292
rect 6404 3236 6408 3292
rect 6344 3232 6408 3236
rect 16407 3292 16471 3296
rect 16407 3236 16411 3292
rect 16411 3236 16467 3292
rect 16467 3236 16471 3292
rect 16407 3232 16471 3236
rect 16487 3292 16551 3296
rect 16487 3236 16491 3292
rect 16491 3236 16547 3292
rect 16547 3236 16551 3292
rect 16487 3232 16551 3236
rect 16567 3292 16631 3296
rect 16567 3236 16571 3292
rect 16571 3236 16627 3292
rect 16627 3236 16631 3292
rect 16567 3232 16631 3236
rect 16647 3292 16711 3296
rect 16647 3236 16651 3292
rect 16651 3236 16707 3292
rect 16707 3236 16711 3292
rect 16647 3232 16711 3236
rect 26711 3292 26775 3296
rect 26711 3236 26715 3292
rect 26715 3236 26771 3292
rect 26771 3236 26775 3292
rect 26711 3232 26775 3236
rect 26791 3292 26855 3296
rect 26791 3236 26795 3292
rect 26795 3236 26851 3292
rect 26851 3236 26855 3292
rect 26791 3232 26855 3236
rect 26871 3292 26935 3296
rect 26871 3236 26875 3292
rect 26875 3236 26931 3292
rect 26931 3236 26935 3292
rect 26871 3232 26935 3236
rect 26951 3292 27015 3296
rect 26951 3236 26955 3292
rect 26955 3236 27011 3292
rect 27011 3236 27015 3292
rect 26951 3232 27015 3236
rect 11255 2748 11319 2752
rect 11255 2692 11259 2748
rect 11259 2692 11315 2748
rect 11315 2692 11319 2748
rect 11255 2688 11319 2692
rect 11335 2748 11399 2752
rect 11335 2692 11339 2748
rect 11339 2692 11395 2748
rect 11395 2692 11399 2748
rect 11335 2688 11399 2692
rect 11415 2748 11479 2752
rect 11415 2692 11419 2748
rect 11419 2692 11475 2748
rect 11475 2692 11479 2748
rect 11415 2688 11479 2692
rect 11495 2748 11559 2752
rect 11495 2692 11499 2748
rect 11499 2692 11555 2748
rect 11555 2692 11559 2748
rect 11495 2688 11559 2692
rect 21559 2748 21623 2752
rect 21559 2692 21563 2748
rect 21563 2692 21619 2748
rect 21619 2692 21623 2748
rect 21559 2688 21623 2692
rect 21639 2748 21703 2752
rect 21639 2692 21643 2748
rect 21643 2692 21699 2748
rect 21699 2692 21703 2748
rect 21639 2688 21703 2692
rect 21719 2748 21783 2752
rect 21719 2692 21723 2748
rect 21723 2692 21779 2748
rect 21779 2692 21783 2748
rect 21719 2688 21783 2692
rect 21799 2748 21863 2752
rect 21799 2692 21803 2748
rect 21803 2692 21859 2748
rect 21859 2692 21863 2748
rect 21799 2688 21863 2692
rect 6104 2204 6168 2208
rect 6104 2148 6108 2204
rect 6108 2148 6164 2204
rect 6164 2148 6168 2204
rect 6104 2144 6168 2148
rect 6184 2204 6248 2208
rect 6184 2148 6188 2204
rect 6188 2148 6244 2204
rect 6244 2148 6248 2204
rect 6184 2144 6248 2148
rect 6264 2204 6328 2208
rect 6264 2148 6268 2204
rect 6268 2148 6324 2204
rect 6324 2148 6328 2204
rect 6264 2144 6328 2148
rect 6344 2204 6408 2208
rect 6344 2148 6348 2204
rect 6348 2148 6404 2204
rect 6404 2148 6408 2204
rect 6344 2144 6408 2148
rect 16407 2204 16471 2208
rect 16407 2148 16411 2204
rect 16411 2148 16467 2204
rect 16467 2148 16471 2204
rect 16407 2144 16471 2148
rect 16487 2204 16551 2208
rect 16487 2148 16491 2204
rect 16491 2148 16547 2204
rect 16547 2148 16551 2204
rect 16487 2144 16551 2148
rect 16567 2204 16631 2208
rect 16567 2148 16571 2204
rect 16571 2148 16627 2204
rect 16627 2148 16631 2204
rect 16567 2144 16631 2148
rect 16647 2204 16711 2208
rect 16647 2148 16651 2204
rect 16651 2148 16707 2204
rect 16707 2148 16711 2204
rect 16647 2144 16711 2148
rect 26711 2204 26775 2208
rect 26711 2148 26715 2204
rect 26715 2148 26771 2204
rect 26771 2148 26775 2204
rect 26711 2144 26775 2148
rect 26791 2204 26855 2208
rect 26791 2148 26795 2204
rect 26795 2148 26851 2204
rect 26851 2148 26855 2204
rect 26791 2144 26855 2148
rect 26871 2204 26935 2208
rect 26871 2148 26875 2204
rect 26875 2148 26931 2204
rect 26931 2148 26935 2204
rect 26871 2144 26935 2148
rect 26951 2204 27015 2208
rect 26951 2148 26955 2204
rect 26955 2148 27011 2204
rect 27011 2148 27015 2204
rect 26951 2144 27015 2148
rect 11255 1660 11319 1664
rect 11255 1604 11259 1660
rect 11259 1604 11315 1660
rect 11315 1604 11319 1660
rect 11255 1600 11319 1604
rect 11335 1660 11399 1664
rect 11335 1604 11339 1660
rect 11339 1604 11395 1660
rect 11395 1604 11399 1660
rect 11335 1600 11399 1604
rect 11415 1660 11479 1664
rect 11415 1604 11419 1660
rect 11419 1604 11475 1660
rect 11475 1604 11479 1660
rect 11415 1600 11479 1604
rect 11495 1660 11559 1664
rect 11495 1604 11499 1660
rect 11499 1604 11555 1660
rect 11555 1604 11559 1660
rect 11495 1600 11559 1604
rect 21559 1660 21623 1664
rect 21559 1604 21563 1660
rect 21563 1604 21619 1660
rect 21619 1604 21623 1660
rect 21559 1600 21623 1604
rect 21639 1660 21703 1664
rect 21639 1604 21643 1660
rect 21643 1604 21699 1660
rect 21699 1604 21703 1660
rect 21639 1600 21703 1604
rect 21719 1660 21783 1664
rect 21719 1604 21723 1660
rect 21723 1604 21779 1660
rect 21779 1604 21783 1660
rect 21719 1600 21783 1604
rect 21799 1660 21863 1664
rect 21799 1604 21803 1660
rect 21803 1604 21859 1660
rect 21859 1604 21863 1660
rect 21799 1600 21863 1604
rect 6104 1116 6168 1120
rect 6104 1060 6108 1116
rect 6108 1060 6164 1116
rect 6164 1060 6168 1116
rect 6104 1056 6168 1060
rect 6184 1116 6248 1120
rect 6184 1060 6188 1116
rect 6188 1060 6244 1116
rect 6244 1060 6248 1116
rect 6184 1056 6248 1060
rect 6264 1116 6328 1120
rect 6264 1060 6268 1116
rect 6268 1060 6324 1116
rect 6324 1060 6328 1116
rect 6264 1056 6328 1060
rect 6344 1116 6408 1120
rect 6344 1060 6348 1116
rect 6348 1060 6404 1116
rect 6404 1060 6408 1116
rect 6344 1056 6408 1060
rect 16407 1116 16471 1120
rect 16407 1060 16411 1116
rect 16411 1060 16467 1116
rect 16467 1060 16471 1116
rect 16407 1056 16471 1060
rect 16487 1116 16551 1120
rect 16487 1060 16491 1116
rect 16491 1060 16547 1116
rect 16547 1060 16551 1116
rect 16487 1056 16551 1060
rect 16567 1116 16631 1120
rect 16567 1060 16571 1116
rect 16571 1060 16627 1116
rect 16627 1060 16631 1116
rect 16567 1056 16631 1060
rect 16647 1116 16711 1120
rect 16647 1060 16651 1116
rect 16651 1060 16707 1116
rect 16707 1060 16711 1116
rect 16647 1056 16711 1060
rect 26711 1116 26775 1120
rect 26711 1060 26715 1116
rect 26715 1060 26771 1116
rect 26771 1060 26775 1116
rect 26711 1056 26775 1060
rect 26791 1116 26855 1120
rect 26791 1060 26795 1116
rect 26795 1060 26851 1116
rect 26851 1060 26855 1116
rect 26791 1056 26855 1060
rect 26871 1116 26935 1120
rect 26871 1060 26875 1116
rect 26875 1060 26931 1116
rect 26931 1060 26935 1116
rect 26871 1056 26935 1060
rect 26951 1116 27015 1120
rect 26951 1060 26955 1116
rect 26955 1060 27011 1116
rect 27011 1060 27015 1116
rect 26951 1056 27015 1060
rect 11255 572 11319 576
rect 11255 516 11259 572
rect 11259 516 11315 572
rect 11315 516 11319 572
rect 11255 512 11319 516
rect 11335 572 11399 576
rect 11335 516 11339 572
rect 11339 516 11395 572
rect 11395 516 11399 572
rect 11335 512 11399 516
rect 11415 572 11479 576
rect 11415 516 11419 572
rect 11419 516 11475 572
rect 11475 516 11479 572
rect 11415 512 11479 516
rect 11495 572 11559 576
rect 11495 516 11499 572
rect 11499 516 11555 572
rect 11555 516 11559 572
rect 11495 512 11559 516
rect 21559 572 21623 576
rect 21559 516 21563 572
rect 21563 516 21619 572
rect 21619 516 21623 572
rect 21559 512 21623 516
rect 21639 572 21703 576
rect 21639 516 21643 572
rect 21643 516 21699 572
rect 21699 516 21703 572
rect 21639 512 21703 516
rect 21719 572 21783 576
rect 21719 516 21723 572
rect 21723 516 21779 572
rect 21779 516 21783 572
rect 21719 512 21783 516
rect 21799 572 21863 576
rect 21799 516 21803 572
rect 21803 516 21859 572
rect 21859 516 21863 572
rect 21799 512 21863 516
<< metal4 >>
rect 6095 47904 6416 48464
rect 6095 47840 6104 47904
rect 6168 47840 6184 47904
rect 6248 47840 6264 47904
rect 6328 47840 6344 47904
rect 6408 47840 6416 47904
rect 6095 46816 6416 47840
rect 6095 46752 6104 46816
rect 6168 46752 6184 46816
rect 6248 46752 6264 46816
rect 6328 46752 6344 46816
rect 6408 46752 6416 46816
rect 6095 45728 6416 46752
rect 6095 45664 6104 45728
rect 6168 45664 6184 45728
rect 6248 45664 6264 45728
rect 6328 45664 6344 45728
rect 6408 45664 6416 45728
rect 6095 44640 6416 45664
rect 6095 44576 6104 44640
rect 6168 44576 6184 44640
rect 6248 44576 6264 44640
rect 6328 44576 6344 44640
rect 6408 44576 6416 44640
rect 6095 43552 6416 44576
rect 6095 43488 6104 43552
rect 6168 43488 6184 43552
rect 6248 43488 6264 43552
rect 6328 43488 6344 43552
rect 6408 43488 6416 43552
rect 6095 42464 6416 43488
rect 6095 42400 6104 42464
rect 6168 42400 6184 42464
rect 6248 42400 6264 42464
rect 6328 42400 6344 42464
rect 6408 42400 6416 42464
rect 6095 41376 6416 42400
rect 6095 41312 6104 41376
rect 6168 41312 6184 41376
rect 6248 41312 6264 41376
rect 6328 41312 6344 41376
rect 6408 41312 6416 41376
rect 6095 40288 6416 41312
rect 6095 40224 6104 40288
rect 6168 40224 6184 40288
rect 6248 40224 6264 40288
rect 6328 40224 6344 40288
rect 6408 40224 6416 40288
rect 6095 39200 6416 40224
rect 6095 39136 6104 39200
rect 6168 39136 6184 39200
rect 6248 39136 6264 39200
rect 6328 39136 6344 39200
rect 6408 39136 6416 39200
rect 6095 38112 6416 39136
rect 6095 38048 6104 38112
rect 6168 38048 6184 38112
rect 6248 38048 6264 38112
rect 6328 38048 6344 38112
rect 6408 38048 6416 38112
rect 6095 37024 6416 38048
rect 6095 36960 6104 37024
rect 6168 36960 6184 37024
rect 6248 36960 6264 37024
rect 6328 36960 6344 37024
rect 6408 36960 6416 37024
rect 6095 35936 6416 36960
rect 6095 35872 6104 35936
rect 6168 35872 6184 35936
rect 6248 35872 6264 35936
rect 6328 35872 6344 35936
rect 6408 35872 6416 35936
rect 6095 34848 6416 35872
rect 6095 34784 6104 34848
rect 6168 34784 6184 34848
rect 6248 34784 6264 34848
rect 6328 34784 6344 34848
rect 6408 34784 6416 34848
rect 6095 33760 6416 34784
rect 6095 33696 6104 33760
rect 6168 33696 6184 33760
rect 6248 33696 6264 33760
rect 6328 33696 6344 33760
rect 6408 33696 6416 33760
rect 6095 32672 6416 33696
rect 6095 32608 6104 32672
rect 6168 32608 6184 32672
rect 6248 32608 6264 32672
rect 6328 32608 6344 32672
rect 6408 32608 6416 32672
rect 6095 31584 6416 32608
rect 6095 31520 6104 31584
rect 6168 31520 6184 31584
rect 6248 31520 6264 31584
rect 6328 31520 6344 31584
rect 6408 31520 6416 31584
rect 6095 30496 6416 31520
rect 6095 30432 6104 30496
rect 6168 30432 6184 30496
rect 6248 30432 6264 30496
rect 6328 30432 6344 30496
rect 6408 30432 6416 30496
rect 6095 29408 6416 30432
rect 6095 29344 6104 29408
rect 6168 29344 6184 29408
rect 6248 29344 6264 29408
rect 6328 29344 6344 29408
rect 6408 29344 6416 29408
rect 6095 28320 6416 29344
rect 6095 28256 6104 28320
rect 6168 28256 6184 28320
rect 6248 28256 6264 28320
rect 6328 28256 6344 28320
rect 6408 28256 6416 28320
rect 6095 27232 6416 28256
rect 6095 27168 6104 27232
rect 6168 27168 6184 27232
rect 6248 27168 6264 27232
rect 6328 27168 6344 27232
rect 6408 27168 6416 27232
rect 6095 26144 6416 27168
rect 6095 26080 6104 26144
rect 6168 26080 6184 26144
rect 6248 26080 6264 26144
rect 6328 26080 6344 26144
rect 6408 26080 6416 26144
rect 6095 25056 6416 26080
rect 6095 24992 6104 25056
rect 6168 24992 6184 25056
rect 6248 24992 6264 25056
rect 6328 24992 6344 25056
rect 6408 24992 6416 25056
rect 6095 23968 6416 24992
rect 6095 23904 6104 23968
rect 6168 23904 6184 23968
rect 6248 23904 6264 23968
rect 6328 23904 6344 23968
rect 6408 23904 6416 23968
rect 6095 22880 6416 23904
rect 6095 22816 6104 22880
rect 6168 22816 6184 22880
rect 6248 22816 6264 22880
rect 6328 22816 6344 22880
rect 6408 22816 6416 22880
rect 6095 21792 6416 22816
rect 6095 21728 6104 21792
rect 6168 21728 6184 21792
rect 6248 21728 6264 21792
rect 6328 21728 6344 21792
rect 6408 21728 6416 21792
rect 6095 20704 6416 21728
rect 6095 20640 6104 20704
rect 6168 20640 6184 20704
rect 6248 20640 6264 20704
rect 6328 20640 6344 20704
rect 6408 20640 6416 20704
rect 6095 19616 6416 20640
rect 6095 19552 6104 19616
rect 6168 19552 6184 19616
rect 6248 19552 6264 19616
rect 6328 19552 6344 19616
rect 6408 19552 6416 19616
rect 6095 18528 6416 19552
rect 6095 18464 6104 18528
rect 6168 18464 6184 18528
rect 6248 18464 6264 18528
rect 6328 18464 6344 18528
rect 6408 18464 6416 18528
rect 6095 17440 6416 18464
rect 6095 17376 6104 17440
rect 6168 17376 6184 17440
rect 6248 17376 6264 17440
rect 6328 17376 6344 17440
rect 6408 17376 6416 17440
rect 6095 16352 6416 17376
rect 6095 16288 6104 16352
rect 6168 16288 6184 16352
rect 6248 16288 6264 16352
rect 6328 16288 6344 16352
rect 6408 16288 6416 16352
rect 6095 15264 6416 16288
rect 6095 15200 6104 15264
rect 6168 15200 6184 15264
rect 6248 15200 6264 15264
rect 6328 15200 6344 15264
rect 6408 15200 6416 15264
rect 6095 14176 6416 15200
rect 6095 14112 6104 14176
rect 6168 14112 6184 14176
rect 6248 14112 6264 14176
rect 6328 14112 6344 14176
rect 6408 14112 6416 14176
rect 6095 13088 6416 14112
rect 6095 13024 6104 13088
rect 6168 13024 6184 13088
rect 6248 13024 6264 13088
rect 6328 13024 6344 13088
rect 6408 13024 6416 13088
rect 6095 12000 6416 13024
rect 6095 11936 6104 12000
rect 6168 11936 6184 12000
rect 6248 11936 6264 12000
rect 6328 11936 6344 12000
rect 6408 11936 6416 12000
rect 6095 10912 6416 11936
rect 6095 10848 6104 10912
rect 6168 10848 6184 10912
rect 6248 10848 6264 10912
rect 6328 10848 6344 10912
rect 6408 10848 6416 10912
rect 6095 9824 6416 10848
rect 6095 9760 6104 9824
rect 6168 9760 6184 9824
rect 6248 9760 6264 9824
rect 6328 9760 6344 9824
rect 6408 9760 6416 9824
rect 6095 8736 6416 9760
rect 6095 8672 6104 8736
rect 6168 8672 6184 8736
rect 6248 8672 6264 8736
rect 6328 8672 6344 8736
rect 6408 8672 6416 8736
rect 6095 7648 6416 8672
rect 6095 7584 6104 7648
rect 6168 7584 6184 7648
rect 6248 7584 6264 7648
rect 6328 7584 6344 7648
rect 6408 7584 6416 7648
rect 6095 6560 6416 7584
rect 6095 6496 6104 6560
rect 6168 6496 6184 6560
rect 6248 6496 6264 6560
rect 6328 6496 6344 6560
rect 6408 6496 6416 6560
rect 6095 5472 6416 6496
rect 6095 5408 6104 5472
rect 6168 5408 6184 5472
rect 6248 5408 6264 5472
rect 6328 5408 6344 5472
rect 6408 5408 6416 5472
rect 6095 4384 6416 5408
rect 6095 4320 6104 4384
rect 6168 4320 6184 4384
rect 6248 4320 6264 4384
rect 6328 4320 6344 4384
rect 6408 4320 6416 4384
rect 6095 3296 6416 4320
rect 6095 3232 6104 3296
rect 6168 3232 6184 3296
rect 6248 3232 6264 3296
rect 6328 3232 6344 3296
rect 6408 3232 6416 3296
rect 6095 2208 6416 3232
rect 6095 2144 6104 2208
rect 6168 2144 6184 2208
rect 6248 2144 6264 2208
rect 6328 2144 6344 2208
rect 6408 2144 6416 2208
rect 6095 1120 6416 2144
rect 6095 1056 6104 1120
rect 6168 1056 6184 1120
rect 6248 1056 6264 1120
rect 6328 1056 6344 1120
rect 6408 1056 6416 1120
rect 6095 496 6416 1056
rect 11247 48448 11567 48464
rect 11247 48384 11255 48448
rect 11319 48384 11335 48448
rect 11399 48384 11415 48448
rect 11479 48384 11495 48448
rect 11559 48384 11567 48448
rect 11247 47360 11567 48384
rect 11247 47296 11255 47360
rect 11319 47296 11335 47360
rect 11399 47296 11415 47360
rect 11479 47296 11495 47360
rect 11559 47296 11567 47360
rect 11247 46272 11567 47296
rect 11247 46208 11255 46272
rect 11319 46208 11335 46272
rect 11399 46208 11415 46272
rect 11479 46208 11495 46272
rect 11559 46208 11567 46272
rect 11247 45184 11567 46208
rect 11247 45120 11255 45184
rect 11319 45120 11335 45184
rect 11399 45120 11415 45184
rect 11479 45120 11495 45184
rect 11559 45120 11567 45184
rect 11247 44096 11567 45120
rect 11247 44032 11255 44096
rect 11319 44032 11335 44096
rect 11399 44032 11415 44096
rect 11479 44032 11495 44096
rect 11559 44032 11567 44096
rect 11247 43008 11567 44032
rect 11247 42944 11255 43008
rect 11319 42944 11335 43008
rect 11399 42944 11415 43008
rect 11479 42944 11495 43008
rect 11559 42944 11567 43008
rect 11247 41920 11567 42944
rect 11247 41856 11255 41920
rect 11319 41856 11335 41920
rect 11399 41856 11415 41920
rect 11479 41856 11495 41920
rect 11559 41856 11567 41920
rect 11247 40832 11567 41856
rect 11247 40768 11255 40832
rect 11319 40768 11335 40832
rect 11399 40768 11415 40832
rect 11479 40768 11495 40832
rect 11559 40768 11567 40832
rect 11247 39744 11567 40768
rect 11247 39680 11255 39744
rect 11319 39680 11335 39744
rect 11399 39680 11415 39744
rect 11479 39680 11495 39744
rect 11559 39680 11567 39744
rect 11247 38656 11567 39680
rect 11247 38592 11255 38656
rect 11319 38592 11335 38656
rect 11399 38592 11415 38656
rect 11479 38592 11495 38656
rect 11559 38592 11567 38656
rect 11247 37568 11567 38592
rect 11247 37504 11255 37568
rect 11319 37504 11335 37568
rect 11399 37504 11415 37568
rect 11479 37504 11495 37568
rect 11559 37504 11567 37568
rect 11247 36480 11567 37504
rect 11247 36416 11255 36480
rect 11319 36416 11335 36480
rect 11399 36416 11415 36480
rect 11479 36416 11495 36480
rect 11559 36416 11567 36480
rect 11247 35392 11567 36416
rect 11247 35328 11255 35392
rect 11319 35328 11335 35392
rect 11399 35328 11415 35392
rect 11479 35328 11495 35392
rect 11559 35328 11567 35392
rect 11247 34304 11567 35328
rect 11247 34240 11255 34304
rect 11319 34240 11335 34304
rect 11399 34240 11415 34304
rect 11479 34240 11495 34304
rect 11559 34240 11567 34304
rect 11247 33216 11567 34240
rect 11247 33152 11255 33216
rect 11319 33152 11335 33216
rect 11399 33152 11415 33216
rect 11479 33152 11495 33216
rect 11559 33152 11567 33216
rect 11247 32128 11567 33152
rect 11247 32064 11255 32128
rect 11319 32064 11335 32128
rect 11399 32064 11415 32128
rect 11479 32064 11495 32128
rect 11559 32064 11567 32128
rect 11247 31040 11567 32064
rect 11247 30976 11255 31040
rect 11319 30976 11335 31040
rect 11399 30976 11415 31040
rect 11479 30976 11495 31040
rect 11559 30976 11567 31040
rect 11247 29952 11567 30976
rect 11247 29888 11255 29952
rect 11319 29888 11335 29952
rect 11399 29888 11415 29952
rect 11479 29888 11495 29952
rect 11559 29888 11567 29952
rect 11247 28864 11567 29888
rect 11247 28800 11255 28864
rect 11319 28800 11335 28864
rect 11399 28800 11415 28864
rect 11479 28800 11495 28864
rect 11559 28800 11567 28864
rect 11247 27776 11567 28800
rect 11247 27712 11255 27776
rect 11319 27712 11335 27776
rect 11399 27712 11415 27776
rect 11479 27712 11495 27776
rect 11559 27712 11567 27776
rect 11247 26688 11567 27712
rect 11247 26624 11255 26688
rect 11319 26624 11335 26688
rect 11399 26624 11415 26688
rect 11479 26624 11495 26688
rect 11559 26624 11567 26688
rect 11247 25600 11567 26624
rect 11247 25536 11255 25600
rect 11319 25536 11335 25600
rect 11399 25536 11415 25600
rect 11479 25536 11495 25600
rect 11559 25536 11567 25600
rect 11247 24512 11567 25536
rect 11247 24448 11255 24512
rect 11319 24448 11335 24512
rect 11399 24448 11415 24512
rect 11479 24448 11495 24512
rect 11559 24448 11567 24512
rect 11247 23424 11567 24448
rect 11247 23360 11255 23424
rect 11319 23360 11335 23424
rect 11399 23360 11415 23424
rect 11479 23360 11495 23424
rect 11559 23360 11567 23424
rect 11247 22336 11567 23360
rect 11247 22272 11255 22336
rect 11319 22272 11335 22336
rect 11399 22272 11415 22336
rect 11479 22272 11495 22336
rect 11559 22272 11567 22336
rect 11247 21248 11567 22272
rect 11247 21184 11255 21248
rect 11319 21184 11335 21248
rect 11399 21184 11415 21248
rect 11479 21184 11495 21248
rect 11559 21184 11567 21248
rect 11247 20160 11567 21184
rect 11247 20096 11255 20160
rect 11319 20096 11335 20160
rect 11399 20096 11415 20160
rect 11479 20096 11495 20160
rect 11559 20096 11567 20160
rect 11247 19072 11567 20096
rect 11247 19008 11255 19072
rect 11319 19008 11335 19072
rect 11399 19008 11415 19072
rect 11479 19008 11495 19072
rect 11559 19008 11567 19072
rect 11247 17984 11567 19008
rect 11247 17920 11255 17984
rect 11319 17920 11335 17984
rect 11399 17920 11415 17984
rect 11479 17920 11495 17984
rect 11559 17920 11567 17984
rect 11247 16896 11567 17920
rect 11247 16832 11255 16896
rect 11319 16832 11335 16896
rect 11399 16832 11415 16896
rect 11479 16832 11495 16896
rect 11559 16832 11567 16896
rect 11247 15808 11567 16832
rect 11247 15744 11255 15808
rect 11319 15744 11335 15808
rect 11399 15744 11415 15808
rect 11479 15744 11495 15808
rect 11559 15744 11567 15808
rect 11247 14720 11567 15744
rect 11247 14656 11255 14720
rect 11319 14656 11335 14720
rect 11399 14656 11415 14720
rect 11479 14656 11495 14720
rect 11559 14656 11567 14720
rect 11247 13632 11567 14656
rect 11247 13568 11255 13632
rect 11319 13568 11335 13632
rect 11399 13568 11415 13632
rect 11479 13568 11495 13632
rect 11559 13568 11567 13632
rect 11247 12544 11567 13568
rect 11247 12480 11255 12544
rect 11319 12480 11335 12544
rect 11399 12480 11415 12544
rect 11479 12480 11495 12544
rect 11559 12480 11567 12544
rect 11247 11456 11567 12480
rect 11247 11392 11255 11456
rect 11319 11392 11335 11456
rect 11399 11392 11415 11456
rect 11479 11392 11495 11456
rect 11559 11392 11567 11456
rect 11247 10368 11567 11392
rect 11247 10304 11255 10368
rect 11319 10304 11335 10368
rect 11399 10304 11415 10368
rect 11479 10304 11495 10368
rect 11559 10304 11567 10368
rect 11247 9280 11567 10304
rect 11247 9216 11255 9280
rect 11319 9216 11335 9280
rect 11399 9216 11415 9280
rect 11479 9216 11495 9280
rect 11559 9216 11567 9280
rect 11247 8192 11567 9216
rect 11247 8128 11255 8192
rect 11319 8128 11335 8192
rect 11399 8128 11415 8192
rect 11479 8128 11495 8192
rect 11559 8128 11567 8192
rect 11247 7104 11567 8128
rect 11247 7040 11255 7104
rect 11319 7040 11335 7104
rect 11399 7040 11415 7104
rect 11479 7040 11495 7104
rect 11559 7040 11567 7104
rect 11247 6016 11567 7040
rect 11247 5952 11255 6016
rect 11319 5952 11335 6016
rect 11399 5952 11415 6016
rect 11479 5952 11495 6016
rect 11559 5952 11567 6016
rect 11247 4928 11567 5952
rect 11247 4864 11255 4928
rect 11319 4864 11335 4928
rect 11399 4864 11415 4928
rect 11479 4864 11495 4928
rect 11559 4864 11567 4928
rect 11247 3840 11567 4864
rect 11247 3776 11255 3840
rect 11319 3776 11335 3840
rect 11399 3776 11415 3840
rect 11479 3776 11495 3840
rect 11559 3776 11567 3840
rect 11247 2752 11567 3776
rect 11247 2688 11255 2752
rect 11319 2688 11335 2752
rect 11399 2688 11415 2752
rect 11479 2688 11495 2752
rect 11559 2688 11567 2752
rect 11247 1664 11567 2688
rect 11247 1600 11255 1664
rect 11319 1600 11335 1664
rect 11399 1600 11415 1664
rect 11479 1600 11495 1664
rect 11559 1600 11567 1664
rect 11247 576 11567 1600
rect 11247 512 11255 576
rect 11319 512 11335 576
rect 11399 512 11415 576
rect 11479 512 11495 576
rect 11559 512 11567 576
rect 11247 496 11567 512
rect 16399 47904 16719 48464
rect 16399 47840 16407 47904
rect 16471 47840 16487 47904
rect 16551 47840 16567 47904
rect 16631 47840 16647 47904
rect 16711 47840 16719 47904
rect 16399 46816 16719 47840
rect 16399 46752 16407 46816
rect 16471 46752 16487 46816
rect 16551 46752 16567 46816
rect 16631 46752 16647 46816
rect 16711 46752 16719 46816
rect 16399 45728 16719 46752
rect 16399 45664 16407 45728
rect 16471 45664 16487 45728
rect 16551 45664 16567 45728
rect 16631 45664 16647 45728
rect 16711 45664 16719 45728
rect 16399 44640 16719 45664
rect 16399 44576 16407 44640
rect 16471 44576 16487 44640
rect 16551 44576 16567 44640
rect 16631 44576 16647 44640
rect 16711 44576 16719 44640
rect 16399 43552 16719 44576
rect 16399 43488 16407 43552
rect 16471 43488 16487 43552
rect 16551 43488 16567 43552
rect 16631 43488 16647 43552
rect 16711 43488 16719 43552
rect 16399 42464 16719 43488
rect 16399 42400 16407 42464
rect 16471 42400 16487 42464
rect 16551 42400 16567 42464
rect 16631 42400 16647 42464
rect 16711 42400 16719 42464
rect 16399 41376 16719 42400
rect 16399 41312 16407 41376
rect 16471 41312 16487 41376
rect 16551 41312 16567 41376
rect 16631 41312 16647 41376
rect 16711 41312 16719 41376
rect 16399 40288 16719 41312
rect 16399 40224 16407 40288
rect 16471 40224 16487 40288
rect 16551 40224 16567 40288
rect 16631 40224 16647 40288
rect 16711 40224 16719 40288
rect 16399 39200 16719 40224
rect 16399 39136 16407 39200
rect 16471 39136 16487 39200
rect 16551 39136 16567 39200
rect 16631 39136 16647 39200
rect 16711 39136 16719 39200
rect 16399 38112 16719 39136
rect 16399 38048 16407 38112
rect 16471 38048 16487 38112
rect 16551 38048 16567 38112
rect 16631 38048 16647 38112
rect 16711 38048 16719 38112
rect 16399 37024 16719 38048
rect 16399 36960 16407 37024
rect 16471 36960 16487 37024
rect 16551 36960 16567 37024
rect 16631 36960 16647 37024
rect 16711 36960 16719 37024
rect 16399 35936 16719 36960
rect 16399 35872 16407 35936
rect 16471 35872 16487 35936
rect 16551 35872 16567 35936
rect 16631 35872 16647 35936
rect 16711 35872 16719 35936
rect 16399 34848 16719 35872
rect 16399 34784 16407 34848
rect 16471 34784 16487 34848
rect 16551 34784 16567 34848
rect 16631 34784 16647 34848
rect 16711 34784 16719 34848
rect 16399 33760 16719 34784
rect 16399 33696 16407 33760
rect 16471 33696 16487 33760
rect 16551 33696 16567 33760
rect 16631 33696 16647 33760
rect 16711 33696 16719 33760
rect 16399 32672 16719 33696
rect 16399 32608 16407 32672
rect 16471 32608 16487 32672
rect 16551 32608 16567 32672
rect 16631 32608 16647 32672
rect 16711 32608 16719 32672
rect 16399 31584 16719 32608
rect 16399 31520 16407 31584
rect 16471 31520 16487 31584
rect 16551 31520 16567 31584
rect 16631 31520 16647 31584
rect 16711 31520 16719 31584
rect 16399 30496 16719 31520
rect 16399 30432 16407 30496
rect 16471 30432 16487 30496
rect 16551 30432 16567 30496
rect 16631 30432 16647 30496
rect 16711 30432 16719 30496
rect 16399 29408 16719 30432
rect 16399 29344 16407 29408
rect 16471 29344 16487 29408
rect 16551 29344 16567 29408
rect 16631 29344 16647 29408
rect 16711 29344 16719 29408
rect 16399 28320 16719 29344
rect 16399 28256 16407 28320
rect 16471 28256 16487 28320
rect 16551 28256 16567 28320
rect 16631 28256 16647 28320
rect 16711 28256 16719 28320
rect 16399 27232 16719 28256
rect 16399 27168 16407 27232
rect 16471 27168 16487 27232
rect 16551 27168 16567 27232
rect 16631 27168 16647 27232
rect 16711 27168 16719 27232
rect 16399 26144 16719 27168
rect 16399 26080 16407 26144
rect 16471 26080 16487 26144
rect 16551 26080 16567 26144
rect 16631 26080 16647 26144
rect 16711 26080 16719 26144
rect 16399 25056 16719 26080
rect 16399 24992 16407 25056
rect 16471 24992 16487 25056
rect 16551 24992 16567 25056
rect 16631 24992 16647 25056
rect 16711 24992 16719 25056
rect 16399 23968 16719 24992
rect 16399 23904 16407 23968
rect 16471 23904 16487 23968
rect 16551 23904 16567 23968
rect 16631 23904 16647 23968
rect 16711 23904 16719 23968
rect 16399 22880 16719 23904
rect 16399 22816 16407 22880
rect 16471 22816 16487 22880
rect 16551 22816 16567 22880
rect 16631 22816 16647 22880
rect 16711 22816 16719 22880
rect 16399 21792 16719 22816
rect 16399 21728 16407 21792
rect 16471 21728 16487 21792
rect 16551 21728 16567 21792
rect 16631 21728 16647 21792
rect 16711 21728 16719 21792
rect 16399 20704 16719 21728
rect 16399 20640 16407 20704
rect 16471 20640 16487 20704
rect 16551 20640 16567 20704
rect 16631 20640 16647 20704
rect 16711 20640 16719 20704
rect 16399 19616 16719 20640
rect 16399 19552 16407 19616
rect 16471 19552 16487 19616
rect 16551 19552 16567 19616
rect 16631 19552 16647 19616
rect 16711 19552 16719 19616
rect 16399 18528 16719 19552
rect 16399 18464 16407 18528
rect 16471 18464 16487 18528
rect 16551 18464 16567 18528
rect 16631 18464 16647 18528
rect 16711 18464 16719 18528
rect 16399 17440 16719 18464
rect 16399 17376 16407 17440
rect 16471 17376 16487 17440
rect 16551 17376 16567 17440
rect 16631 17376 16647 17440
rect 16711 17376 16719 17440
rect 16399 16352 16719 17376
rect 16399 16288 16407 16352
rect 16471 16288 16487 16352
rect 16551 16288 16567 16352
rect 16631 16288 16647 16352
rect 16711 16288 16719 16352
rect 16399 15264 16719 16288
rect 16399 15200 16407 15264
rect 16471 15200 16487 15264
rect 16551 15200 16567 15264
rect 16631 15200 16647 15264
rect 16711 15200 16719 15264
rect 16399 14176 16719 15200
rect 16399 14112 16407 14176
rect 16471 14112 16487 14176
rect 16551 14112 16567 14176
rect 16631 14112 16647 14176
rect 16711 14112 16719 14176
rect 16399 13088 16719 14112
rect 16399 13024 16407 13088
rect 16471 13024 16487 13088
rect 16551 13024 16567 13088
rect 16631 13024 16647 13088
rect 16711 13024 16719 13088
rect 16399 12000 16719 13024
rect 16399 11936 16407 12000
rect 16471 11936 16487 12000
rect 16551 11936 16567 12000
rect 16631 11936 16647 12000
rect 16711 11936 16719 12000
rect 16399 10912 16719 11936
rect 16399 10848 16407 10912
rect 16471 10848 16487 10912
rect 16551 10848 16567 10912
rect 16631 10848 16647 10912
rect 16711 10848 16719 10912
rect 16399 9824 16719 10848
rect 16399 9760 16407 9824
rect 16471 9760 16487 9824
rect 16551 9760 16567 9824
rect 16631 9760 16647 9824
rect 16711 9760 16719 9824
rect 16399 8736 16719 9760
rect 16399 8672 16407 8736
rect 16471 8672 16487 8736
rect 16551 8672 16567 8736
rect 16631 8672 16647 8736
rect 16711 8672 16719 8736
rect 16399 7648 16719 8672
rect 16399 7584 16407 7648
rect 16471 7584 16487 7648
rect 16551 7584 16567 7648
rect 16631 7584 16647 7648
rect 16711 7584 16719 7648
rect 16399 6560 16719 7584
rect 16399 6496 16407 6560
rect 16471 6496 16487 6560
rect 16551 6496 16567 6560
rect 16631 6496 16647 6560
rect 16711 6496 16719 6560
rect 16399 5472 16719 6496
rect 16399 5408 16407 5472
rect 16471 5408 16487 5472
rect 16551 5408 16567 5472
rect 16631 5408 16647 5472
rect 16711 5408 16719 5472
rect 16399 4384 16719 5408
rect 16399 4320 16407 4384
rect 16471 4320 16487 4384
rect 16551 4320 16567 4384
rect 16631 4320 16647 4384
rect 16711 4320 16719 4384
rect 16399 3296 16719 4320
rect 16399 3232 16407 3296
rect 16471 3232 16487 3296
rect 16551 3232 16567 3296
rect 16631 3232 16647 3296
rect 16711 3232 16719 3296
rect 16399 2208 16719 3232
rect 16399 2144 16407 2208
rect 16471 2144 16487 2208
rect 16551 2144 16567 2208
rect 16631 2144 16647 2208
rect 16711 2144 16719 2208
rect 16399 1120 16719 2144
rect 16399 1056 16407 1120
rect 16471 1056 16487 1120
rect 16551 1056 16567 1120
rect 16631 1056 16647 1120
rect 16711 1056 16719 1120
rect 16399 496 16719 1056
rect 21551 48448 21871 48464
rect 21551 48384 21559 48448
rect 21623 48384 21639 48448
rect 21703 48384 21719 48448
rect 21783 48384 21799 48448
rect 21863 48384 21871 48448
rect 21551 47360 21871 48384
rect 21551 47296 21559 47360
rect 21623 47296 21639 47360
rect 21703 47296 21719 47360
rect 21783 47296 21799 47360
rect 21863 47296 21871 47360
rect 21551 46272 21871 47296
rect 21551 46208 21559 46272
rect 21623 46208 21639 46272
rect 21703 46208 21719 46272
rect 21783 46208 21799 46272
rect 21863 46208 21871 46272
rect 21551 45184 21871 46208
rect 21551 45120 21559 45184
rect 21623 45120 21639 45184
rect 21703 45120 21719 45184
rect 21783 45120 21799 45184
rect 21863 45120 21871 45184
rect 21551 44096 21871 45120
rect 21551 44032 21559 44096
rect 21623 44032 21639 44096
rect 21703 44032 21719 44096
rect 21783 44032 21799 44096
rect 21863 44032 21871 44096
rect 21551 43008 21871 44032
rect 21551 42944 21559 43008
rect 21623 42944 21639 43008
rect 21703 42944 21719 43008
rect 21783 42944 21799 43008
rect 21863 42944 21871 43008
rect 21551 41920 21871 42944
rect 21551 41856 21559 41920
rect 21623 41856 21639 41920
rect 21703 41856 21719 41920
rect 21783 41856 21799 41920
rect 21863 41856 21871 41920
rect 21551 40832 21871 41856
rect 21551 40768 21559 40832
rect 21623 40768 21639 40832
rect 21703 40768 21719 40832
rect 21783 40768 21799 40832
rect 21863 40768 21871 40832
rect 21551 39744 21871 40768
rect 21551 39680 21559 39744
rect 21623 39680 21639 39744
rect 21703 39680 21719 39744
rect 21783 39680 21799 39744
rect 21863 39680 21871 39744
rect 21551 38656 21871 39680
rect 21551 38592 21559 38656
rect 21623 38592 21639 38656
rect 21703 38592 21719 38656
rect 21783 38592 21799 38656
rect 21863 38592 21871 38656
rect 21551 37568 21871 38592
rect 21551 37504 21559 37568
rect 21623 37504 21639 37568
rect 21703 37504 21719 37568
rect 21783 37504 21799 37568
rect 21863 37504 21871 37568
rect 21551 36480 21871 37504
rect 21551 36416 21559 36480
rect 21623 36416 21639 36480
rect 21703 36416 21719 36480
rect 21783 36416 21799 36480
rect 21863 36416 21871 36480
rect 21551 35392 21871 36416
rect 21551 35328 21559 35392
rect 21623 35328 21639 35392
rect 21703 35328 21719 35392
rect 21783 35328 21799 35392
rect 21863 35328 21871 35392
rect 21551 34304 21871 35328
rect 21551 34240 21559 34304
rect 21623 34240 21639 34304
rect 21703 34240 21719 34304
rect 21783 34240 21799 34304
rect 21863 34240 21871 34304
rect 21551 33216 21871 34240
rect 21551 33152 21559 33216
rect 21623 33152 21639 33216
rect 21703 33152 21719 33216
rect 21783 33152 21799 33216
rect 21863 33152 21871 33216
rect 21551 32128 21871 33152
rect 21551 32064 21559 32128
rect 21623 32064 21639 32128
rect 21703 32064 21719 32128
rect 21783 32064 21799 32128
rect 21863 32064 21871 32128
rect 21551 31040 21871 32064
rect 21551 30976 21559 31040
rect 21623 30976 21639 31040
rect 21703 30976 21719 31040
rect 21783 30976 21799 31040
rect 21863 30976 21871 31040
rect 21551 29952 21871 30976
rect 21551 29888 21559 29952
rect 21623 29888 21639 29952
rect 21703 29888 21719 29952
rect 21783 29888 21799 29952
rect 21863 29888 21871 29952
rect 21551 28864 21871 29888
rect 21551 28800 21559 28864
rect 21623 28800 21639 28864
rect 21703 28800 21719 28864
rect 21783 28800 21799 28864
rect 21863 28800 21871 28864
rect 21551 27776 21871 28800
rect 21551 27712 21559 27776
rect 21623 27712 21639 27776
rect 21703 27712 21719 27776
rect 21783 27712 21799 27776
rect 21863 27712 21871 27776
rect 21551 26688 21871 27712
rect 21551 26624 21559 26688
rect 21623 26624 21639 26688
rect 21703 26624 21719 26688
rect 21783 26624 21799 26688
rect 21863 26624 21871 26688
rect 21551 25600 21871 26624
rect 21551 25536 21559 25600
rect 21623 25536 21639 25600
rect 21703 25536 21719 25600
rect 21783 25536 21799 25600
rect 21863 25536 21871 25600
rect 21551 24512 21871 25536
rect 21551 24448 21559 24512
rect 21623 24448 21639 24512
rect 21703 24448 21719 24512
rect 21783 24448 21799 24512
rect 21863 24448 21871 24512
rect 21551 23424 21871 24448
rect 21551 23360 21559 23424
rect 21623 23360 21639 23424
rect 21703 23360 21719 23424
rect 21783 23360 21799 23424
rect 21863 23360 21871 23424
rect 21551 22336 21871 23360
rect 21551 22272 21559 22336
rect 21623 22272 21639 22336
rect 21703 22272 21719 22336
rect 21783 22272 21799 22336
rect 21863 22272 21871 22336
rect 21551 21248 21871 22272
rect 21551 21184 21559 21248
rect 21623 21184 21639 21248
rect 21703 21184 21719 21248
rect 21783 21184 21799 21248
rect 21863 21184 21871 21248
rect 21551 20160 21871 21184
rect 21551 20096 21559 20160
rect 21623 20096 21639 20160
rect 21703 20096 21719 20160
rect 21783 20096 21799 20160
rect 21863 20096 21871 20160
rect 21551 19072 21871 20096
rect 21551 19008 21559 19072
rect 21623 19008 21639 19072
rect 21703 19008 21719 19072
rect 21783 19008 21799 19072
rect 21863 19008 21871 19072
rect 21551 17984 21871 19008
rect 21551 17920 21559 17984
rect 21623 17920 21639 17984
rect 21703 17920 21719 17984
rect 21783 17920 21799 17984
rect 21863 17920 21871 17984
rect 21551 16896 21871 17920
rect 21551 16832 21559 16896
rect 21623 16832 21639 16896
rect 21703 16832 21719 16896
rect 21783 16832 21799 16896
rect 21863 16832 21871 16896
rect 21551 15808 21871 16832
rect 21551 15744 21559 15808
rect 21623 15744 21639 15808
rect 21703 15744 21719 15808
rect 21783 15744 21799 15808
rect 21863 15744 21871 15808
rect 21551 14720 21871 15744
rect 21551 14656 21559 14720
rect 21623 14656 21639 14720
rect 21703 14656 21719 14720
rect 21783 14656 21799 14720
rect 21863 14656 21871 14720
rect 21551 13632 21871 14656
rect 21551 13568 21559 13632
rect 21623 13568 21639 13632
rect 21703 13568 21719 13632
rect 21783 13568 21799 13632
rect 21863 13568 21871 13632
rect 21551 12544 21871 13568
rect 21551 12480 21559 12544
rect 21623 12480 21639 12544
rect 21703 12480 21719 12544
rect 21783 12480 21799 12544
rect 21863 12480 21871 12544
rect 21551 11456 21871 12480
rect 21551 11392 21559 11456
rect 21623 11392 21639 11456
rect 21703 11392 21719 11456
rect 21783 11392 21799 11456
rect 21863 11392 21871 11456
rect 21551 10368 21871 11392
rect 21551 10304 21559 10368
rect 21623 10304 21639 10368
rect 21703 10304 21719 10368
rect 21783 10304 21799 10368
rect 21863 10304 21871 10368
rect 21551 9280 21871 10304
rect 21551 9216 21559 9280
rect 21623 9216 21639 9280
rect 21703 9216 21719 9280
rect 21783 9216 21799 9280
rect 21863 9216 21871 9280
rect 21551 8192 21871 9216
rect 21551 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21799 8192
rect 21863 8128 21871 8192
rect 21551 7104 21871 8128
rect 21551 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21799 7104
rect 21863 7040 21871 7104
rect 21551 6016 21871 7040
rect 21551 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21799 6016
rect 21863 5952 21871 6016
rect 21551 4928 21871 5952
rect 21551 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21799 4928
rect 21863 4864 21871 4928
rect 21551 3840 21871 4864
rect 21551 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21799 3840
rect 21863 3776 21871 3840
rect 21551 2752 21871 3776
rect 21551 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21799 2752
rect 21863 2688 21871 2752
rect 21551 1664 21871 2688
rect 21551 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21799 1664
rect 21863 1600 21871 1664
rect 21551 576 21871 1600
rect 21551 512 21559 576
rect 21623 512 21639 576
rect 21703 512 21719 576
rect 21783 512 21799 576
rect 21863 512 21871 576
rect 21551 496 21871 512
rect 26703 47904 27023 48464
rect 26703 47840 26711 47904
rect 26775 47840 26791 47904
rect 26855 47840 26871 47904
rect 26935 47840 26951 47904
rect 27015 47840 27023 47904
rect 26703 46816 27023 47840
rect 26703 46752 26711 46816
rect 26775 46752 26791 46816
rect 26855 46752 26871 46816
rect 26935 46752 26951 46816
rect 27015 46752 27023 46816
rect 26703 45728 27023 46752
rect 26703 45664 26711 45728
rect 26775 45664 26791 45728
rect 26855 45664 26871 45728
rect 26935 45664 26951 45728
rect 27015 45664 27023 45728
rect 26703 44640 27023 45664
rect 26703 44576 26711 44640
rect 26775 44576 26791 44640
rect 26855 44576 26871 44640
rect 26935 44576 26951 44640
rect 27015 44576 27023 44640
rect 26703 43552 27023 44576
rect 26703 43488 26711 43552
rect 26775 43488 26791 43552
rect 26855 43488 26871 43552
rect 26935 43488 26951 43552
rect 27015 43488 27023 43552
rect 26703 42464 27023 43488
rect 26703 42400 26711 42464
rect 26775 42400 26791 42464
rect 26855 42400 26871 42464
rect 26935 42400 26951 42464
rect 27015 42400 27023 42464
rect 26703 41376 27023 42400
rect 26703 41312 26711 41376
rect 26775 41312 26791 41376
rect 26855 41312 26871 41376
rect 26935 41312 26951 41376
rect 27015 41312 27023 41376
rect 26703 40288 27023 41312
rect 26703 40224 26711 40288
rect 26775 40224 26791 40288
rect 26855 40224 26871 40288
rect 26935 40224 26951 40288
rect 27015 40224 27023 40288
rect 26703 39200 27023 40224
rect 26703 39136 26711 39200
rect 26775 39136 26791 39200
rect 26855 39136 26871 39200
rect 26935 39136 26951 39200
rect 27015 39136 27023 39200
rect 26703 38112 27023 39136
rect 26703 38048 26711 38112
rect 26775 38048 26791 38112
rect 26855 38048 26871 38112
rect 26935 38048 26951 38112
rect 27015 38048 27023 38112
rect 26703 37024 27023 38048
rect 26703 36960 26711 37024
rect 26775 36960 26791 37024
rect 26855 36960 26871 37024
rect 26935 36960 26951 37024
rect 27015 36960 27023 37024
rect 26703 35936 27023 36960
rect 26703 35872 26711 35936
rect 26775 35872 26791 35936
rect 26855 35872 26871 35936
rect 26935 35872 26951 35936
rect 27015 35872 27023 35936
rect 26703 34848 27023 35872
rect 26703 34784 26711 34848
rect 26775 34784 26791 34848
rect 26855 34784 26871 34848
rect 26935 34784 26951 34848
rect 27015 34784 27023 34848
rect 26703 33760 27023 34784
rect 26703 33696 26711 33760
rect 26775 33696 26791 33760
rect 26855 33696 26871 33760
rect 26935 33696 26951 33760
rect 27015 33696 27023 33760
rect 26703 32672 27023 33696
rect 26703 32608 26711 32672
rect 26775 32608 26791 32672
rect 26855 32608 26871 32672
rect 26935 32608 26951 32672
rect 27015 32608 27023 32672
rect 26703 31584 27023 32608
rect 26703 31520 26711 31584
rect 26775 31520 26791 31584
rect 26855 31520 26871 31584
rect 26935 31520 26951 31584
rect 27015 31520 27023 31584
rect 26703 30496 27023 31520
rect 26703 30432 26711 30496
rect 26775 30432 26791 30496
rect 26855 30432 26871 30496
rect 26935 30432 26951 30496
rect 27015 30432 27023 30496
rect 26703 29408 27023 30432
rect 26703 29344 26711 29408
rect 26775 29344 26791 29408
rect 26855 29344 26871 29408
rect 26935 29344 26951 29408
rect 27015 29344 27023 29408
rect 26703 28320 27023 29344
rect 26703 28256 26711 28320
rect 26775 28256 26791 28320
rect 26855 28256 26871 28320
rect 26935 28256 26951 28320
rect 27015 28256 27023 28320
rect 26703 27232 27023 28256
rect 26703 27168 26711 27232
rect 26775 27168 26791 27232
rect 26855 27168 26871 27232
rect 26935 27168 26951 27232
rect 27015 27168 27023 27232
rect 26703 26144 27023 27168
rect 26703 26080 26711 26144
rect 26775 26080 26791 26144
rect 26855 26080 26871 26144
rect 26935 26080 26951 26144
rect 27015 26080 27023 26144
rect 26703 25056 27023 26080
rect 26703 24992 26711 25056
rect 26775 24992 26791 25056
rect 26855 24992 26871 25056
rect 26935 24992 26951 25056
rect 27015 24992 27023 25056
rect 26703 23968 27023 24992
rect 26703 23904 26711 23968
rect 26775 23904 26791 23968
rect 26855 23904 26871 23968
rect 26935 23904 26951 23968
rect 27015 23904 27023 23968
rect 26703 22880 27023 23904
rect 26703 22816 26711 22880
rect 26775 22816 26791 22880
rect 26855 22816 26871 22880
rect 26935 22816 26951 22880
rect 27015 22816 27023 22880
rect 26703 21792 27023 22816
rect 26703 21728 26711 21792
rect 26775 21728 26791 21792
rect 26855 21728 26871 21792
rect 26935 21728 26951 21792
rect 27015 21728 27023 21792
rect 26703 20704 27023 21728
rect 26703 20640 26711 20704
rect 26775 20640 26791 20704
rect 26855 20640 26871 20704
rect 26935 20640 26951 20704
rect 27015 20640 27023 20704
rect 26703 19616 27023 20640
rect 26703 19552 26711 19616
rect 26775 19552 26791 19616
rect 26855 19552 26871 19616
rect 26935 19552 26951 19616
rect 27015 19552 27023 19616
rect 26703 18528 27023 19552
rect 26703 18464 26711 18528
rect 26775 18464 26791 18528
rect 26855 18464 26871 18528
rect 26935 18464 26951 18528
rect 27015 18464 27023 18528
rect 26703 17440 27023 18464
rect 26703 17376 26711 17440
rect 26775 17376 26791 17440
rect 26855 17376 26871 17440
rect 26935 17376 26951 17440
rect 27015 17376 27023 17440
rect 26703 16352 27023 17376
rect 26703 16288 26711 16352
rect 26775 16288 26791 16352
rect 26855 16288 26871 16352
rect 26935 16288 26951 16352
rect 27015 16288 27023 16352
rect 26703 15264 27023 16288
rect 26703 15200 26711 15264
rect 26775 15200 26791 15264
rect 26855 15200 26871 15264
rect 26935 15200 26951 15264
rect 27015 15200 27023 15264
rect 26703 14176 27023 15200
rect 26703 14112 26711 14176
rect 26775 14112 26791 14176
rect 26855 14112 26871 14176
rect 26935 14112 26951 14176
rect 27015 14112 27023 14176
rect 26703 13088 27023 14112
rect 26703 13024 26711 13088
rect 26775 13024 26791 13088
rect 26855 13024 26871 13088
rect 26935 13024 26951 13088
rect 27015 13024 27023 13088
rect 26703 12000 27023 13024
rect 26703 11936 26711 12000
rect 26775 11936 26791 12000
rect 26855 11936 26871 12000
rect 26935 11936 26951 12000
rect 27015 11936 27023 12000
rect 26703 10912 27023 11936
rect 26703 10848 26711 10912
rect 26775 10848 26791 10912
rect 26855 10848 26871 10912
rect 26935 10848 26951 10912
rect 27015 10848 27023 10912
rect 26703 9824 27023 10848
rect 26703 9760 26711 9824
rect 26775 9760 26791 9824
rect 26855 9760 26871 9824
rect 26935 9760 26951 9824
rect 27015 9760 27023 9824
rect 26703 8736 27023 9760
rect 26703 8672 26711 8736
rect 26775 8672 26791 8736
rect 26855 8672 26871 8736
rect 26935 8672 26951 8736
rect 27015 8672 27023 8736
rect 26703 7648 27023 8672
rect 26703 7584 26711 7648
rect 26775 7584 26791 7648
rect 26855 7584 26871 7648
rect 26935 7584 26951 7648
rect 27015 7584 27023 7648
rect 26703 6560 27023 7584
rect 26703 6496 26711 6560
rect 26775 6496 26791 6560
rect 26855 6496 26871 6560
rect 26935 6496 26951 6560
rect 27015 6496 27023 6560
rect 26703 5472 27023 6496
rect 26703 5408 26711 5472
rect 26775 5408 26791 5472
rect 26855 5408 26871 5472
rect 26935 5408 26951 5472
rect 27015 5408 27023 5472
rect 26703 4384 27023 5408
rect 26703 4320 26711 4384
rect 26775 4320 26791 4384
rect 26855 4320 26871 4384
rect 26935 4320 26951 4384
rect 27015 4320 27023 4384
rect 26703 3296 27023 4320
rect 26703 3232 26711 3296
rect 26775 3232 26791 3296
rect 26855 3232 26871 3296
rect 26935 3232 26951 3296
rect 27015 3232 27023 3296
rect 26703 2208 27023 3232
rect 26703 2144 26711 2208
rect 26775 2144 26791 2208
rect 26855 2144 26871 2208
rect 26935 2144 26951 2208
rect 27015 2144 27023 2208
rect 26703 1120 27023 2144
rect 26703 1056 26711 1120
rect 26775 1056 26791 1120
rect 26855 1056 26871 1120
rect 26935 1056 26951 1120
rect 27015 1056 27023 1120
rect 26703 496 27023 1056
use sky130_fd_sc_hd__clkbuf_4  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 1748 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1646674385
transform 1 0 1104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 1380 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 1380 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 1748 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1646674385
transform 1 0 2300 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 2852 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1646674385
transform -1 0 2852 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 2852 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_7
timestamp 1646674385
transform 1 0 1748 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 3588 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1646674385
transform 1 0 3772 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1646674385
transform 1 0 4876 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 1646674385
transform 1 0 3956 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 3680 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1646674385
transform 1 0 5980 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1646674385
transform 1 0 6348 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1646674385
transform 1 0 5060 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1646674385
transform 1 0 6164 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1646674385
transform 1 0 6348 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1646674385
transform 1 0 6256 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1646674385
transform 1 0 6256 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1646674385
transform 1 0 7084 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1646674385
transform -1 0 7360 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1646674385
transform 1 0 7452 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1646674385
transform 1 0 7360 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1646674385
transform -1 0 7912 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1646674385
transform 1 0 8096 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1646674385
transform 1 0 7820 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1646674385
transform 1 0 7912 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_prog_clk_A
timestamp 1646674385
transform 1 0 7912 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1646674385
transform 1 0 8464 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_prog_clk_A
timestamp 1646674385
transform -1 0 8464 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_prog_clk_A
timestamp 1646674385
transform 1 0 8464 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1646674385
transform 1 0 8648 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 9292 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1646674385
transform 1 0 8832 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_88
timestamp 1646674385
transform 1 0 9200 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 9660 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1646674385
transform 1 0 8924 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_prog_clk_A
timestamp 1646674385
transform 1 0 9016 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99
timestamp 1646674385
transform 1 0 10212 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1646674385
transform 1 0 10488 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1646674385
transform -1 0 10488 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2625_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 11040 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1646674385
transform 1 0 11408 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1646674385
transform 1 0 11408 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1646674385
transform 1 0 11040 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1646674385
transform 1 0 11500 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1646674385
transform 1 0 11040 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2497__A2
timestamp 1646674385
transform -1 0 11040 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2483__B1
timestamp 1646674385
transform -1 0 11684 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_121
timestamp 1646674385
transform 1 0 12236 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1646674385
transform 1 0 11684 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2482__C
timestamp 1646674385
transform -1 0 12236 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2481__B2
timestamp 1646674385
transform -1 0 12788 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2623_
timestamp 1646674385
transform -1 0 13248 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1646674385
transform 1 0 13248 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144
timestamp 1646674385
transform 1 0 14352 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1646674385
transform 1 0 12788 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1646674385
transform 1 0 13984 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2601_
timestamp 1646674385
transform 1 0 13156 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 14076 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2481__A2
timestamp 1646674385
transform -1 0 15364 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152
timestamp 1646674385
transform 1 0 15088 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_155
timestamp 1646674385
transform 1 0 15364 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1646674385
transform 1 0 16192 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1646674385
transform 1 0 14628 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1646674385
transform 1 0 16192 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1581_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 16192 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2514_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 15916 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1582_
timestamp 1646674385
transform 1 0 16744 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1646674385
transform 1 0 16560 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1646674385
transform 1 0 16560 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1646674385
transform 1 0 16652 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1646674385
transform 1 0 16652 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_186
timestamp 1646674385
transform 1 0 18216 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1646674385
transform 1 0 18124 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1646674385
transform 1 0 17572 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2430__C
timestamp 1646674385
transform -1 0 18124 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2765_
timestamp 1646674385
transform -1 0 18216 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1646674385
transform 1 0 19136 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_192
timestamp 1646674385
transform 1 0 18768 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1646674385
transform 1 0 19228 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1646674385
transform 1 0 19044 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1646674385
transform 1 0 18676 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2431__B1
timestamp 1646674385
transform -1 0 18676 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1646674385
transform 1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1646674385
transform 1 0 20240 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1646674385
transform 1 0 19688 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2445__B2
timestamp 1646674385
transform -1 0 20240 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2763_
timestamp 1646674385
transform -1 0 20332 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1646674385
transform 1 0 20884 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1646674385
transform 1 0 20332 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_214
timestamp 1646674385
transform 1 0 20792 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2486__A2
timestamp 1646674385
transform -1 0 20792 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2446__C
timestamp 1646674385
transform -1 0 20884 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1646674385
transform 1 0 21712 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1646674385
transform 1 0 21712 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1646674385
transform 1 0 21620 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1646674385
transform 1 0 21344 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2498__C
timestamp 1646674385
transform -1 0 21988 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2488__B1
timestamp 1646674385
transform -1 0 21344 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2486__B2
timestamp 1646674385
transform -1 0 21988 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_227
timestamp 1646674385
transform 1 0 21988 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1646674385
transform 1 0 21988 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2565__A1
timestamp 1646674385
transform -1 0 22540 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2565__A3
timestamp 1646674385
transform -1 0 23092 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2565__B1
timestamp 1646674385
transform -1 0 23644 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1646674385
transform 1 0 22540 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_239
timestamp 1646674385
transform 1 0 23092 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1646674385
transform 1 0 23644 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_244
timestamp 1646674385
transform 1 0 23552 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1606_
timestamp 1646674385
transform -1 0 23552 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1646674385
transform -1 0 25116 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2469_
timestamp 1646674385
transform 1 0 24380 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1646674385
transform 1 0 24288 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_256
timestamp 1646674385
transform 1 0 24656 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_252
timestamp 1646674385
transform 1 0 24288 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1646674385
transform 1 0 24380 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1646674385
transform 1 0 24196 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1611_
timestamp 1646674385
transform -1 0 26312 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_261
timestamp 1646674385
transform 1 0 25116 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2748_
timestamp 1646674385
transform -1 0 26496 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1646674385
transform 1 0 26864 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1646674385
transform 1 0 26864 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_281
timestamp 1646674385
transform 1 0 26956 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1646674385
transform 1 0 26496 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1646674385
transform 1 0 26312 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__A
timestamp 1646674385
transform -1 0 27140 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1646674385
transform 1 0 27692 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_283
timestamp 1646674385
transform 1 0 27140 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2607__CLK
timestamp 1646674385
transform -1 0 27692 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2747_
timestamp 1646674385
transform -1 0 28520 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_298
timestamp 1646674385
transform 1 0 28520 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_295
timestamp 1646674385
transform 1 0 28244 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2608__CLK
timestamp 1646674385
transform -1 0 28244 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1646674385
transform 1 0 29072 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1646674385
transform 1 0 28796 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_prog_clk_A
timestamp 1646674385
transform -1 0 28796 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_prog_clk_A
timestamp 1646674385
transform 1 0 28888 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1646674385
transform 1 0 29440 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1646674385
transform 1 0 29624 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_311
timestamp 1646674385
transform 1 0 29716 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1646674385
transform 1 0 29348 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1646674385
transform -1 0 29716 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_prog_clk_A
timestamp 1646674385
transform 1 0 29440 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_316
timestamp 1646674385
transform 1 0 30176 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1646674385
transform -1 0 30176 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1646674385
transform -1 0 30268 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output29
timestamp 1646674385
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1646674385
transform -1 0 32016 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1646674385
transform -1 0 32016 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_329
timestamp 1646674385
transform 1 0 31372 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_324
timestamp 1646674385
transform 1 0 30912 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_329
timestamp 1646674385
transform 1 0 31372 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_317
timestamp 1646674385
transform 1 0 30268 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1646674385
transform -1 0 1564 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1646674385
transform -1 0 2116 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1646674385
transform -1 0 2668 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1646674385
transform 1 0 2116 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1646674385
transform 1 0 2668 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_5
timestamp 1646674385
transform 1 0 1564 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1646674385
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1646674385
transform -1 0 3220 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1646674385
transform -1 0 3956 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1646674385
transform 1 0 3220 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1646674385
transform 1 0 3588 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_31
timestamp 1646674385
transform 1 0 3956 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1646674385
transform 1 0 3680 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2837__CLK
timestamp 1646674385
transform -1 0 6992 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_prog_clk_A
timestamp 1646674385
transform 1 0 5980 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_43
timestamp 1646674385
transform 1 0 5060 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1646674385
transform 1 0 5796 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_55
timestamp 1646674385
transform 1 0 6164 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1646674385
transform 1 0 6716 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2838__CLK
timestamp 1646674385
transform -1 0 7544 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_prog_clk_A
timestamp 1646674385
transform 1 0 8280 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1646674385
transform 1 0 6992 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_70
timestamp 1646674385
transform 1 0 7544 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1646674385
transform 1 0 8464 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2495__A
timestamp 1646674385
transform -1 0 10212 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2616__CLK
timestamp 1646674385
transform -1 0 9660 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_prog_clk_A
timestamp 1646674385
transform 1 0 8924 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1646674385
transform 1 0 9108 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1646674385
transform 1 0 9660 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1646674385
transform 1 0 10212 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1646674385
transform 1 0 8832 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2624_
timestamp 1646674385
transform -1 0 12052 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2195__C
timestamp 1646674385
transform 1 0 12604 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_119
timestamp 1646674385
transform 1 0 12052 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2199__A2
timestamp 1646674385
transform -1 0 13340 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_127
timestamp 1646674385
transform 1 0 12788 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1646674385
transform 1 0 13340 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1646674385
transform 1 0 13892 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1646674385
transform 1 0 13984 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2600_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 14076 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_160
timestamp 1646674385
transform 1 0 15824 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_168
timestamp 1646674385
transform 1 0 16560 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1646674385
transform 1 0 16928 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2513_
timestamp 1646674385
transform 1 0 16652 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2764_
timestamp 1646674385
transform -1 0 18768 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1646674385
transform 1 0 18768 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1646674385
transform 1 0 19228 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1646674385
transform 1 0 19136 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2762_
timestamp 1646674385
transform -1 0 21068 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1646674385
transform 1 0 21068 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2751_
timestamp 1646674385
transform 1 0 21436 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2497__B2
timestamp 1646674385
transform -1 0 23460 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_237
timestamp 1646674385
transform 1 0 22908 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_243
timestamp 1646674385
transform 1 0 23460 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1646674385
transform 1 0 24196 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_269
timestamp 1646674385
transform 1 0 25852 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1646674385
transform 1 0 24288 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2749_
timestamp 1646674385
transform -1 0 25852 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_276
timestamp 1646674385
transform 1 0 26496 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2460_
timestamp 1646674385
transform 1 0 26220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2746_
timestamp 1646674385
transform 1 0 27048 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2569__A
timestamp 1646674385
transform 1 0 28888 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_prog_clk_A
timestamp 1646674385
transform 1 0 29532 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_298
timestamp 1646674385
transform 1 0 28520 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1646674385
transform 1 0 29072 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_311
timestamp 1646674385
transform 1 0 29716 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1646674385
transform 1 0 29440 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_prog_clk_A
timestamp 1646674385
transform 1 0 30084 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_A
timestamp 1646674385
transform 1 0 30912 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_317
timestamp 1646674385
transform 1 0 30268 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_323
timestamp 1646674385
transform 1 0 30820 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_326
timestamp 1646674385
transform 1 0 31096 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_332
timestamp 1646674385
transform 1 0 31648 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1646674385
transform -1 0 32016 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1646674385
transform -1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1646674385
transform -1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1646674385
transform 1 0 2484 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1646674385
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1646674385
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_7
timestamp 1646674385
transform 1 0 1748 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1646674385
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2823__CLK
timestamp 1646674385
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1646674385
transform -1 0 3312 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_24
timestamp 1646674385
transform 1 0 3312 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_34
timestamp 1646674385
transform 1 0 4232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2835__CLK
timestamp 1646674385
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2836__CLK
timestamp 1646674385
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_46
timestamp 1646674385
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1646674385
transform 1 0 5796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1646674385
transform 1 0 6164 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_59
timestamp 1646674385
transform 1 0 6532 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1646674385
transform 1 0 6256 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2269__A2
timestamp 1646674385
transform -1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1646674385
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_70
timestamp 1646674385
transform 1 0 7544 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_78
timestamp 1646674385
transform 1 0 8280 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2626_
timestamp 1646674385
transform -1 0 9844 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1646674385
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1820_
timestamp 1646674385
transform -1 0 11040 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1646674385
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_122
timestamp 1646674385
transform 1 0 12328 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1646674385
transform 1 0 11408 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1822_
timestamp 1646674385
transform 1 0 11500 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1818__A
timestamp 1646674385
transform -1 0 12880 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_128
timestamp 1646674385
transform 1 0 12880 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_137
timestamp 1646674385
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_144
timestamp 1646674385
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2219_
timestamp 1646674385
transform 1 0 14076 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2515_
timestamp 1646674385
transform -1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1646674385
transform 1 0 16192 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2766_
timestamp 1646674385
transform 1 0 14720 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1646674385
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1646674385
transform 1 0 16560 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1580_
timestamp 1646674385
transform -1 0 17480 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1583_
timestamp 1646674385
transform 1 0 17848 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1646674385
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_204
timestamp 1646674385
transform 1 0 19872 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1586_
timestamp 1646674385
transform 1 0 19044 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1646674385
transform 1 0 21344 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1646674385
transform 1 0 21712 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 21344 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2752_
timestamp 1646674385
transform 1 0 21804 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_241
timestamp 1646674385
transform 1 0 23276 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_245
timestamp 1646674385
transform 1 0 23644 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2750_
timestamp 1646674385
transform -1 0 25208 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_262
timestamp 1646674385
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1604_
timestamp 1646674385
transform 1 0 25576 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1646674385
transform 1 0 26496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_291
timestamp 1646674385
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1646674385
transform 1 0 26864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1612_
timestamp 1646674385
transform 1 0 26956 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_3_304
timestamp 1646674385
transform 1 0 29072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_311
timestamp 1646674385
transform 1 0 29716 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1614_
timestamp 1646674385
transform 1 0 28244 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2462_
timestamp 1646674385
transform 1 0 29440 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2570__A
timestamp 1646674385
transform -1 0 30452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_prog_clk_A
timestamp 1646674385
transform -1 0 31004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_319
timestamp 1646674385
transform 1 0 30452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp 1646674385
transform 1 0 31004 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1646674385
transform -1 0 32016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2822__CLK
timestamp 1646674385
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_prog_clk_A
timestamp 1646674385
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1646674385
transform -1 0 1656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1646674385
transform 1 0 2208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1646674385
transform 1 0 2760 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1646674385
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_6
timestamp 1646674385
transform 1 0 1656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1646674385
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2817__CLK
timestamp 1646674385
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2819__CLK
timestamp 1646674385
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2820__CLK
timestamp 1646674385
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1646674385
transform 1 0 3312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_31
timestamp 1646674385
transform 1 0 3956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1646674385
transform 1 0 4508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_41
timestamp 1646674385
transform 1 0 4876 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1646674385
transform 1 0 3680 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2206__A2
timestamp 1646674385
transform -1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2270__A2
timestamp 1646674385
transform -1 0 6900 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2830__CLK
timestamp 1646674385
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2834__CLK
timestamp 1646674385
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 1646674385
transform 1 0 5152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_50
timestamp 1646674385
transform 1 0 5704 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1646674385
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1646674385
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2267__A2
timestamp 1646674385
transform -1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2268__A2
timestamp 1646674385
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1646674385
transform 1 0 6900 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_69
timestamp 1646674385
transform 1 0 7452 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1646674385
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1646674385
transform 1 0 8464 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_104
timestamp 1646674385
transform 1 0 10672 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1646674385
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_91
timestamp 1646674385
transform 1 0 9476 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1646674385
transform 1 0 8832 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1821_
timestamp 1646674385
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2216_
timestamp 1646674385
transform -1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_112
timestamp 1646674385
transform 1 0 11408 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1646674385
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2214_
timestamp 1646674385
transform -1 0 11776 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2622_
timestamp 1646674385
transform -1 0 13616 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1646674385
transform 1 0 13616 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1646674385
transform 1 0 14076 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1646674385
transform 1 0 14444 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1646674385
transform 1 0 13984 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_162
timestamp 1646674385
transform 1 0 16008 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2767_
timestamp 1646674385
transform 1 0 14536 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_168
timestamp 1646674385
transform 1 0 16560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1646674385
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1646674385
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1589_
timestamp 1646674385
transform -1 0 18768 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2503_
timestamp 1646674385
transform 1 0 17296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2508_
timestamp 1646674385
transform -1 0 16928 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1646674385
transform 1 0 18768 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_200
timestamp 1646674385
transform 1 0 19504 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1646674385
transform 1 0 19136 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2505_
timestamp 1646674385
transform 1 0 19228 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2761_
timestamp 1646674385
transform -1 0 21528 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_222
timestamp 1646674385
transform 1 0 21528 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1587_
timestamp 1646674385
transform 1 0 21896 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_230
timestamp 1646674385
transform 1 0 22264 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1646674385
transform 1 0 23736 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1600_
timestamp 1646674385
transform -1 0 23736 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_4_262
timestamp 1646674385
transform 1 0 25208 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1646674385
transform 1 0 24288 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1605_
timestamp 1646674385
transform -1 0 25208 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1615_
timestamp 1646674385
transform 1 0 25760 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_277
timestamp 1646674385
transform 1 0 26588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 1646674385
transform 1 0 27876 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1610_
timestamp 1646674385
transform 1 0 26956 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1646674385
transform 1 0 29072 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1646674385
transform 1 0 29440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1613_
timestamp 1646674385
transform -1 0 29072 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2471_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 30176 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2568__A
timestamp 1646674385
transform 1 0 30912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_316
timestamp 1646674385
transform 1 0 30176 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_326
timestamp 1646674385
transform 1 0 31096 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_332
timestamp 1646674385
transform 1 0 31648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1646674385
transform -1 0 32016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2816__CLK
timestamp 1646674385
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_13
timestamp 1646674385
transform 1 0 2300 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1646674385
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1646674385
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input13
timestamp 1646674385
transform 1 0 1748 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2207__A1
timestamp 1646674385
transform -1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2815__CLK
timestamp 1646674385
transform 1 0 3864 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_21
timestamp 1646674385
transform 1 0 3036 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_29
timestamp 1646674385
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1646674385
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1646674385
transform 1 0 4600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2203__A2
timestamp 1646674385
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2204__A2
timestamp 1646674385
transform -1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2205__A1
timestamp 1646674385
transform -1 0 5888 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_44
timestamp 1646674385
transform 1 0 5152 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1646674385
transform 1 0 5888 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_59
timestamp 1646674385
transform 1 0 6532 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1646674385
transform 1 0 6256 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2184__A2
timestamp 1646674385
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_67
timestamp 1646674385
transform 1 0 7268 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_70
timestamp 1646674385
transform 1 0 7544 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2627_
timestamp 1646674385
transform -1 0 9384 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1646674385
transform 1 0 10580 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_90
timestamp 1646674385
transform 1 0 9384 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1819_
timestamp 1646674385
transform -1 0 10580 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1815__A
timestamp 1646674385
transform -1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1646674385
transform 1 0 11316 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1646674385
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1646674385
transform 1 0 11408 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_prog_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 12052 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1646674385
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2621_
timestamp 1646674385
transform 1 0 14260 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_159
timestamp 1646674385
transform 1 0 15732 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1646674385
transform 1 0 16468 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_172
timestamp 1646674385
transform 1 0 16928 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_187
timestamp 1646674385
transform 1 0 18308 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1646674385
transform 1 0 16560 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2237_
timestamp 1646674385
transform 1 0 16652 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2510_
timestamp 1646674385
transform 1 0 17664 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_5_191
timestamp 1646674385
transform 1 0 18676 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1646674385
transform 1 0 19044 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1646674385
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1588_
timestamp 1646674385
transform 1 0 19504 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2507_
timestamp 1646674385
transform -1 0 19044 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2429__A2
timestamp 1646674385
transform -1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_209
timestamp 1646674385
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1646674385
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1646674385
transform 1 0 21620 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1646674385
transform 1 0 21804 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1646674385
transform 1 0 21712 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2470_
timestamp 1646674385
transform -1 0 22448 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_232
timestamp 1646674385
transform 1 0 22448 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_248
timestamp 1646674385
transform 1 0 23920 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1595_
timestamp 1646674385
transform -1 0 23920 0 -1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_5_252
timestamp 1646674385
transform 1 0 24288 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_262
timestamp 1646674385
transform 1 0 25208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1607_
timestamp 1646674385
transform -1 0 25208 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1608_
timestamp 1646674385
transform 1 0 25576 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1646674385
transform 1 0 26404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1646674385
transform 1 0 26772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_281
timestamp 1646674385
transform 1 0 26956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_285
timestamp 1646674385
transform 1 0 27324 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1646674385
transform 1 0 26864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2461_
timestamp 1646674385
transform 1 0 27048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2745_
timestamp 1646674385
transform 1 0 27692 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2557__C
timestamp 1646674385
transform -1 0 29716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1646674385
transform 1 0 29164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_311
timestamp 1646674385
transform 1 0 29716 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2567__A
timestamp 1646674385
transform -1 0 30728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_319
timestamp 1646674385
transform 1 0 30452 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_322
timestamp 1646674385
transform 1 0 30728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_329
timestamp 1646674385
transform 1 0 31372 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1646674385
transform -1 0 32016 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output41
timestamp 1646674385
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1646674385
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1646674385
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1646674385
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1646674385
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1646674385
transform 1 0 1840 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1646674385
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2818__CLK
timestamp 1646674385
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1646674385
transform 1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1646674385
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1646674385
transform 1 0 2392 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2173__A2
timestamp 1646674385
transform -1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2088__A2
timestamp 1646674385
transform 1 0 2484 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1646674385
transform 1 0 2944 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2171__A2
timestamp 1646674385
transform -1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1646674385
transform 1 0 3680 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_29
timestamp 1646674385
transform 1 0 3772 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1646674385
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_31
timestamp 1646674385
transform 1 0 3956 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2169__A2
timestamp 1646674385
transform -1 0 3956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2168__B
timestamp 1646674385
transform -1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2089__A1
timestamp 1646674385
transform -1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1458_
timestamp 1646674385
transform -1 0 5244 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp 1646674385
transform 1 0 4324 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1646674385
transform 1 0 4324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2831_
timestamp 1646674385
transform -1 0 5888 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2202__B
timestamp 1646674385
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2203__A1
timestamp 1646674385
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_52
timestamp 1646674385
transform 1 0 5888 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1646674385
transform 1 0 6624 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_45
timestamp 1646674385
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_49
timestamp 1646674385
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1646674385
transform 1 0 5888 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1646674385
transform 1 0 6256 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1457_
timestamp 1646674385
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__A1
timestamp 1646674385
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1646674385
transform 1 0 7176 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_73
timestamp 1646674385
transform 1 0 7820 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1646674385
transform 1 0 8464 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1646674385
transform 1 0 7176 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1646674385
transform 1 0 7544 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2225_
timestamp 1646674385
transform -1 0 8464 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2226_
timestamp 1646674385
transform -1 0 7820 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2628_
timestamp 1646674385
transform 1 0 7636 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__o221a_1  _1817_
timestamp 1646674385
transform -1 0 9936 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1646674385
transform 1 0 8832 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1646674385
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_87
timestamp 1646674385
transform 1 0 9108 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1646674385
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _2218_
timestamp 1646674385
transform -1 0 10580 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1646674385
transform 1 0 10672 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1646674385
transform 1 0 9936 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1646674385
transform 1 0 10580 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1815_
timestamp 1646674385
transform -1 0 10672 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1646674385
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_122
timestamp 1646674385
transform 1 0 12328 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1646674385
transform 1 0 11408 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1818_
timestamp 1646674385
transform 1 0 10948 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1825_
timestamp 1646674385
transform 1 0 12236 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1829_
timestamp 1646674385
transform 1 0 11500 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1816__A
timestamp 1646674385
transform -1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1646674385
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1646674385
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1646674385
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_143
timestamp 1646674385
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1646674385
transform 1 0 13984 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1827_
timestamp 1646674385
transform -1 0 13524 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2221_
timestamp 1646674385
transform -1 0 14720 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2768_
timestamp 1646674385
transform -1 0 15824 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_6_148
timestamp 1646674385
transform 1 0 14720 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1646674385
transform 1 0 16284 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1646674385
transform 1 0 15824 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1577_
timestamp 1646674385
transform -1 0 16284 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_176
timestamp 1646674385
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1646674385
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1646674385
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1646674385
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1575_
timestamp 1646674385
transform -1 0 18308 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1576_
timestamp 1646674385
transform -1 0 17572 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _2511_
timestamp 1646674385
transform 1 0 17664 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2516_
timestamp 1646674385
transform 1 0 16652 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1646674385
transform 1 0 18492 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1646674385
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1646674385
transform 1 0 20148 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1646674385
transform 1 0 19504 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1646674385
transform 1 0 19136 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1585_
timestamp 1646674385
transform 1 0 19228 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1591_
timestamp 1646674385
transform 1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2760_
timestamp 1646674385
transform 1 0 19872 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_214
timestamp 1646674385
transform 1 0 20792 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1646674385
transform 1 0 21344 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1646674385
transform 1 0 21712 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1594_
timestamp 1646674385
transform -1 0 22632 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2526_
timestamp 1646674385
transform 1 0 20516 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_prog_clk
timestamp 1646674385
transform 1 0 21160 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_6_238
timestamp 1646674385
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_244
timestamp 1646674385
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1646674385
transform 1 0 23920 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_234
timestamp 1646674385
transform 1 0 22632 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2467_
timestamp 1646674385
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2753_
timestamp 1646674385
transform -1 0 24472 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1646674385
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1646674385
transform 1 0 25484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_254
timestamp 1646674385
transform 1 0 24472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_268
timestamp 1646674385
transform 1 0 25760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1646674385
transform 1 0 24288 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1602_
timestamp 1646674385
transform 1 0 24840 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1609_
timestamp 1646674385
transform 1 0 24564 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_prog_clk
timestamp 1646674385
transform 1 0 25852 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1646674385
transform 1 0 27692 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1646674385
transform 1 0 26404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1646674385
transform 1 0 26772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_284
timestamp 1646674385
transform 1 0 27232 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1646674385
transform 1 0 26864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2451_
timestamp 1646674385
transform -1 0 27232 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2463_
timestamp 1646674385
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2744_
timestamp 1646674385
transform -1 0 29072 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2550__A3
timestamp 1646674385
transform 1 0 29808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2553__C
timestamp 1646674385
transform -1 0 29716 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_300
timestamp 1646674385
transform 1 0 28704 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_311
timestamp 1646674385
transform 1 0 29716 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_304
timestamp 1646674385
transform 1 0 29072 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1646674385
transform 1 0 29440 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _2464_
timestamp 1646674385
transform 1 0 28060 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_7_314
timestamp 1646674385
transform 1 0 29992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_317
timestamp 1646674385
transform 1 0 30268 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2556__C
timestamp 1646674385
transform -1 0 30268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2542__C
timestamp 1646674385
transform 1 0 30360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_326
timestamp 1646674385
transform 1 0 31096 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1646674385
transform 1 0 30544 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_326
timestamp 1646674385
transform 1 0 31096 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_323
timestamp 1646674385
transform 1 0 30820 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2566__A
timestamp 1646674385
transform 1 0 30912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2549__C
timestamp 1646674385
transform -1 0 31096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1646674385
transform -1 0 32016 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1646674385
transform -1 0 32016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_332
timestamp 1646674385
transform 1 0 31648 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_332
timestamp 1646674385
transform 1 0 31648 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1646674385
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1646674385
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2817_
timestamp 1646674385
transform 1 0 1656 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1646674385
transform 1 0 3128 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1646674385
transform 1 0 3680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2830_
timestamp 1646674385
transform 1 0 3772 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_45
timestamp 1646674385
transform 1 0 5244 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_53
timestamp 1646674385
transform 1 0 5980 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2832_
timestamp 1646674385
transform -1 0 7544 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1646674385
transform 1 0 7544 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1646674385
transform 1 0 8280 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1456_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_103
timestamp 1646674385
transform 1 0 10580 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1646674385
transform 1 0 8924 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_89
timestamp 1646674385
transform 1 0 9292 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1646674385
transform 1 0 8832 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1810_
timestamp 1646674385
transform -1 0 10580 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2224_
timestamp 1646674385
transform -1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_117
timestamp 1646674385
transform 1 0 11868 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1816_
timestamp 1646674385
transform 1 0 10948 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1828_
timestamp 1646674385
transform 1 0 12604 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1646674385
transform 1 0 13432 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1646674385
transform 1 0 14076 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1646674385
transform 1 0 13984 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2769_
timestamp 1646674385
transform 1 0 14352 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_160
timestamp 1646674385
transform 1 0 15824 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_166
timestamp 1646674385
transform 1 0 16376 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_176
timestamp 1646674385
transform 1 0 17296 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_182
timestamp 1646674385
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2517_
timestamp 1646674385
transform 1 0 16468 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2528_
timestamp 1646674385
transform 1 0 17940 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1646674385
transform 1 0 18768 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 1646674385
transform 1 0 19228 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_208
timestamp 1646674385
transform 1 0 20240 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1646674385
transform 1 0 19136 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1584_
timestamp 1646674385
transform 1 0 19320 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_8_212
timestamp 1646674385
transform 1 0 20608 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1646674385
transform 1 0 22172 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2758_
timestamp 1646674385
transform -1 0 22172 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1646674385
transform 1 0 23460 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1592_
timestamp 1646674385
transform 1 0 22540 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1646674385
transform 1 0 24196 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_262
timestamp 1646674385
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1646674385
transform 1 0 24288 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1603_
timestamp 1646674385
transform -1 0 25208 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2465_
timestamp 1646674385
transform -1 0 26404 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_275
timestamp 1646674385
transform 1 0 26404 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_290
timestamp 1646674385
transform 1 0 27784 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1616_
timestamp 1646674385
transform 1 0 26956 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1602__A
timestamp 1646674385
transform 1 0 28152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2499__B1
timestamp 1646674385
transform -1 0 28888 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2536__A
timestamp 1646674385
transform -1 0 29716 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_296
timestamp 1646674385
transform 1 0 28336 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1646674385
transform 1 0 28888 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_311
timestamp 1646674385
transform 1 0 29716 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1646674385
transform 1 0 29440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2541__C
timestamp 1646674385
transform 1 0 30544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_319
timestamp 1646674385
transform 1 0 30452 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_322
timestamp 1646674385
transform 1 0 30728 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_329
timestamp 1646674385
transform 1 0 31372 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1646674385
transform -1 0 32016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output32
timestamp 1646674385
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1646674385
transform 1 0 2392 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1646674385
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1646674385
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1646674385
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1908_
timestamp 1646674385
transform -1 0 2392 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1910_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 1748 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2084_
timestamp 1646674385
transform -1 0 3036 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__B2
timestamp 1646674385
transform -1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1646674385
transform 1 0 3036 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1646674385
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1646674385
transform 1 0 4784 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1460_
timestamp 1646674385
transform -1 0 4784 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1646674385
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1646674385
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_2  _2203_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 6348 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _2206_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 5152 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_67
timestamp 1646674385
transform 1 0 7268 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_71
timestamp 1646674385
transform 1 0 7636 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2629_
timestamp 1646674385
transform 1 0 7728 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1646674385
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1646674385
transform 1 0 9844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2222_
timestamp 1646674385
transform 1 0 10212 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2223_
timestamp 1646674385
transform 1 0 9568 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1646674385
transform 1 0 11040 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1646674385
transform 1 0 11500 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_124
timestamp 1646674385
transform 1 0 12512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1646674385
transform 1 0 11408 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1823_
timestamp 1646674385
transform 1 0 11592 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_9_144
timestamp 1646674385
transform 1 0 14352 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2620_
timestamp 1646674385
transform -1 0 14352 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_150
timestamp 1646674385
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1646674385
transform 1 0 15824 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1573_
timestamp 1646674385
transform -1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1646674385
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_175
timestamp 1646674385
transform 1 0 17204 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_186
timestamp 1646674385
transform 1 0 18216 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1646674385
transform 1 0 16560 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2509_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 17204 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2527_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 18216 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_9_194
timestamp 1646674385
transform 1 0 18952 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2759_
timestamp 1646674385
transform -1 0 20516 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__A
timestamp 1646674385
transform -1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1646674385
transform 1 0 20516 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1646674385
transform 1 0 21160 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1646674385
transform 1 0 21804 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1646674385
transform 1 0 21712 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2525_
timestamp 1646674385
transform -1 0 21160 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1646674385
transform 1 0 22264 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_250
timestamp 1646674385
transform 1 0 24104 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2754_
timestamp 1646674385
transform -1 0 24104 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_263
timestamp 1646674385
transform 1 0 25300 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2459_
timestamp 1646674385
transform -1 0 26496 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2472_
timestamp 1646674385
transform -1 0 25300 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1646674385
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_284
timestamp 1646674385
transform 1 0 27232 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_291
timestamp 1646674385
transform 1 0 27876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1646674385
transform 1 0 26864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2453_
timestamp 1646674385
transform -1 0 27232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2455_
timestamp 1646674385
transform 1 0 27600 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2454__B
timestamp 1646674385
transform -1 0 29072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2518__A
timestamp 1646674385
transform 1 0 29440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_298
timestamp 1646674385
transform 1 0 28520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_304
timestamp 1646674385
transform 1 0 29072 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_310
timestamp 1646674385
transform 1 0 29624 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2456_
timestamp 1646674385
transform -1 0 28520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2529__A1
timestamp 1646674385
transform -1 0 30176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2534__A3
timestamp 1646674385
transform 1 0 30544 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2538__C
timestamp 1646674385
transform -1 0 31280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_316
timestamp 1646674385
transform 1 0 30176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_322
timestamp 1646674385
transform 1 0 30728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_328
timestamp 1646674385
transform 1 0 31280 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_332
timestamp 1646674385
transform 1 0 31648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1646674385
transform -1 0 32016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_11
timestamp 1646674385
transform 1 0 2116 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp 1646674385
transform 1 0 2668 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1646674385
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1646674385
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1486_
timestamp 1646674385
transform 1 0 2760 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1646674385
transform 1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1646674385
transform 1 0 3312 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1646674385
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_33
timestamp 1646674385
transform 1 0 4140 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_40
timestamp 1646674385
transform 1 0 4784 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1646674385
transform 1 0 3680 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1903_
timestamp 1646674385
transform -1 0 4784 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1904_
timestamp 1646674385
transform -1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1646674385
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _2208_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 7912 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2576_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 5980 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1824__A
timestamp 1646674385
transform -1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_74
timestamp 1646674385
transform 1 0 7912 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1646674385
transform 1 0 8464 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1646674385
transform 1 0 9752 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1646674385
transform 1 0 8832 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1813_
timestamp 1646674385
transform 1 0 8924 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1814_
timestamp 1646674385
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1810__A
timestamp 1646674385
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1646674385
transform 1 0 10948 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_113
timestamp 1646674385
transform 1 0 11500 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1824_
timestamp 1646674385
transform -1 0 12788 0 1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1646674385
transform 1 0 12788 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1646674385
transform 1 0 13432 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1646674385
transform 1 0 13984 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1830_
timestamp 1646674385
transform -1 0 14904 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2236_
timestamp 1646674385
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1823__A
timestamp 1646674385
transform -1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1646674385
transform 1 0 14904 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_156
timestamp 1646674385
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1646674385
transform 1 0 16100 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2500_
timestamp 1646674385
transform -1 0 16100 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1646674385
transform 1 0 16744 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_179
timestamp 1646674385
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1646674385
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2484_
timestamp 1646674385
transform 1 0 17940 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2489_
timestamp 1646674385
transform -1 0 16744 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2490_
timestamp 1646674385
transform 1 0 17112 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2194__A2
timestamp 1646674385
transform -1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1646674385
transform 1 0 18768 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1646674385
transform 1 0 19228 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1646674385
transform 1 0 19136 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1590_
timestamp 1646674385
transform 1 0 19504 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2199__B2
timestamp 1646674385
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1646674385
transform 1 0 20332 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1646674385
transform 1 0 20884 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_229
timestamp 1646674385
transform 1 0 22172 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1578_
timestamp 1646674385
transform -1 0 22172 0 1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__A
timestamp 1646674385
transform 1 0 23736 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_242
timestamp 1646674385
transform 1 0 23368 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1646674385
transform 1 0 23920 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1599_
timestamp 1646674385
transform 1 0 22540 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_263
timestamp 1646674385
transform 1 0 25300 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1646674385
transform 1 0 24288 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1574_
timestamp 1646674385
transform 1 0 24380 0 1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1619__A
timestamp 1646674385
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_278
timestamp 1646674385
transform 1 0 26680 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_284
timestamp 1646674385
transform 1 0 27232 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2458_
timestamp 1646674385
transform 1 0 26036 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2743_
timestamp 1646674385
transform 1 0 27600 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2457__B
timestamp 1646674385
transform 1 0 29532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1646674385
transform 1 0 29072 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_311
timestamp 1646674385
transform 1 0 29716 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1646674385
transform 1 0 29440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2487__C
timestamp 1646674385
transform -1 0 30268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2533__C
timestamp 1646674385
transform 1 0 30820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_317
timestamp 1646674385
transform 1 0 30268 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_325
timestamp 1646674385
transform 1 0 31004 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1646674385
transform -1 0 32016 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1646674385
transform 1 0 2392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1646674385
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1646674385
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2089_
timestamp 1646674385
transform -1 0 2392 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2577_
timestamp 1646674385
transform -1 0 3588 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_27
timestamp 1646674385
transform 1 0 3588 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_35
timestamp 1646674385
transform 1 0 4324 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1646674385
transform 1 0 4784 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2207_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 4416 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2090__A2
timestamp 1646674385
transform -1 0 6532 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1646674385
transform 1 0 5888 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_59
timestamp 1646674385
transform 1 0 6532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1646674385
transform 1 0 6256 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2204_
timestamp 1646674385
transform 1 0 5152 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_prog_clk
timestamp 1646674385
transform 1 0 7268 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_11_87
timestamp 1646674385
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2630_
timestamp 1646674385
transform -1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1646674385
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1646674385
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1646674385
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1646674385
transform 1 0 12512 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1646674385
transform 1 0 11408 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2239_
timestamp 1646674385
transform 1 0 11684 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_144
timestamp 1646674385
transform 1 0 14352 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2619_
timestamp 1646674385
transform -1 0 14352 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_150
timestamp 1646674385
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1646674385
transform 1 0 15824 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1572_
timestamp 1646674385
transform -1 0 15824 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1646674385
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_176
timestamp 1646674385
transform 1 0 17296 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1646674385
transform 1 0 16560 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2501_
timestamp 1646674385
transform 1 0 18032 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2504_
timestamp 1646674385
transform 1 0 16836 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_11_189
timestamp 1646674385
transform 1 0 18492 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_201
timestamp 1646674385
transform 1 0 19596 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_208
timestamp 1646674385
transform 1 0 20240 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2502_
timestamp 1646674385
transform 1 0 19964 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2531_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 19228 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1646674385
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1646674385
transform 1 0 21620 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1646674385
transform 1 0 21804 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1646674385
transform 1 0 21712 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1598_
timestamp 1646674385
transform -1 0 22816 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2512_
timestamp 1646674385
transform 1 0 20608 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_236
timestamp 1646674385
transform 1 0 22816 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_244
timestamp 1646674385
transform 1 0 23552 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1646674385
transform 1 0 23920 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2468_
timestamp 1646674385
transform 1 0 23644 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1646674385
transform 1 0 24748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_269
timestamp 1646674385
transform 1 0 25852 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2466_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 24748 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _2478_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 25852 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1646674385
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1646674385
transform 1 0 26956 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1646674385
transform 1 0 26864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1620_
timestamp 1646674385
transform 1 0 27140 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2443_
timestamp 1646674385
transform 1 0 26220 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2395__B1
timestamp 1646674385
transform 1 0 28336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2436__B1
timestamp 1646674385
transform 1 0 28888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2441__C
timestamp 1646674385
transform -1 0 29624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_292
timestamp 1646674385
transform 1 0 27968 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_298
timestamp 1646674385
transform 1 0 28520 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_304
timestamp 1646674385
transform 1 0 29072 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_310
timestamp 1646674385
transform 1 0 29624 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2447__B1
timestamp 1646674385
transform 1 0 29992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2475__B
timestamp 1646674385
transform -1 0 30728 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_316
timestamp 1646674385
transform 1 0 30176 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_322
timestamp 1646674385
transform 1 0 30728 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_329
timestamp 1646674385
transform 1 0 31372 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1646674385
transform -1 0 32016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2568_
timestamp 1646674385
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_10
timestamp 1646674385
transform 1 0 2024 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1646674385
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1646674385
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _2086_
timestamp 1646674385
transform 1 0 2392 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _2088_
timestamp 1646674385
transform -1 0 2024 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1646674385
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1646674385
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1646674385
transform 1 0 4876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1646674385
transform 1 0 3680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2083_
timestamp 1646674385
transform 1 0 4600 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2085_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 4232 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2086__A1
timestamp 1646674385
transform -1 0 6256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_45
timestamp 1646674385
transform 1 0 5244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_50
timestamp 1646674385
transform 1 0 5704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_56
timestamp 1646674385
transform 1 0 6256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2202_
timestamp 1646674385
transform 1 0 6624 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2205_
timestamp 1646674385
transform -1 0 5704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_65
timestamp 1646674385
transform 1 0 7084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp 1646674385
transform 1 0 7820 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1646674385
transform 1 0 8188 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1646674385
transform 1 0 8740 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1905_
timestamp 1646674385
transform 1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1646674385
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_94
timestamp 1646674385
transform 1 0 9752 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1646674385
transform 1 0 8832 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1812_
timestamp 1646674385
transform -1 0 9752 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2228_
timestamp 1646674385
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_112
timestamp 1646674385
transform 1 0 11408 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1646674385
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _2238_
timestamp 1646674385
transform -1 0 12420 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1646674385
transform 1 0 13248 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1646674385
transform 1 0 13984 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2220_
timestamp 1646674385
transform 1 0 12788 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2229_
timestamp 1646674385
transform 1 0 14076 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_12_146
timestamp 1646674385
transform 1 0 14536 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1646674385
transform 1 0 15732 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_163
timestamp 1646674385
transform 1 0 16100 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1571_
timestamp 1646674385
transform -1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2523_
timestamp 1646674385
transform -1 0 16836 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__A
timestamp 1646674385
transform -1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_171
timestamp 1646674385
transform 1 0 16836 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1646674385
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2529_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 17756 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1646674385
transform 1 0 18492 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1646674385
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1646674385
transform 1 0 19688 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1646674385
transform 1 0 19136 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1593_
timestamp 1646674385
transform 1 0 20056 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1845_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 19228 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_12_216
timestamp 1646674385
transform 1 0 20976 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2755_
timestamp 1646674385
transform 1 0 21344 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2209__C
timestamp 1646674385
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2377__A2
timestamp 1646674385
transform 1 0 23736 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1646674385
transform 1 0 22816 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_242
timestamp 1646674385
transform 1 0 23368 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1646674385
transform 1 0 23920 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_253
timestamp 1646674385
transform 1 0 24380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1646674385
transform 1 0 24840 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_270
timestamp 1646674385
transform 1 0 25944 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1646674385
transform 1 0 24288 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _2477_
timestamp 1646674385
transform 1 0 25208 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _2479_
timestamp 1646674385
transform -1 0 24840 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_284
timestamp 1646674385
transform 1 0 27232 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1619_
timestamp 1646674385
transform 1 0 26312 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2742_
timestamp 1646674385
transform -1 0 29072 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2437__A
timestamp 1646674385
transform 1 0 29532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1646674385
transform 1 0 29072 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_311
timestamp 1646674385
transform 1 0 29716 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1646674385
transform 1 0 29440 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2440__A2
timestamp 1646674385
transform -1 0 30268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_317
timestamp 1646674385
transform 1 0 30268 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_325
timestamp 1646674385
transform 1 0 31004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_329
timestamp 1646674385
transform 1 0 31372 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1646674385
transform -1 0 32016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1646674385
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2087_
timestamp 1646674385
transform 1 0 1748 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1909_
timestamp 1646674385
transform -1 0 1840 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1646674385
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1646674385
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1646674385
transform 1 0 1840 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1646674385
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1646674385
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2090_
timestamp 1646674385
transform 1 0 2208 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1907_
timestamp 1646674385
transform -1 0 3220 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1646674385
transform 1 0 2576 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1646674385
transform 1 0 2852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1646674385
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _2091_
timestamp 1646674385
transform -1 0 4508 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2085__B
timestamp 1646674385
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1646674385
transform 1 0 4508 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1646674385
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1646674385
transform 1 0 3588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1646674385
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1646674385
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2834_
timestamp 1646674385
transform 1 0 3956 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1906_
timestamp 1646674385
transform -1 0 5704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1646674385
transform 1 0 5428 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1646674385
transform 1 0 5704 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1646674385
transform 1 0 5060 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2087__A1
timestamp 1646674385
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _2201_
timestamp 1646674385
transform -1 0 6992 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1646674385
transform 1 0 6256 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_57
timestamp 1646674385
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_53
timestamp 1646674385
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1646674385
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2833_
timestamp 1646674385
transform -1 0 7912 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_64
timestamp 1646674385
transform 1 0 6992 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2200_
timestamp 1646674385
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1646674385
transform 1 0 7728 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_68
timestamp 1646674385
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2232_
timestamp 1646674385
transform -1 0 8464 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_74
timestamp 1646674385
transform 1 0 7912 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_76
timestamp 1646674385
transform 1 0 8096 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1646674385
transform 1 0 8464 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_80
timestamp 1646674385
transform 1 0 8464 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1831__C1
timestamp 1646674385
transform -1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_93
timestamp 1646674385
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_97
timestamp 1646674385
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_104
timestamp 1646674385
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1646674385
transform 1 0 8924 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1646674385
transform 1 0 8832 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1811_
timestamp 1646674385
transform 1 0 8832 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2227_
timestamp 1646674385
transform -1 0 10764 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2632_
timestamp 1646674385
transform 1 0 9200 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1646674385
transform 1 0 10764 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1646674385
transform 1 0 11316 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_120
timestamp 1646674385
transform 1 0 12144 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1646674385
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1646674385
transform 1 0 11408 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2189_
timestamp 1646674385
transform -1 0 12972 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2234_
timestamp 1646674385
transform 1 0 11500 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2235_
timestamp 1646674385
transform 1 0 11040 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _2241_
timestamp 1646674385
transform -1 0 12972 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2212_
timestamp 1646674385
transform -1 0 13800 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2188_
timestamp 1646674385
transform 1 0 13340 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1646674385
transform 1 0 12972 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1646674385
transform 1 0 12972 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1646674385
transform 1 0 13984 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1646674385
transform 1 0 13616 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_142
timestamp 1646674385
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1646674385
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2771_
timestamp 1646674385
transform -1 0 15548 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2770_
timestamp 1646674385
transform -1 0 15732 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1646674385
transform 1 0 15732 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_157
timestamp 1646674385
transform 1 0 15548 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2495_
timestamp 1646674385
transform 1 0 16284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2524_
timestamp 1646674385
transform 1 0 16652 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2506_
timestamp 1646674385
transform -1 0 17388 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1646674385
transform 1 0 16560 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1646674385
transform 1 0 16560 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1646674385
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2592_
timestamp 1646674385
transform -1 0 18768 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _2530_
timestamp 1646674385
transform -1 0 18492 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1646674385
transform 1 0 17388 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1646674385
transform 1 0 17848 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1646674385
transform 1 0 17480 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_192
timestamp 1646674385
transform 1 0 18768 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1646674385
transform 1 0 18492 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1646674385
transform 1 0 19044 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1646674385
transform 1 0 19228 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1646674385
transform 1 0 19596 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1646674385
transform 1 0 19136 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1837_
timestamp 1646674385
transform -1 0 19596 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2610_
timestamp 1646674385
transform 1 0 19136 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2615_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 19964 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2194__B2
timestamp 1646674385
transform 1 0 20976 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_212
timestamp 1646674385
transform 1 0 20608 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1646674385
transform 1 0 21160 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1646674385
transform 1 0 21804 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_222
timestamp 1646674385
transform 1 0 21528 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1646674385
transform 1 0 21712 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1597_
timestamp 1646674385
transform 1 0 21988 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_236
timestamp 1646674385
transform 1 0 22816 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_230
timestamp 1646674385
transform 1 0 22264 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1646674385
transform 1 0 23920 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2756_
timestamp 1646674385
transform 1 0 22356 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2757_
timestamp 1646674385
transform 1 0 23184 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_13_257
timestamp 1646674385
transform 1 0 24748 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_263
timestamp 1646674385
transform 1 0 25300 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_269
timestamp 1646674385
transform 1 0 25852 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1646674385
transform 1 0 24380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_266
timestamp 1646674385
transform 1 0 25576 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1646674385
transform 1 0 24288 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2449_
timestamp 1646674385
transform 1 0 25392 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2450_
timestamp 1646674385
transform 1 0 25944 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2591_
timestamp 1646674385
transform 1 0 24748 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2448_
timestamp 1646674385
transform 1 0 26220 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1626_
timestamp 1646674385
transform 1 0 26588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1646674385
transform 1 0 26864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_273
timestamp 1646674385
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1646674385
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2473_
timestamp 1646674385
transform 1 0 27784 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1623_
timestamp 1646674385
transform 1 0 27048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1646674385
transform 1 0 27416 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 1646674385
transform 1 0 26956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_291
timestamp 1646674385
transform 1 0 27876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2382__A2
timestamp 1646674385
transform -1 0 28612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2390__B1
timestamp 1646674385
transform -1 0 29716 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_311
timestamp 1646674385
transform 1 0 29716 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_293
timestamp 1646674385
transform 1 0 28060 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_299
timestamp 1646674385
transform 1 0 28612 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1646674385
transform 1 0 29348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_311
timestamp 1646674385
transform 1 0 29716 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1646674385
transform 1 0 29440 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2741_
timestamp 1646674385
transform -1 0 29716 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_317
timestamp 1646674385
transform 1 0 30268 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_317
timestamp 1646674385
transform 1 0 30268 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2434__A2
timestamp 1646674385
transform -1 0 30268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2393__B2
timestamp 1646674385
transform 1 0 30084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2440__B2
timestamp 1646674385
transform -1 0 30820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2429__B2
timestamp 1646674385
transform -1 0 30820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_323
timestamp 1646674385
transform 1 0 30820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_323
timestamp 1646674385
transform 1 0 30820 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2445__A2
timestamp 1646674385
transform -1 0 31372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2434__B2
timestamp 1646674385
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_329
timestamp 1646674385
transform 1 0 31372 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_329
timestamp 1646674385
transform 1 0 31372 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1646674385
transform -1 0 32016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1646674385
transform -1 0 32016 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2086__A2
timestamp 1646674385
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_11
timestamp 1646674385
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1646674385
transform 1 0 2668 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1646674385
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1646674385
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1646674385
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1957__A2
timestamp 1646674385
transform -1 0 3864 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1960__A2
timestamp 1646674385
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1646674385
transform 1 0 3036 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1646674385
transform 1 0 3312 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1646674385
transform 1 0 3864 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1454_
timestamp 1646674385
transform -1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_43
timestamp 1646674385
transform 1 0 5060 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1646674385
transform 1 0 5704 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1646674385
transform 1 0 6256 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1455_
timestamp 1646674385
transform 1 0 6348 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1915_
timestamp 1646674385
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1646674385
transform 1 0 7176 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 1646674385
transform 1 0 7544 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2631_
timestamp 1646674385
transform 1 0 7636 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1646674385
transform 1 0 10396 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1646674385
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1646674385
transform 1 0 9752 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2230_
timestamp 1646674385
transform 1 0 10120 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2233_
timestamp 1646674385
transform 1 0 9476 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1646674385
transform 1 0 11040 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1646674385
transform 1 0 11960 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1646674385
transform 1 0 11408 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2165_
timestamp 1646674385
transform -1 0 11040 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2215_
timestamp 1646674385
transform -1 0 11960 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _2240_
timestamp 1646674385
transform -1 0 13064 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_130
timestamp 1646674385
transform 1 0 13064 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_134
timestamp 1646674385
transform 1 0 13432 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1646674385
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2197_
timestamp 1646674385
transform -1 0 13800 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_prog_clk
timestamp 1646674385
transform 1 0 14168 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1646674385
transform 1 0 16008 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1646674385
transform 1 0 16928 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_185
timestamp 1646674385
transform 1 0 18124 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1646674385
transform 1 0 16560 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2211_
timestamp 1646674385
transform 1 0 16652 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2518_
timestamp 1646674385
transform 1 0 17664 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_prog_clk
timestamp 1646674385
transform 1 0 18860 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1836__A
timestamp 1646674385
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_213
timestamp 1646674385
transform 1 0 20700 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_217
timestamp 1646674385
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1646674385
transform 1 0 21344 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1646674385
transform 1 0 21712 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _1836_
timestamp 1646674385
transform -1 0 22264 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1646674385
transform 1 0 22264 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1646674385
transform 1 0 23460 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1596_
timestamp 1646674385
transform 1 0 22632 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1852_
timestamp 1646674385
transform 1 0 23828 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1852__B
timestamp 1646674385
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1646674385
transform 1 0 24288 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_258
timestamp 1646674385
transform 1 0 24840 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_266
timestamp 1646674385
transform 1 0 25576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2476_
timestamp 1646674385
transform -1 0 26496 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1646674385
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1646674385
transform 1 0 26956 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1646674385
transform 1 0 26864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1624_
timestamp 1646674385
transform 1 0 27324 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2382__B2
timestamp 1646674385
transform 1 0 29164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2384__B1
timestamp 1646674385
transform -1 0 29900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_294
timestamp 1646674385
transform 1 0 28152 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_301
timestamp 1646674385
transform 1 0 28796 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_307
timestamp 1646674385
transform 1 0 29348 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2474_
timestamp 1646674385
transform 1 0 28520 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2393__A2
timestamp 1646674385
transform 1 0 30268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2394__C
timestamp 1646674385
transform -1 0 31004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_313
timestamp 1646674385
transform 1 0 29900 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1646674385
transform 1 0 30452 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_325
timestamp 1646674385
transform 1 0 31004 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1646674385
transform -1 0 32016 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1646674385
transform 1 0 2852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1646674385
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2816_
timestamp 1646674385
transform -1 0 2852 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1646674385
transform 1 0 3588 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1646674385
transform 1 0 3772 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1646674385
transform 1 0 4140 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1646674385
transform 1 0 3680 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1960_
timestamp 1646674385
transform -1 0 4968 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1956__B
timestamp 1646674385
transform -1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_42
timestamp 1646674385
transform 1 0 4968 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_48
timestamp 1646674385
transform 1 0 5520 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1646674385
transform 1 0 6256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1449_
timestamp 1646674385
transform -1 0 6256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1453_
timestamp 1646674385
transform -1 0 6992 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__A
timestamp 1646674385
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1807__A
timestamp 1646674385
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1646674385
transform 1 0 6992 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_70
timestamp 1646674385
transform 1 0 7544 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1646674385
transform 1 0 8464 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1806__C1
timestamp 1646674385
transform -1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_100
timestamp 1646674385
transform 1 0 10304 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_103
timestamp 1646674385
transform 1 0 10580 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1646674385
transform 1 0 8924 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1646674385
transform 1 0 9936 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1646674385
transform 1 0 8832 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1807_
timestamp 1646674385
transform 1 0 9016 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_16_109
timestamp 1646674385
transform 1 0 11132 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_115
timestamp 1646674385
transform 1 0 11684 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2217_
timestamp 1646674385
transform -1 0 11684 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2595_
timestamp 1646674385
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1646674385
transform 1 0 13248 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_145
timestamp 1646674385
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1646674385
transform 1 0 13984 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _2242_
timestamp 1646674385
transform 1 0 14076 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1646674385
transform 1 0 15640 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1568_
timestamp 1646674385
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1570_
timestamp 1646674385
transform -1 0 15640 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1646674385
transform 1 0 16836 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1646674385
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1646674385
transform 1 0 18308 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1558_
timestamp 1646674385
transform 1 0 17204 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1559_
timestamp 1646674385
transform -1 0 18308 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1646674385
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1646674385
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1646674385
transform 1 0 19688 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1646674385
transform 1 0 19136 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1846_
timestamp 1646674385
transform 1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2519_
timestamp 1646674385
transform 1 0 20056 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1646674385
transform 1 0 20332 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1646674385
transform 1 0 20700 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2911_
timestamp 1646674385
transform 1 0 20792 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__A1
timestamp 1646674385
transform 1 0 23460 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1646674385
transform 1 0 22264 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_237
timestamp 1646674385
transform 1 0 22908 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1646674385
transform 1 0 23644 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2563_
timestamp 1646674385
transform -1 0 22908 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1646674385
transform 1 0 24196 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 1646674385
transform 1 0 24380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_259
timestamp 1646674385
transform 1 0 24932 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_268
timestamp 1646674385
transform 1 0 25760 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1646674385
transform 1 0 24288 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2432_
timestamp 1646674385
transform 1 0 24656 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2438_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 25300 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1646674385
transform 1 0 26312 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_284
timestamp 1646674385
transform 1 0 27232 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1625_
timestamp 1646674385
transform 1 0 26404 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2740_
timestamp 1646674385
transform -1 0 29072 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2379__B1
timestamp 1646674385
transform 1 0 29532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1646674385
transform 1 0 29072 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_311
timestamp 1646674385
transform 1 0 29716 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1646674385
transform 1 0 29440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2383__C
timestamp 1646674385
transform -1 0 30268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_317
timestamp 1646674385
transform 1 0 30268 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_325
timestamp 1646674385
transform 1 0 31004 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_329
timestamp 1646674385
transform 1 0 31372 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1646674385
transform -1 0 32016 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output33
timestamp 1646674385
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1958__A2
timestamp 1646674385
transform -1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_10
timestamp 1646674385
transform 1 0 2024 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1646674385
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1646674385
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1646674385
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2815_
timestamp 1646674385
transform -1 0 3864 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1646674385
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1646674385
transform 1 0 4232 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1646674385
transform 1 0 4692 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1452_
timestamp 1646674385
transform -1 0 4692 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1646674385
transform 1 0 5888 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1646674385
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2580_
timestamp 1646674385
transform -1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2835_
timestamp 1646674385
transform 1 0 6348 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1806__B2
timestamp 1646674385
transform -1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_73
timestamp 1646674385
transform 1 0 7820 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1646674385
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_101
timestamp 1646674385
transform 1 0 10396 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2633_
timestamp 1646674385
transform 1 0 8924 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1646674385
transform 1 0 11040 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1646674385
transform 1 0 11500 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1646674385
transform 1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1646674385
transform 1 0 12604 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1646674385
transform 1 0 11408 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1826_
timestamp 1646674385
transform 1 0 12236 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2231_
timestamp 1646674385
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2522_
timestamp 1646674385
transform -1 0 11868 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1808__A
timestamp 1646674385
transform -1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1646674385
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1646674385
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1831_
timestamp 1646674385
transform 1 0 13524 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1646674385
transform 1 0 16192 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2772_
timestamp 1646674385
transform 1 0 14720 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1646674385
transform 1 0 17572 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_183
timestamp 1646674385
transform 1 0 17940 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1646674385
transform 1 0 16560 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1567_
timestamp 1646674385
transform -1 0 17572 0 -1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2775_
timestamp 1646674385
transform 1 0 18032 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_17_200
timestamp 1646674385
transform 1 0 19504 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1851_
timestamp 1646674385
transform -1 0 20332 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1646674385
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1646674385
transform 1 0 20976 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1646674385
transform 1 0 21712 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2520_
timestamp 1646674385
transform 1 0 20700 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2565_
timestamp 1646674385
transform 1 0 21804 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_233
timestamp 1646674385
transform 1 0 22540 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_239
timestamp 1646674385
transform 1 0 23092 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_243
timestamp 1646674385
transform 1 0 23460 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1854_
timestamp 1646674385
transform 1 0 23184 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2437_
timestamp 1646674385
transform 1 0 24012 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_252
timestamp 1646674385
transform 1 0 24288 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1646674385
transform 1 0 25116 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2452_
timestamp 1646674385
transform 1 0 24656 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2475_
timestamp 1646674385
transform 1 0 25484 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1646674385
transform 1 0 26128 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1646674385
transform 1 0 26864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2739_
timestamp 1646674385
transform -1 0 28428 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2377__B2
timestamp 1646674385
transform 1 0 28796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_297
timestamp 1646674385
transform 1 0 28428 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_303
timestamp 1646674385
transform 1 0 28980 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2784_
timestamp 1646674385
transform 1 0 29532 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1646674385
transform 1 0 31004 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1646674385
transform -1 0 32016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_10
timestamp 1646674385
transform 1 0 2024 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1646674385
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1646674385
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1482_
timestamp 1646674385
transform -1 0 3312 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1916_
timestamp 1646674385
transform -1 0 2024 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1646674385
transform 1 0 3312 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_33
timestamp 1646674385
transform 1 0 4140 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1646674385
transform 1 0 3680 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1958_
timestamp 1646674385
transform 1 0 4508 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1959_
timestamp 1646674385
transform 1 0 3772 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1646674385
transform 1 0 5244 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 1646674385
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_59
timestamp 1646674385
transform 1 0 6532 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1451_
timestamp 1646674385
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_66
timestamp 1646674385
transform 1 0 7176 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_70
timestamp 1646674385
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1646674385
transform 1 0 8464 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1809_
timestamp 1646674385
transform -1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1955_
timestamp 1646674385
transform -1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp 1646674385
transform 1 0 10396 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_95
timestamp 1646674385
transform 1 0 9844 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1646674385
transform 1 0 8832 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1808_
timestamp 1646674385
transform -1 0 9844 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_2  _2636_
timestamp 1646674385
transform -1 0 12052 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1646674385
transform 1 0 12052 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2213_
timestamp 1646674385
transform -1 0 12696 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_126
timestamp 1646674385
transform 1 0 12696 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 1646674385
transform 1 0 13248 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1646674385
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1646674385
transform 1 0 13984 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2521_
timestamp 1646674385
transform -1 0 13616 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2618_
timestamp 1646674385
transform 1 0 14076 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_157
timestamp 1646674385
transform 1 0 15548 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2773_
timestamp 1646674385
transform 1 0 16100 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1646674385
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1564_
timestamp 1646674385
transform 1 0 17940 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1646674385
transform 1 0 18768 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1646674385
transform 1 0 19688 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1646674385
transform 1 0 19136 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1849_
timestamp 1646674385
transform 1 0 19228 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2608_
timestamp 1646674385
transform 1 0 20056 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_222
timestamp 1646674385
transform 1 0 21528 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2564_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 22080 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1646674385
transform 1 0 22632 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_238
timestamp 1646674385
transform 1 0 23000 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_244
timestamp 1646674385
transform 1 0 23552 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1853_
timestamp 1646674385
transform 1 0 23092 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1882__A_N
timestamp 1646674385
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1646674385
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1646674385
transform 1 0 25392 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1646674385
transform 1 0 24288 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2454_
timestamp 1646674385
transform 1 0 24932 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2457_
timestamp 1646674385
transform 1 0 25760 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_18_273
timestamp 1646674385
transform 1 0 26220 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1646674385
transform 1 0 26864 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1618_
timestamp 1646674385
transform 1 0 27232 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _2562_
timestamp 1646674385
transform 1 0 26588 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__A
timestamp 1646674385
transform 1 0 28520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1646674385
transform 1 0 28152 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1646674385
transform 1 0 28704 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1646674385
transform 1 0 29440 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2783_
timestamp 1646674385
transform 1 0 29532 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_325
timestamp 1646674385
transform 1 0 31004 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1646674385
transform -1 0 32016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1488_
timestamp 1646674385
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1487_
timestamp 1646674385
transform -1 0 2576 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1646674385
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1646674385
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1646674385
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1646674385
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1646674385
transform 1 0 2760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1646674385
transform 1 0 2392 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_16
timestamp 1646674385
transform 1 0 2576 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1490_
timestamp 1646674385
transform -1 0 3772 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_29
timestamp 1646674385
transform 1 0 3772 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1646674385
transform 1 0 4508 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1646674385
transform 1 0 3128 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1646674385
transform 1 0 3772 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1646674385
transform 1 0 3680 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_2  _1957_
timestamp 1646674385
transform 1 0 4600 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_prog_clk
timestamp 1646674385
transform 1 0 4140 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1646674385
transform 1 0 5520 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_62
timestamp 1646674385
transform 1 0 6808 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_53
timestamp 1646674385
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1646674385
transform 1 0 6624 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1646674385
transform 1 0 6256 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1918_
timestamp 1646674385
transform -1 0 6624 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1956_
timestamp 1646674385
transform -1 0 6808 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1646674385
transform 1 0 8464 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2837_
timestamp 1646674385
transform 1 0 6992 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2838_
timestamp 1646674385
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__o221a_1  _1806_
timestamp 1646674385
transform -1 0 10396 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1400_
timestamp 1646674385
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1646674385
transform 1 0 8832 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1646674385
transform 1 0 9200 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1646674385
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_92
timestamp 1646674385
transform 1 0 9568 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1646674385
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1804__B2
timestamp 1646674385
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_101
timestamp 1646674385
transform 1 0 10396 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1802_
timestamp 1646674385
transform 1 0 10120 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1834_
timestamp 1646674385
transform 1 0 11132 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1646674385
transform 1 0 11408 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1646674385
transform 1 0 11592 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1646674385
transform 1 0 11500 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1646674385
transform 1 0 11040 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1835_
timestamp 1646674385
transform -1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1646674385
transform 1 0 12236 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1646674385
transform 1 0 11868 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1802__A
timestamp 1646674385
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2616_
timestamp 1646674385
transform 1 0 11960 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_19_127
timestamp 1646674385
transform 1 0 12788 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1646674385
transform 1 0 13432 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_135
timestamp 1646674385
transform 1 0 13524 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__A
timestamp 1646674385
transform -1 0 13524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1646674385
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1646674385
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_145
timestamp 1646674385
transform 1 0 14444 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1646674385
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1646674385
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1646674385
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1646674385
transform 1 0 14996 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1646674385
transform 1 0 15732 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1646674385
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_161
timestamp 1646674385
transform 1 0 15916 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1302_
timestamp 1646674385
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1386_
timestamp 1646674385
transform 1 0 15364 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1566_
timestamp 1646674385
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1569_
timestamp 1646674385
transform -1 0 15916 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1389_
timestamp 1646674385
transform -1 0 17112 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1646674385
transform 1 0 16560 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_169
timestamp 1646674385
transform 1 0 16652 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1646674385
transform 1 0 17112 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1646674385
transform 1 0 16652 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1646674385
transform 1 0 16468 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1646674385
transform 1 0 18216 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1646674385
transform 1 0 17664 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__A
timestamp 1646674385
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2774_
timestamp 1646674385
transform 1 0 17480 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1561_
timestamp 1646674385
transform 1 0 16744 0 1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1561__A
timestamp 1646674385
transform -1 0 18768 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1646674385
transform 1 0 18952 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1646674385
transform 1 0 18768 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1646674385
transform 1 0 20056 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1646674385
transform 1 0 19136 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1563_
timestamp 1646674385
transform 1 0 19228 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _2776_
timestamp 1646674385
transform 1 0 19320 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1646674385
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1646674385
transform 1 0 21620 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1646674385
transform 1 0 21804 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1646674385
transform 1 0 21160 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_229
timestamp 1646674385
transform 1 0 22172 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1646674385
transform 1 0 21712 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1601_
timestamp 1646674385
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _1870_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 20424 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1871_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 21528 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_19_232
timestamp 1646674385
transform 1 0 22448 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_236
timestamp 1646674385
transform 1 0 22816 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_237
timestamp 1646674385
transform 1 0 22908 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1646674385
transform 1 0 23920 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1838_
timestamp 1646674385
transform 1 0 23000 0 1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2607_
timestamp 1646674385
transform 1 0 22908 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 1646674385
transform 1 0 24380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_265
timestamp 1646674385
transform 1 0 25484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_260
timestamp 1646674385
transform 1 0 25024 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_266
timestamp 1646674385
transform 1 0 25576 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1646674385
transform 1 0 24288 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _1882_
timestamp 1646674385
transform -1 0 25484 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1883_
timestamp 1646674385
transform -1 0 25024 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2560_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 26128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2561_
timestamp 1646674385
transform -1 0 26404 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_275
timestamp 1646674385
transform 1 0 26404 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1646674385
transform 1 0 26128 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2547_
timestamp 1646674385
transform -1 0 27232 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2546_
timestamp 1646674385
transform 1 0 27140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2545_
timestamp 1646674385
transform -1 0 27876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1646674385
transform 1 0 26864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_284
timestamp 1646674385
transform 1 0 27232 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1646674385
transform 1 0 26956 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1646674385
transform 1 0 27876 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_291
timestamp 1646674385
transform 1 0 27876 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1646674385
transform 1 0 29072 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1646674385
transform 1 0 29440 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1551_
timestamp 1646674385
transform 1 0 29532 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1553_
timestamp 1646674385
transform 1 0 28244 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_prog_clk
timestamp 1646674385
transform 1 0 28244 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1646674385
transform 1 0 30360 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_315
timestamp 1646674385
transform 1 0 30084 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2378__C
timestamp 1646674385
transform -1 0 30636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1646674385
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2543_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 31372 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_322
timestamp 1646674385
transform 1 0 30728 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_325
timestamp 1646674385
transform 1 0 31004 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_321
timestamp 1646674385
transform 1 0 30636 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1646674385
transform -1 0 32016 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1646674385
transform -1 0 32016 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_329
timestamp 1646674385
transform 1 0 31372 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_329
timestamp 1646674385
transform 1 0 31372 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__A1
timestamp 1646674385
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1646674385
transform 1 0 2484 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1646674385
transform 1 0 2760 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_7
timestamp 1646674385
transform 1 0 1748 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1646674385
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1646674385
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__B2
timestamp 1646674385
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1646674385
transform 1 0 3312 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_31
timestamp 1646674385
transform 1 0 3956 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1942_
timestamp 1646674385
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _1962_
timestamp 1646674385
transform -1 0 5888 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1646674385
transform 1 0 5888 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1646674385
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1646674385
transform 1 0 6256 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1443_
timestamp 1646674385
transform -1 0 7360 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_21_68
timestamp 1646674385
transform 1 0 7360 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_76
timestamp 1646674385
transform 1 0 8096 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_81
timestamp 1646674385
transform 1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1445_
timestamp 1646674385
transform -1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__A
timestamp 1646674385
transform 1 0 9568 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__A
timestamp 1646674385
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1646674385
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_91
timestamp 1646674385
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_94
timestamp 1646674385
transform 1 0 9752 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_98
timestamp 1646674385
transform 1 0 10120 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1804_
timestamp 1646674385
transform 1 0 10212 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1646674385
transform 1 0 11040 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1646674385
transform 1 0 11500 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1646674385
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1646674385
transform 1 0 11408 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1833_
timestamp 1646674385
transform 1 0 11868 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_21_133
timestamp 1646674385
transform 1 0 13340 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1993_
timestamp 1646674385
transform 1 0 12696 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2909_
timestamp 1646674385
transform 1 0 14076 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__A
timestamp 1646674385
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1646674385
transform 1 0 15548 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1646674385
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1566__A
timestamp 1646674385
transform -1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1646674385
transform 1 0 16468 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_171
timestamp 1646674385
transform 1 0 16836 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_177
timestamp 1646674385
transform 1 0 17388 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_187
timestamp 1646674385
transform 1 0 18308 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1646674385
transform 1 0 16560 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1565_
timestamp 1646674385
transform -1 0 18308 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1831__B1
timestamp 1646674385
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_193
timestamp 1646674385
transform 1 0 18860 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1646674385
transform 1 0 20056 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1850_
timestamp 1646674385
transform 1 0 19596 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__A
timestamp 1646674385
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1849__B
timestamp 1646674385
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_212
timestamp 1646674385
transform 1 0 20608 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1646674385
transform 1 0 21344 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1646674385
transform 1 0 21712 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1872_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 21804 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1646674385
transform 1 0 23000 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_242
timestamp 1646674385
transform 1 0 23368 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_249
timestamp 1646674385
transform 1 0 24012 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1884_
timestamp 1646674385
transform 1 0 23460 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_255
timestamp 1646674385
transform 1 0 24564 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2794_
timestamp 1646674385
transform -1 0 26128 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1883__B
timestamp 1646674385
transform -1 0 27968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1646674385
transform 1 0 26128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1646674385
transform 1 0 27416 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1646674385
transform 1 0 26864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _2556_
timestamp 1646674385
transform 1 0 26956 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_21_292
timestamp 1646674385
transform 1 0 27968 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_299
timestamp 1646674385
transform 1 0 28612 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_305
timestamp 1646674385
transform 1 0 29164 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_309
timestamp 1646674385
transform 1 0 29532 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2540_
timestamp 1646674385
transform 1 0 29256 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2544_
timestamp 1646674385
transform -1 0 28612 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_329
timestamp 1646674385
transform 1 0 31372 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1646674385
transform -1 0 32016 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2781_
timestamp 1646674385
transform 1 0 29900 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1646674385
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1646674385
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1646674385
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2819_
timestamp 1646674385
transform 1 0 1840 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1646674385
transform 1 0 3312 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1646674385
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1646674385
transform 1 0 4140 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_37
timestamp 1646674385
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1646674385
transform 1 0 3680 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1917_
timestamp 1646674385
transform -1 0 4508 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1939_
timestamp 1646674385
transform -1 0 5152 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_44
timestamp 1646674385
transform 1 0 5152 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_56
timestamp 1646674385
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1446_
timestamp 1646674385
transform 1 0 6624 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1961_
timestamp 1646674385
transform -1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1646674385
transform 1 0 7452 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_76
timestamp 1646674385
transform 1 0 8096 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1954_
timestamp 1646674385
transform 1 0 7820 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_101
timestamp 1646674385
transform 1 0 10396 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1646674385
transform 1 0 8832 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2634_
timestamp 1646674385
transform 1 0 8924 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_114
timestamp 1646674385
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1803_
timestamp 1646674385
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_4  _1994_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 12328 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1646674385
transform 1 0 13616 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1646674385
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1646674385
transform 1 0 13984 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1305_
timestamp 1646674385
transform -1 0 15088 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_22_152
timestamp 1646674385
transform 1 0 15088 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2910_
timestamp 1646674385
transform -1 0 17112 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1569__A
timestamp 1646674385
transform 1 0 18124 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1646674385
transform 1 0 17112 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1646674385
transform 1 0 17756 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1646674385
transform 1 0 18308 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2485_
timestamp 1646674385
transform 1 0 17480 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1646674385
transform 1 0 19044 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_206
timestamp 1646674385
transform 1 0 20056 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1646674385
transform 1 0 19136 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1562_
timestamp 1646674385
transform 1 0 19228 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1529__B1
timestamp 1646674385
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1884__B1
timestamp 1646674385
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_214
timestamp 1646674385
transform 1 0 20792 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1646674385
transform 1 0 21344 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_229
timestamp 1646674385
transform 1 0 22172 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1839_
timestamp 1646674385
transform 1 0 21712 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1872__B1
timestamp 1646674385
transform 1 0 23552 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_240
timestamp 1646674385
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1646674385
transform 1 0 23736 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  _1873_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 23184 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_22_262
timestamp 1646674385
transform 1 0 25208 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1646674385
transform 1 0 24288 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _1885_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 24380 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _2536_
timestamp 1646674385
transform 1 0 25760 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_272
timestamp 1646674385
transform 1 0 26128 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_284
timestamp 1646674385
transform 1 0 27232 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2558_
timestamp 1646674385
transform 1 0 26680 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2786_
timestamp 1646674385
transform 1 0 27600 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1646674385
transform 1 0 29072 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_309
timestamp 1646674385
transform 1 0 29532 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1646674385
transform 1 0 29440 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1555_
timestamp 1646674385
transform 1 0 29624 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_319
timestamp 1646674385
transform 1 0 30452 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1646674385
transform 1 0 31280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_332
timestamp 1646674385
transform 1 0 31648 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1646674385
transform -1 0 32016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2541_
timestamp 1646674385
transform -1 0 31280 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_23_19
timestamp 1646674385
transform 1 0 2852 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1646674385
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2818_
timestamp 1646674385
transform -1 0 2852 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp 1646674385
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 1646674385
transform 1 0 4692 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1485_
timestamp 1646674385
transform -1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1940_
timestamp 1646674385
transform -1 0 4692 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2008__A2
timestamp 1646674385
transform -1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_46
timestamp 1646674385
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1646674385
transform 1 0 5888 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1646674385
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1646674385
transform 1 0 6256 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1447_
timestamp 1646674385
transform 1 0 6532 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1941_
timestamp 1646674385
transform 1 0 5060 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1804__C1
timestamp 1646674385
transform -1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 1646674385
transform 1 0 7360 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_75
timestamp 1646674385
transform 1 0 8004 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 1646674385
transform 1 0 8556 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1892_
timestamp 1646674385
transform -1 0 8004 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1803__C1
timestamp 1646674385
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1646674385
transform 1 0 10580 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1646674385
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_90
timestamp 1646674385
transform 1 0 9384 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1805_
timestamp 1646674385
transform -1 0 10580 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1646674385
transform 1 0 11316 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1646674385
transform 1 0 11408 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2637_
timestamp 1646674385
transform 1 0 11500 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_129
timestamp 1646674385
transform 1 0 12972 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1646674385
transform 1 0 13708 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1646674385
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1290_
timestamp 1646674385
transform 1 0 13340 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1992_
timestamp 1646674385
transform -1 0 14352 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1646674385
transform 1 0 16192 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2907_
timestamp 1646674385
transform -1 0 16192 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1646674385
transform 1 0 17480 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1646674385
transform 1 0 16560 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1304_
timestamp 1646674385
transform -1 0 17480 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2898_
timestamp 1646674385
transform -1 0 19320 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1832__A
timestamp 1646674385
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2158__A2
timestamp 1646674385
transform -1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1646674385
transform 1 0 19320 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_204
timestamp 1646674385
transform 1 0 19872 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1529__A1
timestamp 1646674385
transform -1 0 21344 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_210
timestamp 1646674385
transform 1 0 20424 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1646674385
transform 1 0 21344 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1646674385
transform 1 0 21804 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1646674385
transform 1 0 21712 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1847_
timestamp 1646674385
transform 1 0 22172 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1842__A
timestamp 1646674385
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_234
timestamp 1646674385
transform 1 0 22632 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_242
timestamp 1646674385
transform 1 0 23368 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1646674385
transform 1 0 23644 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2793_
timestamp 1646674385
transform -1 0 25484 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1646674385
transform 1 0 25484 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2559_
timestamp 1646674385
transform 1 0 25852 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2186__C
timestamp 1646674385
transform 1 0 27692 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1646674385
transform 1 0 26128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_285
timestamp 1646674385
transform 1 0 27324 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_291
timestamp 1646674385
transform 1 0 27876 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1646674385
transform 1 0 26864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _2557_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 27324 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_295
timestamp 1646674385
transform 1 0 28244 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_312
timestamp 1646674385
transform 1 0 29808 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2785_
timestamp 1646674385
transform -1 0 29808 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_324
timestamp 1646674385
transform 1 0 30912 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_332
timestamp 1646674385
transform 1 0 31648 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1646674385
transform -1 0 32016 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2542_
timestamp 1646674385
transform 1 0 30544 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2157__A2
timestamp 1646674385
transform -1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_18
timestamp 1646674385
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_5
timestamp 1646674385
transform 1 0 1564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1646674385
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1484_
timestamp 1646674385
transform -1 0 2760 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A
timestamp 1646674385
transform -1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1646674385
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_37
timestamp 1646674385
transform 1 0 4508 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1646674385
transform 1 0 3680 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2009_
timestamp 1646674385
transform -1 0 4508 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1646674385
transform 1 0 5428 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1450_
timestamp 1646674385
transform -1 0 5428 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2836_
timestamp 1646674385
transform 1 0 5796 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__B1
timestamp 1646674385
transform -1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 1646674385
transform 1 0 7268 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_74
timestamp 1646674385
transform 1 0 7912 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1646674385
transform 1 0 8464 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1891_
timestamp 1646674385
transform 1 0 7636 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1646674385
transform 1 0 9200 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1646674385
transform 1 0 8832 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2155_
timestamp 1646674385
transform 1 0 8924 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2635_
timestamp 1646674385
transform 1 0 9568 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1803__B2
timestamp 1646674385
transform -1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1805__C1
timestamp 1646674385
transform -1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 1646674385
transform 1 0 11040 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1646674385
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_120
timestamp 1646674385
transform 1 0 12144 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A
timestamp 1646674385
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_126
timestamp 1646674385
transform 1 0 12696 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1646674385
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_143
timestamp 1646674385
transform 1 0 14260 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1646674385
transform 1 0 13984 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1415_
timestamp 1646674385
transform 1 0 12788 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_159
timestamp 1646674385
transform 1 0 15732 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1303_
timestamp 1646674385
transform -1 0 15732 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1646674385
transform 1 0 16468 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_177
timestamp 1646674385
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2486_
timestamp 1646674385
transform 1 0 16560 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2488_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 17756 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1646674385
transform 1 0 18400 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1646674385
transform 1 0 19228 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1646674385
transform 1 0 19136 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2777_
timestamp 1646674385
transform 1 0 19504 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1646674385
transform 1 0 20976 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_228
timestamp 1646674385
transform 1 0 22080 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1529_
timestamp 1646674385
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1646674385
transform 1 0 23000 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1646674385
transform 1 0 23644 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1528_
timestamp 1646674385
transform 1 0 22448 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1848_
timestamp 1646674385
transform 1 0 23368 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1646674385
transform 1 0 24196 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_262
timestamp 1646674385
transform 1 0 25208 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1646674385
transform 1 0 24288 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1536_
timestamp 1646674385
transform 1 0 24380 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2791_
timestamp 1646674385
transform 1 0 25760 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_24_284
timestamp 1646674385
transform 1 0 27232 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_290
timestamp 1646674385
transform 1 0 27784 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1547_
timestamp 1646674385
transform -1 0 28704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2187__B1
timestamp 1646674385
transform 1 0 29532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1646674385
transform 1 0 28704 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_311
timestamp 1646674385
transform 1 0 29716 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1646674385
transform 1 0 29440 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_318
timestamp 1646674385
transform 1 0 30360 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_326
timestamp 1646674385
transform 1 0 31096 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_332
timestamp 1646674385
transform 1 0 31648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1646674385
transform -1 0 32016 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2537_
timestamp 1646674385
transform 1 0 30728 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output34
timestamp 1646674385
transform -1 0 30360 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_17
timestamp 1646674385
transform 1 0 2668 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1646674385
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1646674385
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1483_
timestamp 1646674385
transform -1 0 2668 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_25_21
timestamp 1646674385
transform 1 0 3036 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1646674385
transform 1 0 3864 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _2008_
timestamp 1646674385
transform -1 0 5152 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _2011_
timestamp 1646674385
transform -1 0 3864 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_44
timestamp 1646674385
transform 1 0 5152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1646674385
transform 1 0 5888 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1646674385
transform 1 0 6256 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1439_
timestamp 1646674385
transform 1 0 5520 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1448_
timestamp 1646674385
transform -1 0 7176 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1646674385
transform 1 0 7176 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_73
timestamp 1646674385
transform 1 0 7820 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1890_
timestamp 1646674385
transform -1 0 7820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2586_
timestamp 1646674385
transform -1 0 9016 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A
timestamp 1646674385
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1805__B2
timestamp 1646674385
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1646674385
transform 1 0 9016 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1646674385
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1646674385
transform 1 0 10212 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1893_
timestamp 1646674385
transform 1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1826__A
timestamp 1646674385
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1833__B
timestamp 1646674385
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1646674385
transform 1 0 10764 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1646674385
transform 1 0 11316 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1646674385
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_121
timestamp 1646674385
transform 1 0 12236 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1646674385
transform 1 0 11408 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1646674385
transform 1 0 12972 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2846_
timestamp 1646674385
transform 1 0 13064 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1646674385
transform 1 0 14536 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1646674385
transform 1 0 15732 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1307_
timestamp 1646674385
transform 1 0 14904 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1646674385
transform 1 0 16468 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1646674385
transform 1 0 17296 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_180
timestamp 1646674385
transform 1 0 17664 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1646674385
transform 1 0 16560 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _2487_
timestamp 1646674385
transform 1 0 16652 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2897_
timestamp 1646674385
transform 1 0 17756 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_197
timestamp 1646674385
transform 1 0 19228 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2617_
timestamp 1646674385
transform 1 0 19780 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1646674385
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1646674385
transform 1 0 21620 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_228
timestamp 1646674385
transform 1 0 22080 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1646674385
transform 1 0 21712 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1527_
timestamp 1646674385
transform -1 0 22080 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1646674385
transform 1 0 24104 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2609_
timestamp 1646674385
transform 1 0 22632 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_263
timestamp 1646674385
transform 1 0 25300 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1534_
timestamp 1646674385
transform 1 0 24472 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1538_
timestamp 1646674385
transform 1 0 25668 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2179__B
timestamp 1646674385
transform -1 0 27784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1646674385
transform 1 0 26496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_284
timestamp 1646674385
transform 1 0 27232 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_290
timestamp 1646674385
transform 1 0 27784 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1646674385
transform 1 0 26864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2555_
timestamp 1646674385
transform 1 0 26956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_296
timestamp 1646674385
transform 1 0 28336 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_306
timestamp 1646674385
transform 1 0 29256 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1549_
timestamp 1646674385
transform 1 0 28428 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1554_
timestamp 1646674385
transform 1 0 29624 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_319
timestamp 1646674385
transform 1 0 30452 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_329
timestamp 1646674385
transform 1 0 31372 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1646674385
transform -1 0 32016 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2539_
timestamp 1646674385
transform -1 0 31372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1646674385
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1646674385
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1646674385
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1646674385
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_6
timestamp 1646674385
transform 1 0 1656 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1646674385
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2007__B
timestamp 1646674385
transform -1 0 1656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_11
timestamp 1646674385
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_20
timestamp 1646674385
transform 1 0 2944 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2820_
timestamp 1646674385
transform 1 0 2208 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1480_
timestamp 1646674385
transform -1 0 2944 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1646674385
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_35
timestamp 1646674385
transform 1 0 4324 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_28
timestamp 1646674385
transform 1 0 3680 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1646674385
transform 1 0 4876 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1646674385
transform 1 0 3680 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _2007_
timestamp 1646674385
transform 1 0 3864 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _2013_
timestamp 1646674385
transform 1 0 4692 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2584_
timestamp 1646674385
transform -1 0 4876 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_56
timestamp 1646674385
transform 1 0 6256 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1646674385
transform 1 0 5612 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1646674385
transform 1 0 6164 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1646674385
transform 1 0 6348 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1646674385
transform 1 0 6256 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _2012_
timestamp 1646674385
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2156_
timestamp 1646674385
transform 1 0 6624 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1646674385
transform 1 0 7360 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1646674385
transform 1 0 8464 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_65
timestamp 1646674385
transform 1 0 7084 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_77
timestamp 1646674385
transform 1 0 8188 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2158_
timestamp 1646674385
transform -1 0 8464 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2159_
timestamp 1646674385
transform 1 0 8556 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2160_
timestamp 1646674385
transform 1 0 7452 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2161_
timestamp 1646674385
transform 1 0 6992 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1800__A
timestamp 1646674385
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1646674385
transform 1 0 9108 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_95
timestamp 1646674385
transform 1 0 9844 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1646674385
transform 1 0 8924 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1646674385
transform 1 0 8832 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1409_
timestamp 1646674385
transform 1 0 10212 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1800_
timestamp 1646674385
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2852_
timestamp 1646674385
transform 1 0 9292 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_26_109
timestamp 1646674385
transform 1 0 11132 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1646674385
transform 1 0 11684 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1646674385
transform 1 0 10764 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1646674385
transform 1 0 11316 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1646674385
transform 1 0 11408 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1408_
timestamp 1646674385
transform 1 0 11776 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2849_
timestamp 1646674385
transform 1 0 11500 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1646674385
transform 1 0 12972 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_132
timestamp 1646674385
transform 1 0 13248 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_126
timestamp 1646674385
transform 1 0 12696 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2209_
timestamp 1646674385
transform 1 0 13340 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2198_
timestamp 1646674385
transform -1 0 13616 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1646674385
transform 1 0 13984 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_140
timestamp 1646674385
transform 1 0 13984 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1646674385
transform 1 0 13616 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_143
timestamp 1646674385
transform 1 0 14260 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A
timestamp 1646674385
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1306_
timestamp 1646674385
transform 1 0 14628 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_146
timestamp 1646674385
transform 1 0 14536 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_149
timestamp 1646674385
transform 1 0 14812 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1831__B2
timestamp 1646674385
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_prog_clk
timestamp 1646674385
transform 1 0 16192 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2480_
timestamp 1646674385
transform 1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1646674385
transform 1 0 16100 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1646674385
transform 1 0 15456 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_160
timestamp 1646674385
transform 1 0 15824 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 1646674385
transform 1 0 15548 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1646674385
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  _1291_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 17112 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1646674385
transform 1 0 16560 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1646674385
transform 1 0 16928 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1646674385
transform 1 0 16652 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1646674385
transform 1 0 16468 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_168
timestamp 1646674385
transform 1 0 16560 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A
timestamp 1646674385
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _2444_
timestamp 1646674385
transform -1 0 17572 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1646674385
transform 1 0 17572 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1646674385
transform 1 0 17664 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2446_
timestamp 1646674385
transform 1 0 18124 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1299_
timestamp 1646674385
transform -1 0 18308 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1646674385
transform 1 0 18308 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1646674385
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1646674385
transform 1 0 18768 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_200
timestamp 1646674385
transform 1 0 19504 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_200
timestamp 1646674385
transform 1 0 19504 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1646674385
transform 1 0 19136 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1832_
timestamp 1646674385
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2441_
timestamp 1646674385
transform 1 0 19872 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2442_
timestamp 1646674385
transform -1 0 21252 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__o221a_1  _2445_
timestamp 1646674385
transform 1 0 18676 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_26_211
timestamp 1646674385
transform 1 0 20516 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_217
timestamp 1646674385
transform 1 0 21068 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1646674385
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1646674385
transform 1 0 21620 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1646674385
transform 1 0 21804 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1646674385
transform 1 0 21712 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1843_
timestamp 1646674385
transform -1 0 22540 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2795_
timestamp 1646674385
transform 1 0 21160 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_234
timestamp 1646674385
transform 1 0 22632 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1646674385
transform 1 0 23276 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1646674385
transform 1 0 23920 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_233
timestamp 1646674385
transform 1 0 22540 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1646674385
transform 1 0 23644 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1419_
timestamp 1646674385
transform -1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1423_
timestamp 1646674385
transform -1 0 23644 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1842_
timestamp 1646674385
transform -1 0 23920 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1530_
timestamp 1646674385
transform 1 0 24380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1646674385
transform 1 0 24288 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_253
timestamp 1646674385
transform 1 0 24380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_256
timestamp 1646674385
transform 1 0 24656 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__B1
timestamp 1646674385
transform -1 0 25208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1537_
timestamp 1646674385
transform -1 0 26588 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_270
timestamp 1646674385
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_264
timestamp 1646674385
transform 1 0 25392 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_262
timestamp 1646674385
transform 1 0 25208 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__C1
timestamp 1646674385
transform -1 0 25944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1533_
timestamp 1646674385
transform 1 0 24472 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1646674385
transform 1 0 26864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1646674385
transform 1 0 26496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1646674385
transform 1 0 26588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2160__A2
timestamp 1646674385
transform -1 0 26496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1543_
timestamp 1646674385
transform 1 0 26956 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1646674385
transform 1 0 27784 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_289
timestamp 1646674385
transform 1 0 27692 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1646674385
transform 1 0 27140 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2164__B1
timestamp 1646674385
transform 1 0 27508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2163__C
timestamp 1646674385
transform 1 0 26956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1646674385
transform -1 0 28428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2569_
timestamp 1646674385
transform 1 0 28796 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1542_
timestamp 1646674385
transform -1 0 28520 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_298
timestamp 1646674385
transform 1 0 28520 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_297
timestamp 1646674385
transform 1 0 28428 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_293
timestamp 1646674385
transform 1 0 28060 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1646674385
transform 1 0 29440 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_309
timestamp 1646674385
transform 1 0 29532 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1646674385
transform 1 0 29072 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2782_
timestamp 1646674385
transform -1 0 31096 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1548_
timestamp 1646674385
transform 1 0 29256 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_26_326
timestamp 1646674385
transform 1 0 31096 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_332
timestamp 1646674385
transform 1 0 31648 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_316
timestamp 1646674385
transform 1 0 30176 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_322
timestamp 1646674385
transform 1 0 30728 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_328
timestamp 1646674385
transform 1 0 31280 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_332
timestamp 1646674385
transform 1 0 31648 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1646674385
transform -1 0 32016 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1646674385
transform -1 0 32016 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2538_
timestamp 1646674385
transform 1 0 30820 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_28_16
timestamp 1646674385
transform 1 0 2576 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1646674385
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1646674385
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1472_
timestamp 1646674385
transform -1 0 3312 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1473_
timestamp 1646674385
transform -1 0 2576 0 1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1646674385
transform 1 0 3312 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1646674385
transform 1 0 3772 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1646674385
transform 1 0 4508 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1646674385
transform 1 0 3680 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1479_
timestamp 1646674385
transform 1 0 4140 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2010_
timestamp 1646674385
transform -1 0 5244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2010__A2
timestamp 1646674385
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 1646674385
transform 1 0 5244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_51
timestamp 1646674385
transform 1 0 5796 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1444_
timestamp 1646674385
transform 1 0 6164 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_64
timestamp 1646674385
transform 1 0 6992 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1646674385
transform 1 0 8464 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _2157_
timestamp 1646674385
transform 1 0 7544 0 1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_28_102
timestamp 1646674385
transform 1 0 10488 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1646674385
transform 1 0 8832 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_4  _2162_
timestamp 1646674385
transform 1 0 8924 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_28_106
timestamp 1646674385
transform 1 0 10856 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_116
timestamp 1646674385
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1410_
timestamp 1646674385
transform 1 0 10948 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2850_
timestamp 1646674385
transform 1 0 12144 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1646674385
transform 1 0 13616 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1646674385
transform 1 0 14076 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1646674385
transform 1 0 13984 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2908_
timestamp 1646674385
transform -1 0 15916 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1646674385
transform 1 0 15916 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _2483_
timestamp 1646674385
transform 1 0 16284 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_28_172
timestamp 1646674385
transform 1 0 16928 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1646674385
transform 1 0 18308 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1326_
timestamp 1646674385
transform 1 0 17480 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1646674385
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1646674385
transform 1 0 19228 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1646674385
transform 1 0 19136 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_prog_clk
timestamp 1646674385
transform 1 0 19596 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1646674385
transform 1 0 21436 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1646674385
transform 1 0 22080 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1844_
timestamp 1646674385
transform 1 0 21804 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1646674385
transform 1 0 23920 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2612_
timestamp 1646674385
transform -1 0 23920 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1646674385
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1646674385
transform 1 0 24840 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1646674385
transform 1 0 24288 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1531_
timestamp 1646674385
transform 1 0 24564 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2792_
timestamp 1646674385
transform 1 0 25208 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1646674385
transform 1 0 26680 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2789_
timestamp 1646674385
transform 1 0 27048 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__A
timestamp 1646674385
transform -1 0 29072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_298
timestamp 1646674385
transform 1 0 28520 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1646674385
transform 1 0 29072 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1646674385
transform 1 0 29532 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1646674385
transform 1 0 29440 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_317
timestamp 1646674385
transform 1 0 30268 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_324
timestamp 1646674385
transform 1 0 30912 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_332
timestamp 1646674385
transform 1 0 31648 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1646674385
transform -1 0 32016 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1550_
timestamp 1646674385
transform 1 0 29900 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2535_
timestamp 1646674385
transform 1 0 30636 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__A
timestamp 1646674385
transform -1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_18
timestamp 1646674385
transform 1 0 2760 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_5
timestamp 1646674385
transform 1 0 1564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1646674385
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1481_
timestamp 1646674385
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_26
timestamp 1646674385
transform 1 0 3496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_34
timestamp 1646674385
transform 1 0 4232 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_38
timestamp 1646674385
transform 1 0 4600 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1459_
timestamp 1646674385
transform 1 0 3128 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1463_
timestamp 1646674385
transform -1 0 4232 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2005_
timestamp 1646674385
transform 1 0 4692 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_42
timestamp 1646674385
transform 1 0 4968 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1646674385
transform 1 0 5704 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1646674385
transform 1 0 6256 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1442_
timestamp 1646674385
transform 1 0 5336 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2839_
timestamp 1646674385
transform -1 0 7912 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_29_74
timestamp 1646674385
transform 1 0 7912 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_82
timestamp 1646674385
transform 1 0 8648 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2154_
timestamp 1646674385
transform -1 0 9016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_86
timestamp 1646674385
transform 1 0 9016 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1646674385
transform 1 0 9752 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1512_
timestamp 1646674385
transform 1 0 9384 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2163_
timestamp 1646674385
transform 1 0 10120 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1646674385
transform 1 0 10764 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1646674385
transform 1 0 11316 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_123
timestamp 1646674385
transform 1 0 12420 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1646674385
transform 1 0 11408 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1406_
timestamp 1646674385
transform 1 0 11500 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1646674385
transform 1 0 13156 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_141
timestamp 1646674385
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_145
timestamp 1646674385
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2199_
timestamp 1646674385
transform 1 0 13248 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_150
timestamp 1646674385
transform 1 0 14904 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_154
timestamp 1646674385
transform 1 0 15272 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1646674385
transform 1 0 16192 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1301_
timestamp 1646674385
transform -1 0 14904 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2481_
timestamp 1646674385
transform 1 0 15364 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_185
timestamp 1646674385
transform 1 0 18124 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1646674385
transform 1 0 16560 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2900_
timestamp 1646674385
transform 1 0 16652 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_198
timestamp 1646674385
transform 1 0 19320 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_202
timestamp 1646674385
transform 1 0 19688 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1325_
timestamp 1646674385
transform 1 0 18492 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2895_
timestamp 1646674385
transform 1 0 19780 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1646674385
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1646674385
transform 1 0 21620 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1646674385
transform 1 0 21712 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _1426_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 22264 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__A
timestamp 1646674385
transform -1 0 23920 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_230
timestamp 1646674385
transform 1 0 22264 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_242
timestamp 1646674385
transform 1 0 23368 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_248
timestamp 1646674385
transform 1 0 23920 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1424_
timestamp 1646674385
transform 1 0 22632 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_262
timestamp 1646674385
transform 1 0 25208 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1532_
timestamp 1646674385
transform 1 0 25576 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1539_
timestamp 1646674385
transform 1 0 24288 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__B1
timestamp 1646674385
transform -1 0 27140 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1646674385
transform 1 0 26496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_283
timestamp 1646674385
transform 1 0 27140 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp 1646674385
transform 1 0 27508 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1646674385
transform 1 0 26864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1540_
timestamp 1646674385
transform 1 0 27600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_292
timestamp 1646674385
transform 1 0 27968 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1646674385
transform 1 0 28520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_305
timestamp 1646674385
transform 1 0 29164 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1557_
timestamp 1646674385
transform 1 0 29532 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2554_
timestamp 1646674385
transform -1 0 29164 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_318
timestamp 1646674385
transform 1 0 30360 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_329
timestamp 1646674385
transform 1 0 31372 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1646674385
transform -1 0 32016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2566_
timestamp 1646674385
transform 1 0 31096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2156__B
timestamp 1646674385
transform -1 0 1656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_14
timestamp 1646674385
transform 1 0 2392 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1646674385
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_6
timestamp 1646674385
transform 1 0 1656 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1646674385
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1470_
timestamp 1646674385
transform -1 0 2392 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1646674385
transform 1 0 2760 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A
timestamp 1646674385
transform -1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1646674385
transform 1 0 3128 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1646674385
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1646674385
transform 1 0 4232 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_41
timestamp 1646674385
transform 1 0 4876 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1646674385
transform 1 0 3680 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2006_
timestamp 1646674385
transform 1 0 4600 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _2031_
timestamp 1646674385
transform -1 0 6992 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2153__A2
timestamp 1646674385
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_64
timestamp 1646674385
transform 1 0 6992 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_71
timestamp 1646674385
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_77
timestamp 1646674385
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1646674385
transform 1 0 8464 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2249_
timestamp 1646674385
transform 1 0 7360 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A
timestamp 1646674385
transform -1 0 9568 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1646674385
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1646674385
transform 1 0 9292 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_92
timestamp 1646674385
transform 1 0 9568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1646674385
transform 1 0 8832 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2153_
timestamp 1646674385
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_105
timestamp 1646674385
transform 1 0 10764 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1646674385
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1411_
timestamp 1646674385
transform 1 0 11132 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1412_
timestamp 1646674385
transform 1 0 12328 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 1646674385
transform 1 0 13156 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1646674385
transform 1 0 13892 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1646674385
transform 1 0 13984 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _2164_
timestamp 1646674385
transform 1 0 14076 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1646674385
transform 1 0 14720 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1646674385
transform 1 0 15732 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_163
timestamp 1646674385
transform 1 0 16100 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1399_
timestamp 1646674385
transform 1 0 16192 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _2210_
timestamp 1646674385
transform 1 0 15088 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_168
timestamp 1646674385
transform 1 0 16560 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1646674385
transform 1 0 17756 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1323_
timestamp 1646674385
transform -1 0 17756 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _2430_
timestamp 1646674385
transform 1 0 18124 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1646674385
transform 1 0 18768 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1646674385
transform 1 0 19136 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2447_
timestamp 1646674385
transform 1 0 19228 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1646674385
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2611_
timestamp 1646674385
transform 1 0 20792 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_230
timestamp 1646674385
transform 1 0 22264 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_238
timestamp 1646674385
transform 1 0 23000 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1646674385
transform 1 0 23920 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1560_
timestamp 1646674385
transform 1 0 23092 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_269
timestamp 1646674385
transform 1 0 25852 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1646674385
transform 1 0 24288 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2778_
timestamp 1646674385
transform -1 0 25852 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__A
timestamp 1646674385
transform 1 0 27508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_283
timestamp 1646674385
transform 1 0 27140 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_289
timestamp 1646674385
transform 1 0 27692 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1535_
timestamp 1646674385
transform 1 0 26220 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_30_293
timestamp 1646674385
transform 1 0 28060 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1646674385
transform 1 0 29072 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1646674385
transform 1 0 29440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1552_
timestamp 1646674385
transform 1 0 28152 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1556_
timestamp 1646674385
transform 1 0 29532 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_318
timestamp 1646674385
transform 1 0 30360 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_326
timestamp 1646674385
transform 1 0 31096 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_332
timestamp 1646674385
transform 1 0 31648 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1646674385
transform -1 0 32016 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2552_
timestamp 1646674385
transform 1 0 30728 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_12
timestamp 1646674385
transform 1 0 2208 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1646674385
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1476_
timestamp 1646674385
transform 1 0 1380 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2823_
timestamp 1646674385
transform 1 0 2576 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_32
timestamp 1646674385
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1646674385
transform 1 0 4784 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1475_
timestamp 1646674385
transform -1 0 4784 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp 1646674385
transform 1 0 5520 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1646674385
transform 1 0 6348 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1646674385
transform 1 0 6256 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1438_
timestamp 1646674385
transform -1 0 7084 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2028_
timestamp 1646674385
transform -1 0 5520 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A
timestamp 1646674385
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_65
timestamp 1646674385
transform 1 0 7084 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 1646674385
transform 1 0 7636 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_80
timestamp 1646674385
transform 1 0 8464 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2265_
timestamp 1646674385
transform 1 0 8004 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_31_94
timestamp 1646674385
transform 1 0 9752 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1405_
timestamp 1646674385
transform -1 0 10948 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1773_
timestamp 1646674385
transform -1 0 9752 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1646674385
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1646674385
transform 1 0 11316 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_116
timestamp 1646674385
transform 1 0 11776 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1646674385
transform 1 0 11408 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2152_
timestamp 1646674385
transform 1 0 11500 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2848_
timestamp 1646674385
transform 1 0 12328 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1646674385
transform 1 0 13800 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_prog_clk
timestamp 1646674385
transform 1 0 14168 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1646674385
transform 1 0 16008 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1646674385
transform 1 0 16652 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_182
timestamp 1646674385
transform 1 0 17848 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1646674385
transform 1 0 16560 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2429_
timestamp 1646674385
transform 1 0 17020 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1646674385
transform 1 0 18216 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1646674385
transform 1 0 20056 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1646674385
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1646674385
transform 1 0 21620 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1646674385
transform 1 0 21804 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1646674385
transform 1 0 22172 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1646674385
transform 1 0 21712 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2440_
timestamp 1646674385
transform 1 0 20424 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1646674385
transform 1 0 23828 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2845_
timestamp 1646674385
transform 1 0 22264 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_31_254
timestamp 1646674385
transform 1 0 24472 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2439_
timestamp 1646674385
transform 1 0 24196 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2738_
timestamp 1646674385
transform 1 0 25024 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1646674385
transform 1 0 26496 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_290
timestamp 1646674385
transform 1 0 27784 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1646674385
transform 1 0 26864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1541_
timestamp 1646674385
transform 1 0 26956 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_296
timestamp 1646674385
transform 1 0 28336 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_302
timestamp 1646674385
transform 1 0 28888 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_309
timestamp 1646674385
transform 1 0 29532 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2551_
timestamp 1646674385
transform 1 0 29256 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2553_
timestamp 1646674385
transform -1 0 28888 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_31_329
timestamp 1646674385
transform 1 0 31372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1646674385
transform -1 0 32016 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2779_
timestamp 1646674385
transform 1 0 29900 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1646674385
transform 1 0 2852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1646674385
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2822_
timestamp 1646674385
transform -1 0 2852 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2012__A2
timestamp 1646674385
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2026__A2
timestamp 1646674385
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1646674385
transform 1 0 3588 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 1646674385
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1646674385
transform 1 0 4048 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_38
timestamp 1646674385
transform 1 0 4600 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1646674385
transform 1 0 3680 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_46
timestamp 1646674385
transform 1 0 5336 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_55
timestamp 1646674385
transform 1 0 6164 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1646674385
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2023_
timestamp 1646674385
transform -1 0 6164 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2030_
timestamp 1646674385
transform -1 0 5336 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2248_
timestamp 1646674385
transform -1 0 7084 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_65
timestamp 1646674385
transform 1 0 7084 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1646674385
transform 1 0 8188 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1646674385
transform 1 0 8740 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2267_
timestamp 1646674385
transform -1 0 8188 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1773__A
timestamp 1646674385
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_88
timestamp 1646674385
transform 1 0 9200 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_96
timestamp 1646674385
transform 1 0 9936 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1646674385
transform 1 0 8832 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _2250_
timestamp 1646674385
transform 1 0 8924 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_prog_clk
timestamp 1646674385
transform 1 0 10488 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_32_122
timestamp 1646674385
transform 1 0 12328 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A
timestamp 1646674385
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__A
timestamp 1646674385
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_128
timestamp 1646674385
transform 1 0 12880 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1646674385
transform 1 0 13616 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_143
timestamp 1646674385
transform 1 0 14260 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1646674385
transform 1 0 13984 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1421_
timestamp 1646674385
transform -1 0 13616 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_153
timestamp 1646674385
transform 1 0 15180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1646674385
transform 1 0 16192 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1420_
timestamp 1646674385
transform 1 0 14628 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2482_
timestamp 1646674385
transform 1 0 15548 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1646674385
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp 1646674385
transform 1 0 17204 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1646674385
transform 1 0 17756 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _2431_
timestamp 1646674385
transform 1 0 18124 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2498_
timestamp 1646674385
transform 1 0 16560 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1646674385
transform 1 0 18768 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1646674385
transform 1 0 20056 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1646674385
transform 1 0 19136 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1331_
timestamp 1646674385
transform 1 0 19228 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__A
timestamp 1646674385
transform -1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1646674385
transform 1 0 20700 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1646674385
transform 1 0 21252 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_229
timestamp 1646674385
transform 1 0 22172 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1926_
timestamp 1646674385
transform 1 0 21620 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2428_
timestamp 1646674385
transform 1 0 20424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_235
timestamp 1646674385
transform 1 0 22724 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_240
timestamp 1646674385
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1646674385
transform 1 0 23920 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1418_
timestamp 1646674385
transform -1 0 23184 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1422_
timestamp 1646674385
transform -1 0 23920 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A
timestamp 1646674385
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_255
timestamp 1646674385
transform 1 0 24564 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1646674385
transform 1 0 24288 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_prog_clk
timestamp 1646674385
transform 1 0 25300 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_32_283
timestamp 1646674385
transform 1 0 27140 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2790_
timestamp 1646674385
transform 1 0 27508 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1646674385
transform 1 0 28980 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1646674385
transform 1 0 29348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1646674385
transform 1 0 29532 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1646674385
transform 1 0 29440 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_329
timestamp 1646674385
transform 1 0 31372 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1646674385
transform -1 0 32016 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2780_
timestamp 1646674385
transform 1 0 29900 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1875_
timestamp 1646674385
transform 1 0 1840 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1477_
timestamp 1646674385
transform 1 0 1472 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1646674385
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1646674385
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_7
timestamp 1646674385
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1646674385
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1646674385
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2172_
timestamp 1646674385
transform -1 0 3220 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1877_
timestamp 1646674385
transform -1 0 2944 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_11
timestamp 1646674385
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1646674385
transform 1 0 2300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_20
timestamp 1646674385
transform 1 0 2944 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_31
timestamp 1646674385
transform 1 0 3956 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_38
timestamp 1646674385
transform 1 0 4600 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1646674385
transform 1 0 3220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1646674385
transform 1 0 3588 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_38
timestamp 1646674385
transform 1 0 4600 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1646674385
transform 1 0 3680 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1902_
timestamp 1646674385
transform -1 0 4600 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2167_
timestamp 1646674385
transform -1 0 3956 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2579_
timestamp 1646674385
transform -1 0 4600 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_33_50
timestamp 1646674385
transform 1 0 5704 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_46
timestamp 1646674385
transform 1 0 5336 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_57
timestamp 1646674385
transform 1 0 6348 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1646674385
transform 1 0 6256 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _2025_
timestamp 1646674385
transform -1 0 7176 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _2026_
timestamp 1646674385
transform 1 0 5428 0 1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _2027_
timestamp 1646674385
transform 1 0 4968 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2590_
timestamp 1646674385
transform 1 0 6348 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_66
timestamp 1646674385
transform 1 0 7176 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_73
timestamp 1646674385
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_66
timestamp 1646674385
transform 1 0 7176 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1646674385
transform 1 0 8464 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2247_
timestamp 1646674385
transform -1 0 7820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _2266_
timestamp 1646674385
transform 1 0 7544 0 1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2587_
timestamp 1646674385
transform -1 0 9016 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1646674385
transform 1 0 9016 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_102
timestamp 1646674385
transform 1 0 10488 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1646674385
transform 1 0 8832 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_4  _2271_
timestamp 1646674385
transform -1 0 10488 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2851_
timestamp 1646674385
transform 1 0 9384 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2153__B2
timestamp 1646674385
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1646674385
transform 1 0 10856 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_115
timestamp 1646674385
transform 1 0 11684 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_115
timestamp 1646674385
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_119
timestamp 1646674385
transform 1 0 12052 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1646674385
transform 1 0 11408 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1407_
timestamp 1646674385
transform -1 0 11684 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1413_
timestamp 1646674385
transform 1 0 12144 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2847_
timestamp 1646674385
transform 1 0 12420 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2104__B1
timestamp 1646674385
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1646674385
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1646674385
transform 1 0 12972 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1646674385
transform 1 0 13340 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1646674385
transform 1 0 13616 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1646674385
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1646674385
transform 1 0 14444 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1646674385
transform 1 0 13984 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2906_
timestamp 1646674385
transform 1 0 14260 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1646674385
transform 1 0 15732 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1646674385
transform 1 0 15364 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1646674385
transform 1 0 16100 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1297_
timestamp 1646674385
transform -1 0 16100 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1311_
timestamp 1646674385
transform -1 0 15364 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2499_
timestamp 1646674385
transform -1 0 17296 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1328_
timestamp 1646674385
transform 1 0 16468 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1646674385
transform 1 0 16560 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1646674385
transform 1 0 17296 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_176
timestamp 1646674385
transform 1 0 17296 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1646674385
transform 1 0 16468 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1646674385
transform -1 0 17940 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1646674385
transform 1 0 17940 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2896_
timestamp 1646674385
transform 1 0 18308 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1296_
timestamp 1646674385
transform 1 0 17664 0 1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1646674385
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_203
timestamp 1646674385
transform 1 0 19780 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1646674385
transform 1 0 18584 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_199
timestamp 1646674385
transform 1 0 19412 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1646674385
transform 1 0 19136 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1333_
timestamp 1646674385
transform 1 0 20148 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2894_
timestamp 1646674385
transform -1 0 21620 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1646674385
transform 1 0 20976 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_228
timestamp 1646674385
transform 1 0 22080 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1646674385
transform 1 0 21620 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1646674385
transform 1 0 21712 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2381_
timestamp 1646674385
transform -1 0 22080 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2383_
timestamp 1646674385
transform 1 0 21988 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1840_
timestamp 1646674385
transform 1 0 22540 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1293_
timestamp 1646674385
transform -1 0 23368 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_238
timestamp 1646674385
transform 1 0 23000 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1646674385
transform 1 0 22632 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_236
timestamp 1646674385
transform 1 0 22816 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_232
timestamp 1646674385
transform 1 0 22448 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1629_
timestamp 1646674385
transform 1 0 23368 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1646674385
transform 1 0 23920 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_242
timestamp 1646674385
transform 1 0 23368 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A
timestamp 1646674385
transform 1 0 23736 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1627__A
timestamp 1646674385
transform 1 0 25852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_251
timestamp 1646674385
transform 1 0 24196 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_265
timestamp 1646674385
transform 1 0 25484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_263
timestamp 1646674385
transform 1 0 25300 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1646674385
transform 1 0 24288 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1627_
timestamp 1646674385
transform 1 0 24564 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1628_
timestamp 1646674385
transform 1 0 24380 0 1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1622_
timestamp 1646674385
transform -1 0 26404 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1646674385
transform 1 0 26864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_281
timestamp 1646674385
transform 1 0 26956 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_275
timestamp 1646674385
transform 1 0 26404 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1646674385
transform 1 0 26956 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1646674385
transform 1 0 26772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1646674385
transform 1 0 26036 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1546_
timestamp 1646674385
transform 1 0 27048 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1646674385
transform 1 0 27876 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_285
timestamp 1646674385
transform 1 0 27324 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1544__A
timestamp 1646674385
transform 1 0 27140 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2788_
timestamp 1646674385
transform -1 0 29164 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_305
timestamp 1646674385
transform 1 0 29164 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1646674385
transform 1 0 29072 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1646674385
transform 1 0 29440 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1545_
timestamp 1646674385
transform 1 0 28244 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2787_
timestamp 1646674385
transform 1 0 29532 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_prog_clk
timestamp 1646674385
transform 1 0 29532 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_33_325
timestamp 1646674385
transform 1 0 31004 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1646674385
transform 1 0 31372 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1646674385
transform -1 0 32016 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1646674385
transform -1 0 32016 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_9
timestamp 1646674385
transform 1 0 1932 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1646674385
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2170_
timestamp 1646674385
transform -1 0 3036 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1646674385
transform 1 0 1380 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1646674385
transform 1 0 3036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_35
timestamp 1646674385
transform 1 0 4324 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_41
timestamp 1646674385
transform 1 0 4876 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_2  _2169_
timestamp 1646674385
transform 1 0 3404 0 -1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1646674385
transform 1 0 5704 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_60
timestamp 1646674385
transform 1 0 6624 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1646674385
transform 1 0 6256 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1899_
timestamp 1646674385
transform -1 0 6624 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2029_
timestamp 1646674385
transform 1 0 4968 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2025__B
timestamp 1646674385
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_66
timestamp 1646674385
transform 1 0 7176 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_78
timestamp 1646674385
transform 1 0 8280 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2268_
timestamp 1646674385
transform 1 0 8648 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2269_
timestamp 1646674385
transform -1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1646674385
transform 1 0 9016 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_93
timestamp 1646674385
transform 1 0 9660 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _2186_
timestamp 1646674385
transform 1 0 10396 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2263_
timestamp 1646674385
transform 1 0 9384 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1646674385
transform 1 0 11040 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1646674385
transform 1 0 11500 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1646674385
transform 1 0 11408 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2187_
timestamp 1646674385
transform 1 0 11776 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1964__A
timestamp 1646674385
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_129
timestamp 1646674385
transform 1 0 12972 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_136
timestamp 1646674385
transform 1 0 13616 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_142
timestamp 1646674385
transform 1 0 14168 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2190_
timestamp 1646674385
transform 1 0 13340 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_151
timestamp 1646674385
transform 1 0 14996 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1646674385
transform 1 0 16192 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2496_
timestamp 1646674385
transform 1 0 14720 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2497_
timestamp 1646674385
transform 1 0 15364 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_35_169
timestamp 1646674385
transform 1 0 16652 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1646674385
transform 1 0 18216 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1646674385
transform 1 0 16560 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2899_
timestamp 1646674385
transform -1 0 18216 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_199
timestamp 1646674385
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_203
timestamp 1646674385
transform 1 0 19780 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1324_
timestamp 1646674385
transform 1 0 18584 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2893_
timestamp 1646674385
transform 1 0 19872 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1646674385
transform 1 0 21344 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1646674385
transform 1 0 21804 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1646674385
transform 1 0 21712 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2614_
timestamp 1646674385
transform 1 0 22172 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1628__A
timestamp 1646674385
transform 1 0 24012 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_245
timestamp 1646674385
transform 1 0 23644 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1646674385
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2734_
timestamp 1646674385
transform -1 0 26036 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1646674385
transform 1 0 26036 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1646674385
transform 1 0 26772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_291
timestamp 1646674385
transform 1 0 27876 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1646674385
transform 1 0 26864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1636_
timestamp 1646674385
transform -1 0 27876 0 -1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_35_299
timestamp 1646674385
transform 1 0 28612 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_306
timestamp 1646674385
transform 1 0 29256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1544_
timestamp 1646674385
transform -1 0 28612 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output35
timestamp 1646674385
transform -1 0 29256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1646674385
transform -1 0 30084 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_315
timestamp 1646674385
transform 1 0 30084 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_322
timestamp 1646674385
transform 1 0 30728 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_329
timestamp 1646674385
transform 1 0 31372 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1646674385
transform -1 0 32016 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2532_
timestamp 1646674385
transform -1 0 31372 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2570_
timestamp 1646674385
transform 1 0 30452 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2101__A2
timestamp 1646674385
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_16
timestamp 1646674385
transform 1 0 2576 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1646674385
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_9
timestamp 1646674385
transform 1 0 1932 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1646674385
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1874_
timestamp 1646674385
transform -1 0 2576 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2171_
timestamp 1646674385
transform -1 0 3312 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1646674385
transform 1 0 3312 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1646674385
transform 1 0 3680 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_4  _2174_
timestamp 1646674385
transform 1 0 3772 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_46
timestamp 1646674385
transform 1 0 5336 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_53
timestamp 1646674385
transform 1 0 5980 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_60
timestamp 1646674385
transform 1 0 6624 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1900_
timestamp 1646674385
transform -1 0 5980 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1901_
timestamp 1646674385
transform 1 0 6348 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_67
timestamp 1646674385
transform 1 0 7268 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_73
timestamp 1646674385
transform 1 0 7820 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1646674385
transform 1 0 8280 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2024_
timestamp 1646674385
transform 1 0 6992 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2270_
timestamp 1646674385
transform 1 0 7912 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_88
timestamp 1646674385
transform 1 0 9200 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1646674385
transform 1 0 8832 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2264_
timestamp 1646674385
transform 1 0 8924 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2854_
timestamp 1646674385
transform -1 0 11040 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_108
timestamp 1646674385
transform 1 0 11040 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_121
timestamp 1646674385
transform 1 0 12236 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1403_
timestamp 1646674385
transform -1 0 12236 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1646674385
transform 1 0 13432 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1646674385
transform 1 0 13984 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _2195_
timestamp 1646674385
transform 1 0 12788 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2905_
timestamp 1646674385
transform 1 0 14076 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_157
timestamp 1646674385
transform 1 0 15548 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1318_
timestamp 1646674385
transform 1 0 15916 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1646674385
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_170
timestamp 1646674385
transform 1 0 16744 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1646674385
transform 1 0 17296 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1321_
timestamp 1646674385
transform -1 0 18584 0 1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_36_190
timestamp 1646674385
transform 1 0 18584 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1646674385
transform 1 0 20148 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1646674385
transform 1 0 19136 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1327_
timestamp 1646674385
transform 1 0 19228 0 1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_36_220
timestamp 1646674385
transform 1 0 21344 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1332_
timestamp 1646674385
transform 1 0 20516 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2382_
timestamp 1646674385
transform 1 0 21712 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_36_233
timestamp 1646674385
transform 1 0 22540 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1646674385
transform 1 0 23920 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1633_
timestamp 1646674385
transform -1 0 23920 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1646674385
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_261
timestamp 1646674385
transform 1 0 25116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1646674385
transform 1 0 24288 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _1522_
timestamp 1646674385
transform 1 0 24564 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2733_
timestamp 1646674385
transform -1 0 26956 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_281
timestamp 1646674385
transform 1 0 26956 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2732_
timestamp 1646674385
transform 1 0 27324 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1646674385
transform 1 0 28796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1646674385
transform 1 0 29348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1646674385
transform 1 0 29532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1646674385
transform 1 0 29440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2548_
timestamp 1646674385
transform 1 0 29716 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_314
timestamp 1646674385
transform 1 0 29992 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_325
timestamp 1646674385
transform 1 0 31004 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1646674385
transform -1 0 32016 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2550_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 31004 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1646674385
transform 1 0 2116 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_15
timestamp 1646674385
transform 1 0 2484 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1646674385
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1646674385
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1876_
timestamp 1646674385
transform 1 0 2208 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2173_
timestamp 1646674385
transform 1 0 2852 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1646674385
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_23
timestamp 1646674385
transform 1 0 3220 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1646674385
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_39
timestamp 1646674385
transform 1 0 4692 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2166_
timestamp 1646674385
transform -1 0 4692 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2168_
timestamp 1646674385
transform 1 0 3588 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__A
timestamp 1646674385
transform -1 0 6532 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_47
timestamp 1646674385
transform 1 0 5428 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1646674385
transform 1 0 5888 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_59
timestamp 1646674385
transform 1 0 6532 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1646674385
transform 1 0 6256 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1508_
timestamp 1646674385
transform -1 0 5888 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_73
timestamp 1646674385
transform 1 0 7820 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_81
timestamp 1646674385
transform 1 0 8556 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1513_
timestamp 1646674385
transform 1 0 6900 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1516_
timestamp 1646674385
transform -1 0 8556 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A
timestamp 1646674385
transform -1 0 10396 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A
timestamp 1646674385
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_101
timestamp 1646674385
transform 1 0 10396 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1646674385
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_94
timestamp 1646674385
transform 1 0 9752 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_98
timestamp 1646674385
transform 1 0 10120 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2178_
timestamp 1646674385
transform -1 0 9752 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1646674385
transform 1 0 11040 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_122
timestamp 1646674385
transform 1 0 12328 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1646674385
transform 1 0 11408 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2175_
timestamp 1646674385
transform 1 0 10764 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2176_
timestamp 1646674385
transform 1 0 11500 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1646674385
transform 1 0 13708 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1315_
timestamp 1646674385
transform -1 0 14904 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2194_
timestamp 1646674385
transform -1 0 13708 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_150
timestamp 1646674385
transform 1 0 14904 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1646674385
transform 1 0 16192 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1312_
timestamp 1646674385
transform -1 0 16192 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_37_172
timestamp 1646674385
transform 1 0 16928 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_176
timestamp 1646674385
transform 1 0 17296 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_187
timestamp 1646674385
transform 1 0 18308 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1646674385
transform 1 0 16560 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1322_
timestamp 1646674385
transform -1 0 18308 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2491_
timestamp 1646674385
transform 1 0 16652 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_201
timestamp 1646674385
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1329_
timestamp 1646674385
transform 1 0 18676 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1330_
timestamp 1646674385
transform 1 0 19964 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1646674385
transform 1 0 20884 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1646674385
transform 1 0 21620 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1646674385
transform 1 0 21804 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1646674385
transform 1 0 21712 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _2384_
timestamp 1646674385
transform -1 0 22632 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_37_234
timestamp 1646674385
transform 1 0 22632 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2735_
timestamp 1646674385
transform 1 0 23184 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__A
timestamp 1646674385
transform 1 0 25024 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1646674385
transform 1 0 24656 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1646674385
transform 1 0 25208 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1630_
timestamp 1646674385
transform 1 0 25576 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1646674385
transform 1 0 26496 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1646674385
transform 1 0 26956 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1646674385
transform 1 0 26864 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1635_
timestamp 1646674385
transform -1 0 28244 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_37_295
timestamp 1646674385
transform 1 0 28244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2731_
timestamp 1646674385
transform -1 0 30084 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_37_315
timestamp 1646674385
transform 1 0 30084 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_321
timestamp 1646674385
transform 1 0 30636 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_329
timestamp 1646674385
transform 1 0 31372 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1646674385
transform -1 0 32016 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2534_
timestamp 1646674385
transform 1 0 30728 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_38_14
timestamp 1646674385
transform 1 0 2392 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1646674385
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1646674385
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1478_
timestamp 1646674385
transform -1 0 2392 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2027__A2
timestamp 1646674385
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2029__A2
timestamp 1646674385
transform 1 0 4140 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2099__A2
timestamp 1646674385
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1646674385
transform 1 0 3312 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1646674385
transform 1 0 3772 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1646674385
transform 1 0 4324 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1646674385
transform 1 0 4876 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1646674385
transform 1 0 3680 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__A
timestamp 1646674385
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_54
timestamp 1646674385
transform 1 0 6072 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_60
timestamp 1646674385
transform 1 0 6624 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1514_
timestamp 1646674385
transform -1 0 6072 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1646674385
transform 1 0 8464 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2802_
timestamp 1646674385
transform 1 0 6992 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1646674385
transform 1 0 8924 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1646674385
transform 1 0 9476 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_95
timestamp 1646674385
transform 1 0 9844 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1646674385
transform 1 0 8832 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1401_
timestamp 1646674385
transform 1 0 9936 0 1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _2179_
timestamp 1646674385
transform 1 0 9016 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_38_106
timestamp 1646674385
transform 1 0 10856 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_120
timestamp 1646674385
transform 1 0 12144 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1398_
timestamp 1646674385
transform 1 0 11224 0 1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_38_128
timestamp 1646674385
transform 1 0 12880 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1646674385
transform 1 0 13616 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1646674385
transform 1 0 14076 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1646674385
transform 1 0 13984 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1316_
timestamp 1646674385
transform -1 0 15272 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2196_
timestamp 1646674385
transform 1 0 12972 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_38_154
timestamp 1646674385
transform 1 0 15272 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_158
timestamp 1646674385
transform 1 0 15640 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2902_
timestamp 1646674385
transform 1 0 15732 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_175
timestamp 1646674385
transform 1 0 17204 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_179
timestamp 1646674385
transform 1 0 17572 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1646674385
transform 1 0 17940 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1337_
timestamp 1646674385
transform -1 0 18676 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2376_
timestamp 1646674385
transform -1 0 17940 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1646674385
transform 1 0 18676 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1646674385
transform 1 0 19044 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1646674385
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_208
timestamp 1646674385
transform 1 0 20240 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1646674385
transform 1 0 19136 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1336_
timestamp 1646674385
transform -1 0 20240 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1646674385
transform 1 0 20608 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1926__A
timestamp 1646674385
transform 1 0 22172 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2015__A
timestamp 1646674385
transform -1 0 21344 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_214
timestamp 1646674385
transform 1 0 20792 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_220
timestamp 1646674385
transform 1 0 21344 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_228
timestamp 1646674385
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_231
timestamp 1646674385
transform 1 0 22356 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_237
timestamp 1646674385
transform 1 0 22908 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_241
timestamp 1646674385
transform 1 0 23276 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1646674385
transform 1 0 23920 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2385_
timestamp 1646674385
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2416_
timestamp 1646674385
transform -1 0 23276 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_262
timestamp 1646674385
transform 1 0 25208 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1646674385
transform 1 0 24288 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1632_
timestamp 1646674385
transform -1 0 25208 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1634_
timestamp 1646674385
transform 1 0 25576 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_275
timestamp 1646674385
transform 1 0 26404 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1646674385
transform 1 0 27600 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1637_
timestamp 1646674385
transform -1 0 27600 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1635__A
timestamp 1646674385
transform -1 0 29716 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1646674385
transform 1 0 28796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1646674385
transform 1 0 29348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_311
timestamp 1646674385
transform 1 0 29716 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1646674385
transform 1 0 29440 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1639_
timestamp 1646674385
transform -1 0 28796 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_321
timestamp 1646674385
transform 1 0 30636 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_329
timestamp 1646674385
transform 1 0 31372 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1646674385
transform -1 0 32016 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2533_
timestamp 1646674385
transform 1 0 31004 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _2549_
timestamp 1646674385
transform -1 0 30636 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_19
timestamp 1646674385
transform 1 0 2852 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_17
timestamp 1646674385
transform 1 0 2668 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1646674385
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1646674385
transform 1 0 1748 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1646674385
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1646674385
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1474_
timestamp 1646674385
transform 1 0 1840 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2821_
timestamp 1646674385
transform 1 0 1380 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__o221a_1  _1510_
timestamp 1646674385
transform -1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1441_
timestamp 1646674385
transform -1 0 4140 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1646674385
transform 1 0 3680 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1646674385
transform 1 0 3312 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_21
timestamp 1646674385
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2099__A1
timestamp 1646674385
transform -1 0 3312 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_37
timestamp 1646674385
transform 1 0 4508 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_33
timestamp 1646674385
transform 1 0 4140 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_32
timestamp 1646674385
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_prog_clk
timestamp 1646674385
transform 1 0 4600 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2804_
timestamp 1646674385
transform -1 0 5888 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1646674385
transform 1 0 5888 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1646674385
transform 1 0 6348 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_58
timestamp 1646674385
transform 1 0 6440 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1646674385
transform 1 0 6256 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1517_
timestamp 1646674385
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2801_
timestamp 1646674385
transform 1 0 6532 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_39_75
timestamp 1646674385
transform 1 0 8004 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_83
timestamp 1646674385
transform 1 0 8740 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_71
timestamp 1646674385
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_75
timestamp 1646674385
transform 1 0 8004 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1646674385
transform 1 0 8464 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2184_
timestamp 1646674385
transform 1 0 8096 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2581_
timestamp 1646674385
transform -1 0 10120 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1646674385
transform 1 0 8832 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1646674385
transform 1 0 8924 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1404_
timestamp 1646674385
transform 1 0 10212 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1402_
timestamp 1646674385
transform 1 0 10580 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_98
timestamp 1646674385
transform 1 0 10120 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_102
timestamp 1646674385
transform 1 0 10488 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_98
timestamp 1646674385
transform 1 0 10120 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_94
timestamp 1646674385
transform 1 0 9752 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _2180_
timestamp 1646674385
transform -1 0 9752 0 -1 22304
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1646674385
transform 1 0 11040 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_112
timestamp 1646674385
transform 1 0 11408 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1646674385
transform 1 0 11408 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2853_
timestamp 1646674385
transform 1 0 11500 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2855_
timestamp 1646674385
transform 1 0 11776 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1646674385
transform 1 0 12972 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_136
timestamp 1646674385
transform 1 0 13616 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_144
timestamp 1646674385
transform 1 0 14352 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1646674385
transform 1 0 13248 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1646674385
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1646674385
transform 1 0 13984 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1310_
timestamp 1646674385
transform 1 0 14444 0 1 22304
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2262_
timestamp 1646674385
transform 1 0 13340 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2433_
timestamp 1646674385
transform -1 0 14720 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_148
timestamp 1646674385
transform 1 0 14720 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1646674385
transform 1 0 16008 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1646674385
transform 1 0 15364 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1314_
timestamp 1646674385
transform -1 0 16008 0 -1 22304
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2901_
timestamp 1646674385
transform 1 0 15732 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1646674385
transform 1 0 16652 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_179
timestamp 1646674385
transform 1 0 17572 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_187
timestamp 1646674385
transform 1 0 18308 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1646674385
transform 1 0 17204 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1646674385
transform 1 0 16560 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2434_
timestamp 1646674385
transform 1 0 16744 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _2436_
timestamp 1646674385
transform 1 0 17572 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1646674385
transform 1 0 19228 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1646674385
transform 1 0 18768 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1646674385
transform 1 0 19228 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1646674385
transform 1 0 19136 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1334_
timestamp 1646674385
transform 1 0 18400 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2891_
timestamp 1646674385
transform -1 0 21068 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2892_
timestamp 1646674385
transform 1 0 19596 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1646674385
transform 1 0 21068 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1646674385
transform 1 0 21620 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1646674385
transform 1 0 21804 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_217
timestamp 1646674385
transform 1 0 21068 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_223
timestamp 1646674385
transform 1 0 21620 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1646674385
transform 1 0 21712 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2889_
timestamp 1646674385
transform 1 0 21712 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_prog_clk
timestamp 1646674385
transform 1 0 22172 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1631__A1
timestamp 1646674385
transform 1 0 23736 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1646674385
transform 1 0 24012 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_240
timestamp 1646674385
transform 1 0 23184 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1646674385
transform 1 0 23920 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_262
timestamp 1646674385
transform 1 0 25208 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_270
timestamp 1646674385
transform 1 0 25944 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_269
timestamp 1646674385
transform 1 0 25852 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1646674385
transform 1 0 24288 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1631_
timestamp 1646674385
transform 1 0 24380 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2737_
timestamp 1646674385
transform -1 0 25852 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1646674385
transform 1 0 26496 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_284
timestamp 1646674385
transform 1 0 27232 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_275
timestamp 1646674385
transform 1 0 26404 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_285
timestamp 1646674385
transform 1 0 27324 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1646674385
transform 1 0 26864 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2380_
timestamp 1646674385
transform 1 0 26956 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2402_
timestamp 1646674385
transform 1 0 26036 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2420_
timestamp 1646674385
transform -1 0 27324 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1641_
timestamp 1646674385
transform 1 0 28152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1640_
timestamp 1646674385
transform 1 0 28060 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_40_293
timestamp 1646674385
transform 1 0 28060 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_302
timestamp 1646674385
transform 1 0 28888 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_292
timestamp 1646674385
transform 1 0 27968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2415_
timestamp 1646674385
transform 1 0 29256 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1646674385
transform 1 0 29440 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1646674385
transform 1 0 29348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_303
timestamp 1646674385
transform 1 0 28980 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_309
timestamp 1646674385
transform 1 0 29532 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2730_
timestamp 1646674385
transform -1 0 31004 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1636__A
timestamp 1646674385
transform -1 0 30084 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_315
timestamp 1646674385
transform 1 0 30084 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_322
timestamp 1646674385
transform 1 0 30728 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_329
timestamp 1646674385
transform 1 0 31372 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_325
timestamp 1646674385
transform 1 0 31004 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1646674385
transform -1 0 32016 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1646674385
transform -1 0 32016 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2567_
timestamp 1646674385
transform 1 0 31096 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output36
timestamp 1646674385
transform -1 0 30728 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1646674385
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_7
timestamp 1646674385
transform 1 0 1748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1646674385
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2824_
timestamp 1646674385
transform 1 0 1840 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2098__A2
timestamp 1646674385
transform -1 0 3956 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_24
timestamp 1646674385
transform 1 0 3312 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_28
timestamp 1646674385
transform 1 0 3680 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_31
timestamp 1646674385
transform 1 0 3956 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2805_
timestamp 1646674385
transform 1 0 4324 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1646674385
transform 1 0 5796 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1646674385
transform 1 0 6164 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1646674385
transform 1 0 6256 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1518_
timestamp 1646674385
transform 1 0 6348 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_66
timestamp 1646674385
transform 1 0 7176 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_74
timestamp 1646674385
transform 1 0 7912 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_82
timestamp 1646674385
transform 1 0 8648 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1430_
timestamp 1646674385
transform -1 0 7912 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2182_
timestamp 1646674385
transform 1 0 8280 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_103
timestamp 1646674385
transform 1 0 10580 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _2185_
timestamp 1646674385
transform -1 0 10580 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1646674385
transform 1 0 11316 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_116
timestamp 1646674385
transform 1 0 11776 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_124
timestamp 1646674385
transform 1 0 12512 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1646674385
transform 1 0 11408 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _1964_
timestamp 1646674385
transform 1 0 12604 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2177_
timestamp 1646674385
transform 1 0 11500 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_131
timestamp 1646674385
transform 1 0 13156 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2903_
timestamp 1646674385
transform 1 0 13524 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_151
timestamp 1646674385
transform 1 0 14996 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1646674385
transform 1 0 16192 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1320_
timestamp 1646674385
transform 1 0 15364 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1646674385
transform 1 0 16652 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1646674385
transform 1 0 17204 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1646674385
transform 1 0 16560 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1319_
timestamp 1646674385
transform -1 0 17204 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1646674385
transform 1 0 17572 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_41_199
timestamp 1646674385
transform 1 0 19412 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_207
timestamp 1646674385
transform 1 0 20148 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1335_
timestamp 1646674385
transform 1 0 19780 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1646674385
transform 1 0 21344 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1646674385
transform 1 0 21712 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1339_
timestamp 1646674385
transform 1 0 21804 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1340_
timestamp 1646674385
transform 1 0 20516 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A
timestamp 1646674385
transform -1 0 23184 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_234
timestamp 1646674385
transform 1 0 22632 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_240
timestamp 1646674385
transform 1 0 23184 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2736_
timestamp 1646674385
transform 1 0 23552 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_41_261
timestamp 1646674385
transform 1 0 25116 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2423_
timestamp 1646674385
transform 1 0 25852 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1646674385
transform 1 0 26496 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1646674385
transform 1 0 26956 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1646674385
transform 1 0 26864 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _2419_
timestamp 1646674385
transform 1 0 27324 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2176__A2
timestamp 1646674385
transform 1 0 29624 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_292
timestamp 1646674385
transform 1 0 27968 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_299
timestamp 1646674385
transform 1 0 28612 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_306
timestamp 1646674385
transform 1 0 29256 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_312
timestamp 1646674385
transform 1 0 29808 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2417_
timestamp 1646674385
transform -1 0 28612 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2418_
timestamp 1646674385
transform 1 0 28980 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2176__B2
timestamp 1646674385
transform 1 0 30176 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_318
timestamp 1646674385
transform 1 0 30360 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_329
timestamp 1646674385
transform 1 0 31372 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1646674385
transform -1 0 32016 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2571_
timestamp 1646674385
transform -1 0 31372 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2040__A2
timestamp 1646674385
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_13
timestamp 1646674385
transform 1 0 2300 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1646674385
transform 1 0 2852 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1646674385
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1646674385
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1646674385
transform 1 0 1748 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1646674385
transform 1 0 3588 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1646674385
transform 1 0 3680 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2827_
timestamp 1646674385
transform -1 0 5244 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_45
timestamp 1646674385
transform 1 0 5244 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_53
timestamp 1646674385
transform 1 0 5980 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1511_
timestamp 1646674385
transform 1 0 6072 0 1 23392
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_42_64
timestamp 1646674385
transform 1 0 6992 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1646674385
transform 1 0 8188 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1646674385
transform 1 0 8740 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1520_
timestamp 1646674385
transform 1 0 7360 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__A
timestamp 1646674385
transform -1 0 10212 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1646674385
transform 1 0 9660 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1646674385
transform 1 0 10212 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1646674385
transform 1 0 8832 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2183_
timestamp 1646674385
transform 1 0 8924 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2856_
timestamp 1646674385
transform -1 0 12052 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_119
timestamp 1646674385
transform 1 0 12052 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2273_
timestamp 1646674385
transform 1 0 12420 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A
timestamp 1646674385
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_130
timestamp 1646674385
transform 1 0 13064 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1646674385
transform 1 0 13616 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1646674385
transform 1 0 14076 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1646674385
transform 1 0 13984 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1317_
timestamp 1646674385
transform -1 0 15272 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_42_154
timestamp 1646674385
transform 1 0 15272 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_160
timestamp 1646674385
transform 1 0 15824 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_165
timestamp 1646674385
transform 1 0 16284 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _2435_
timestamp 1646674385
transform 1 0 15916 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_175
timestamp 1646674385
transform 1 0 17204 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2015_
timestamp 1646674385
transform 1 0 16652 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2377_
timestamp 1646674385
transform 1 0 17940 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1646674385
transform 1 0 18768 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1646674385
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_206
timestamp 1646674385
transform 1 0 20056 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1646674385
transform 1 0 19136 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _2378_
timestamp 1646674385
transform -1 0 20056 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_42_214
timestamp 1646674385
transform 1 0 20792 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1646674385
transform 1 0 20424 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2890_
timestamp 1646674385
transform -1 0 23000 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_238
timestamp 1646674385
transform 1 0 23000 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1646674385
transform 1 0 23644 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2392_
timestamp 1646674385
transform -1 0 23644 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1646674385
transform 1 0 24196 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_260
timestamp 1646674385
transform 1 0 25024 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1646674385
transform 1 0 25852 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1646674385
transform 1 0 24288 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _2395_
timestamp 1646674385
transform 1 0 24380 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2400_
timestamp 1646674385
transform 1 0 25392 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_42_278
timestamp 1646674385
transform 1 0 26680 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_287
timestamp 1646674385
transform 1 0 27508 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2386_
timestamp 1646674385
transform 1 0 26220 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2405_
timestamp 1646674385
transform 1 0 27048 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1646674385
transform 1 0 28060 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 1646674385
transform 1 0 28980 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1646674385
transform 1 0 29348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1646674385
transform 1 0 29440 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1642_
timestamp 1646674385
transform 1 0 28152 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2729_
timestamp 1646674385
transform -1 0 31004 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_325
timestamp 1646674385
transform 1 0 31004 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1646674385
transform -1 0 32016 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_17
timestamp 1646674385
transform 1 0 2668 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1646674385
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1646674385
transform 1 0 1748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1646674385
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1471_
timestamp 1646674385
transform 1 0 1840 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_43_23
timestamp 1646674385
transform 1 0 3220 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_34
timestamp 1646674385
transform 1 0 4232 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1462_
timestamp 1646674385
transform -1 0 4232 0 -1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_43_42
timestamp 1646674385
transform 1 0 4968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1646674385
transform 1 0 5888 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1646674385
transform 1 0 6348 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1646674385
transform 1 0 6256 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1515_
timestamp 1646674385
transform -1 0 5888 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2800_
timestamp 1646674385
transform -1 0 8004 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_43_75
timestamp 1646674385
transform 1 0 8004 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_81
timestamp 1646674385
transform 1 0 8556 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2181_
timestamp 1646674385
transform 1 0 8648 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_103
timestamp 1646674385
transform 1 0 10580 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_90
timestamp 1646674385
transform 1 0 9384 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_97
timestamp 1646674385
transform 1 0 10028 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1390_
timestamp 1646674385
transform -1 0 11040 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1878_
timestamp 1646674385
transform -1 0 10028 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1646674385
transform 1 0 11040 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_123
timestamp 1646674385
transform 1 0 12420 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1646674385
transform 1 0 11408 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1396_
timestamp 1646674385
transform 1 0 11500 0 -1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_43_140
timestamp 1646674385
transform 1 0 13984 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _2080_
timestamp 1646674385
transform 1 0 14352 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2274_
timestamp 1646674385
transform 1 0 12788 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__A
timestamp 1646674385
transform 1 0 16008 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1646674385
transform 1 0 14904 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1646674385
transform 1 0 15640 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1646674385
transform 1 0 16192 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1313_
timestamp 1646674385
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1646674385
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1646674385
transform 1 0 16560 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1345_
timestamp 1646674385
transform 1 0 17940 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1348_
timestamp 1646674385
transform -1 0 17572 0 -1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_43_192
timestamp 1646674385
transform 1 0 18768 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_196
timestamp 1646674385
transform 1 0 19136 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_204
timestamp 1646674385
transform 1 0 19872 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _2379_
timestamp 1646674385
transform 1 0 19228 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1896__B1
timestamp 1646674385
transform -1 0 21988 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_210
timestamp 1646674385
transform 1 0 20424 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1646674385
transform 1 0 21344 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_227
timestamp 1646674385
transform 1 0 21988 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1646674385
transform 1 0 21712 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1342_
timestamp 1646674385
transform 1 0 20516 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_240
timestamp 1646674385
transform 1 0 23184 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2393_
timestamp 1646674385
transform 1 0 22356 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _2394_
timestamp 1646674385
transform 1 0 23552 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1855__B
timestamp 1646674385
transform 1 0 25484 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1894__A_N
timestamp 1646674385
transform 1 0 24748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_251
timestamp 1646674385
transform 1 0 24196 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_259
timestamp 1646674385
transform 1 0 24932 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_267
timestamp 1646674385
transform 1 0 25668 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1646674385
transform 1 0 26496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_286
timestamp 1646674385
transform 1 0 27416 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1646674385
transform 1 0 26864 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2397_
timestamp 1646674385
transform 1 0 26956 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2414_
timestamp 1646674385
transform -1 0 26496 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2093__B2
timestamp 1646674385
transform 1 0 29348 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_292
timestamp 1646674385
transform 1 0 27968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_296
timestamp 1646674385
transform 1 0 28336 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_303
timestamp 1646674385
transform 1 0 28980 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_309
timestamp 1646674385
transform 1 0 29532 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2409_
timestamp 1646674385
transform -1 0 28336 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2411_
timestamp 1646674385
transform -1 0 28980 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2116__A
timestamp 1646674385
transform 1 0 30544 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2118__C
timestamp 1646674385
transform 1 0 29900 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_315
timestamp 1646674385
transform 1 0 30084 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_319
timestamp 1646674385
transform 1 0 30452 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_322
timestamp 1646674385
transform 1 0 30728 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_329
timestamp 1646674385
transform 1 0 31372 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1646674385
transform -1 0 32016 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output48
timestamp 1646674385
transform -1 0 31372 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1646674385
transform 1 0 2852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1646674385
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2825_
timestamp 1646674385
transform -1 0 2852 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1646674385
transform 1 0 3588 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_38
timestamp 1646674385
transform 1 0 4600 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1646674385
transform 1 0 3680 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1467_
timestamp 1646674385
transform 1 0 3772 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_58
timestamp 1646674385
transform 1 0 6440 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1509_
timestamp 1646674385
transform 1 0 6808 0 1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2803_
timestamp 1646674385
transform 1 0 4968 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_72
timestamp 1646674385
transform 1 0 7728 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1646674385
transform 1 0 8464 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1519_
timestamp 1646674385
transform -1 0 8464 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A
timestamp 1646674385
transform -1 0 10396 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_101
timestamp 1646674385
transform 1 0 10396 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_88
timestamp 1646674385
transform 1 0 9200 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_95
timestamp 1646674385
transform 1 0 9844 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1646674385
transform 1 0 8832 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1879_
timestamp 1646674385
transform 1 0 8924 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1880_
timestamp 1646674385
transform -1 0 9844 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_114
timestamp 1646674385
transform 1 0 11592 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1397_
timestamp 1646674385
transform 1 0 10764 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2272_
timestamp 1646674385
transform 1 0 12328 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_44_131
timestamp 1646674385
transform 1 0 13156 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1646674385
transform 1 0 13892 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1646674385
transform 1 0 13984 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2904_
timestamp 1646674385
transform 1 0 14076 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1646674385
transform 1 0 15548 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_165
timestamp 1646674385
transform 1 0 16284 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1356_
timestamp 1646674385
transform 1 0 15916 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_171
timestamp 1646674385
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk
timestamp 1646674385
transform -1 0 18768 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1646674385
transform 1 0 18768 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1646674385
transform 1 0 19228 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_207
timestamp 1646674385
transform 1 0 20148 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1646674385
transform 1 0 19136 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1341_
timestamp 1646674385
transform 1 0 19320 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_214
timestamp 1646674385
transform 1 0 20792 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_218
timestamp 1646674385
transform 1 0 21160 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2387_
timestamp 1646674385
transform -1 0 20792 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2887_
timestamp 1646674385
transform -1 0 22724 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1841__B
timestamp 1646674385
transform -1 0 23920 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_235
timestamp 1646674385
transform 1 0 22724 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_242
timestamp 1646674385
transform 1 0 23368 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1646674385
transform 1 0 23920 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2326_
timestamp 1646674385
transform -1 0 23368 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_256
timestamp 1646674385
transform 1 0 24656 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_260
timestamp 1646674385
transform 1 0 25024 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_269
timestamp 1646674385
transform 1 0 25852 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1646674385
transform 1 0 24288 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1857_
timestamp 1646674385
transform 1 0 24380 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2426_
timestamp 1646674385
transform 1 0 25116 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_281
timestamp 1646674385
transform 1 0 26956 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_287
timestamp 1646674385
transform 1 0 27508 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2413_
timestamp 1646674385
transform 1 0 27600 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _2425_
timestamp 1646674385
transform 1 0 26220 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_297
timestamp 1646674385
transform 1 0 28428 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1646674385
transform 1 0 29072 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1646674385
transform 1 0 29440 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2408_
timestamp 1646674385
transform -1 0 29072 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2728_
timestamp 1646674385
transform -1 0 31004 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_44_325
timestamp 1646674385
transform 1 0 31004 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1646674385
transform -1 0 32016 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_13
timestamp 1646674385
transform 1 0 2300 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_7
timestamp 1646674385
transform 1 0 1748 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1646674385
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1464_
timestamp 1646674385
transform 1 0 2392 0 -1 25568
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1646674385
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__A
timestamp 1646674385
transform 1 0 3680 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__B1
timestamp 1646674385
transform -1 0 4784 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1646674385
transform 1 0 3312 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_30
timestamp 1646674385
transform 1 0 3864 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1646674385
transform 1 0 4784 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__B2
timestamp 1646674385
transform -1 0 5336 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2093__A2
timestamp 1646674385
transform 1 0 5704 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_46
timestamp 1646674385
transform 1 0 5336 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1646674385
transform 1 0 5888 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp 1646674385
transform 1 0 6348 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1646674385
transform 1 0 6256 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1427_
timestamp 1646674385
transform 1 0 6624 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_64
timestamp 1646674385
transform 1 0 6992 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_68
timestamp 1646674385
transform 1 0 7360 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1646674385
transform 1 0 8372 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1432_
timestamp 1646674385
transform -1 0 8372 0 -1 25568
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1881_
timestamp 1646674385
transform -1 0 9016 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_103
timestamp 1646674385
transform 1 0 10580 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1646674385
transform 1 0 9016 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_90
timestamp 1646674385
transform 1 0 9384 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_95
timestamp 1646674385
transform 1 0 9844 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1387_
timestamp 1646674385
transform -1 0 11040 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1425_
timestamp 1646674385
transform -1 0 9844 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1646674385
transform 1 0 11040 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_123
timestamp 1646674385
transform 1 0 12420 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1646674385
transform 1 0 11408 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1391_
timestamp 1646674385
transform -1 0 12420 0 -1 25568
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_45_134
timestamp 1646674385
transform 1 0 13432 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2287_
timestamp 1646674385
transform 1 0 12788 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2492_
timestamp 1646674385
transform -1 0 14628 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_147
timestamp 1646674385
transform 1 0 14628 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1646674385
transform 1 0 16192 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2494_
timestamp 1646674385
transform 1 0 14996 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_45_173
timestamp 1646674385
transform 1 0 17020 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_177
timestamp 1646674385
transform 1 0 17388 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1646674385
transform 1 0 16560 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1416_
timestamp 1646674385
transform 1 0 16652 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2885_
timestamp 1646674385
transform 1 0 17480 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_194
timestamp 1646674385
transform 1 0 18952 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2886_
timestamp 1646674385
transform -1 0 20792 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A
timestamp 1646674385
transform -1 0 21344 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_214
timestamp 1646674385
transform 1 0 20792 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1646674385
transform 1 0 21344 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1646674385
transform 1 0 21712 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _2390_
timestamp 1646674385
transform 1 0 21804 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_45_232
timestamp 1646674385
transform 1 0 22448 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_238
timestamp 1646674385
transform 1 0 23000 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2606_
timestamp 1646674385
transform 1 0 23092 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_255
timestamp 1646674385
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_267
timestamp 1646674385
transform 1 0 25668 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _1894_
timestamp 1646674385
transform -1 0 25668 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1646674385
transform 1 0 26496 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_288
timestamp 1646674385
transform 1 0 27600 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1646674385
transform 1 0 26864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1855_
timestamp 1646674385
transform -1 0 26496 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2412_
timestamp 1646674385
transform -1 0 27600 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_302
timestamp 1646674385
transform 1 0 28888 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1638_
timestamp 1646674385
transform 1 0 27968 0 -1 25568
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1646_
timestamp 1646674385
transform 1 0 29256 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_315
timestamp 1646674385
transform 1 0 30084 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_322
timestamp 1646674385
transform 1 0 30728 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_329
timestamp 1646674385
transform 1 0 31372 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1646674385
transform -1 0 32016 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2410_
timestamp 1646674385
transform 1 0 30452 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1646674385
transform -1 0 31372 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__B2
timestamp 1646674385
transform -1 0 1656 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_19
timestamp 1646674385
transform 1 0 2852 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_19
timestamp 1646674385
transform 1 0 2852 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_3
timestamp 1646674385
transform 1 0 1380 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_6
timestamp 1646674385
transform 1 0 1656 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1646674385
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1646674385
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1469_
timestamp 1646674385
transform 1 0 2024 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2826_
timestamp 1646674385
transform -1 0 2852 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1646674385
transform 1 0 3588 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_41
timestamp 1646674385
transform 1 0 4876 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1646674385
transform 1 0 3680 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2828_
timestamp 1646674385
transform -1 0 4876 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2829_
timestamp 1646674385
transform 1 0 3772 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1912_
timestamp 1646674385
transform -1 0 5888 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1646674385
transform 1 0 5888 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_51
timestamp 1646674385
transform 1 0 5796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_45
timestamp 1646674385
transform 1 0 5244 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2038__A2
timestamp 1646674385
transform 1 0 5612 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1440_
timestamp 1646674385
transform -1 0 7636 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1646674385
transform 1 0 6256 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1646674385
transform 1 0 6348 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_58
timestamp 1646674385
transform 1 0 6440 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_55
timestamp 1646674385
transform 1 0 6164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A
timestamp 1646674385
transform -1 0 6440 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2840_
timestamp 1646674385
transform 1 0 6716 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_46_71
timestamp 1646674385
transform 1 0 7636 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_79
timestamp 1646674385
transform 1 0 8372 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1646674385
transform 1 0 8740 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_77
timestamp 1646674385
transform 1 0 8188 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1431_
timestamp 1646674385
transform 1 0 8004 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1433_
timestamp 1646674385
transform 1 0 8556 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A
timestamp 1646674385
transform -1 0 9936 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2080__A
timestamp 1646674385
transform -1 0 10488 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_102
timestamp 1646674385
transform 1 0 10488 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1646674385
transform 1 0 8924 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_102
timestamp 1646674385
transform 1 0 10488 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_90
timestamp 1646674385
transform 1 0 9384 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_96
timestamp 1646674385
transform 1 0 9936 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1646674385
transform 1 0 8832 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2844_
timestamp 1646674385
transform 1 0 9016 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__A
timestamp 1646674385
transform -1 0 11224 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2043__A
timestamp 1646674385
transform -1 0 11040 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_110
timestamp 1646674385
transform 1 0 11224 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1646674385
transform 1 0 11040 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1646674385
transform 1 0 12328 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1646674385
transform 1 0 11408 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1394_
timestamp 1646674385
transform 1 0 11500 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2858_
timestamp 1646674385
transform -1 0 13064 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1646674385
transform -1 0 14260 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A
timestamp 1646674385
transform -1 0 13616 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_130
timestamp 1646674385
transform 1 0 13064 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1646674385
transform 1 0 13616 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_143
timestamp 1646674385
transform 1 0 14260 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_129
timestamp 1646674385
transform 1 0 12972 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1646674385
transform 1 0 13984 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2285_
timestamp 1646674385
transform 1 0 12696 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2288_
timestamp 1646674385
transform 1 0 13340 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_46_154
timestamp 1646674385
transform 1 0 15272 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_146
timestamp 1646674385
transform 1 0 14536 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_156
timestamp 1646674385
transform 1 0 15456 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1646674385
transform 1 0 16192 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2016_
timestamp 1646674385
transform 1 0 14904 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2103_
timestamp 1646674385
transform 1 0 15824 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2493_
timestamp 1646674385
transform 1 0 14628 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1646674385
transform -1 0 17480 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_46_178
timestamp 1646674385
transform 1 0 17480 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_169
timestamp 1646674385
transform 1 0 16652 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_183
timestamp 1646674385
transform 1 0 17940 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1646674385
transform 1 0 16560 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2093_
timestamp 1646674385
transform -1 0 18676 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _2104_
timestamp 1646674385
transform 1 0 16744 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_1  _2389_
timestamp 1646674385
transform 1 0 19228 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2322_
timestamp 1646674385
transform 1 0 18492 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1646674385
transform 1 0 19136 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1646674385
transform 1 0 18860 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1646674385
transform 1 0 19228 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1646674385
transform 1 0 19044 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1646674385
transform 1 0 18676 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2388_
timestamp 1646674385
transform 1 0 20240 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_204
timestamp 1646674385
transform 1 0 19872 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1646674385
transform 1 0 19596 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2888_
timestamp 1646674385
transform -1 0 21160 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__A
timestamp 1646674385
transform -1 0 21712 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_218
timestamp 1646674385
transform 1 0 21160 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1646674385
transform 1 0 21712 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1646674385
transform 1 0 21068 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1646674385
transform 1 0 21620 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1646674385
transform 1 0 21804 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1646674385
transform 1 0 21712 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2327_
timestamp 1646674385
transform 1 0 22172 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _2328_
timestamp 1646674385
transform 1 0 22080 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1841__A
timestamp 1646674385
transform 1 0 23736 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_235
timestamp 1646674385
transform 1 0 22724 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_242
timestamp 1646674385
transform 1 0 23368 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1646674385
transform 1 0 23920 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_238
timestamp 1646674385
transform 1 0 23000 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1646674385
transform 1 0 23828 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1841_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 23368 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2321_
timestamp 1646674385
transform 1 0 23092 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1646674385
transform 1 0 24840 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_251
timestamp 1646674385
transform 1 0 24196 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_265
timestamp 1646674385
transform 1 0 25484 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1646674385
transform 1 0 24288 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _1856_
timestamp 1646674385
transform -1 0 24840 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1896_
timestamp 1646674385
transform -1 0 25484 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _2427_
timestamp 1646674385
transform 1 0 25852 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2594_
timestamp 1646674385
transform -1 0 26036 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2424_
timestamp 1646674385
transform -1 0 27232 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1646674385
transform 1 0 26864 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1646674385
transform 1 0 26772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1646674385
transform 1 0 26220 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1646674385
transform 1 0 26036 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2407_
timestamp 1646674385
transform 1 0 27692 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2406_
timestamp 1646674385
transform 1 0 27692 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2391_
timestamp 1646674385
transform 1 0 26956 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_288
timestamp 1646674385
transform 1 0 27600 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_284
timestamp 1646674385
transform 1 0 27232 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_288
timestamp 1646674385
transform 1 0 27600 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_284
timestamp 1646674385
transform 1 0 27232 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2404_
timestamp 1646674385
transform -1 0 28980 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_298
timestamp 1646674385
transform 1 0 28520 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_296
timestamp 1646674385
transform 1 0 28336 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1648_
timestamp 1646674385
transform 1 0 29440 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1646674385
transform 1 0 29440 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_304
timestamp 1646674385
transform 1 0 29072 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1646674385
transform 1 0 29532 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1646674385
transform 1 0 29348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1646674385
transform 1 0 28980 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1652__A
timestamp 1646674385
transform 1 0 28888 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_329
timestamp 1646674385
transform 1 0 31372 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_317
timestamp 1646674385
transform 1 0 30268 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_321
timestamp 1646674385
transform 1 0 30636 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_329
timestamp 1646674385
transform 1 0 31372 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1646674385
transform -1 0 32016 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1646674385
transform -1 0 32016 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _2116_
timestamp 1646674385
transform 1 0 30728 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2727_
timestamp 1646674385
transform -1 0 31372 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2035__B
timestamp 1646674385
transform 1 0 1748 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_17
timestamp 1646674385
transform 1 0 2668 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1646674385
transform 1 0 1380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_9
timestamp 1646674385
transform 1 0 1932 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1646674385
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1468_
timestamp 1646674385
transform 1 0 2300 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__B2
timestamp 1646674385
transform 1 0 3128 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_21
timestamp 1646674385
transform 1 0 3036 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1646674385
transform 1 0 3312 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_38
timestamp 1646674385
transform 1 0 4600 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1646674385
transform 1 0 3680 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1465_
timestamp 1646674385
transform 1 0 3772 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_46
timestamp 1646674385
transform 1 0 5336 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_50
timestamp 1646674385
transform 1 0 5704 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1461_
timestamp 1646674385
transform -1 0 5336 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_prog_clk
timestamp 1646674385
transform -1 0 7636 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__B2
timestamp 1646674385
transform 1 0 8280 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_71
timestamp 1646674385
transform 1 0 7636 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_77
timestamp 1646674385
transform 1 0 8188 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1646674385
transform 1 0 8464 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_101
timestamp 1646674385
transform 1 0 10396 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1646674385
transform 1 0 8832 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2842_
timestamp 1646674385
transform 1 0 8924 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_48_109
timestamp 1646674385
transform 1 0 11132 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_119
timestamp 1646674385
transform 1 0 12052 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1395_
timestamp 1646674385
transform 1 0 11224 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1646674385
transform 1 0 13616 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1646674385
transform 1 0 14076 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1646674385
transform 1 0 13984 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1309_
timestamp 1646674385
transform -1 0 14812 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2286_
timestamp 1646674385
transform 1 0 12788 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_149
timestamp 1646674385
transform 1 0 14812 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_153
timestamp 1646674385
transform 1 0 15180 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2883_
timestamp 1646674385
transform -1 0 16744 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_170
timestamp 1646674385
transform 1 0 16744 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_174
timestamp 1646674385
transform 1 0 17112 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_184
timestamp 1646674385
transform 1 0 18032 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1349_
timestamp 1646674385
transform 1 0 17204 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1646674385
transform 1 0 18676 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1646674385
transform 1 0 19044 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_204
timestamp 1646674385
transform 1 0 19872 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_208
timestamp 1646674385
transform 1 0 20240 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1646674385
transform 1 0 19136 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2092_
timestamp 1646674385
transform -1 0 18676 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2118_
timestamp 1646674385
transform 1 0 19228 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_48_216
timestamp 1646674385
transform 1 0 20976 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_226
timestamp 1646674385
transform 1 0 21896 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1417_
timestamp 1646674385
transform 1 0 21344 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2324_
timestamp 1646674385
transform 1 0 20332 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_48_230
timestamp 1646674385
transform 1 0 22264 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1646674385
transform 1 0 23552 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2329_
timestamp 1646674385
transform 1 0 22356 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_260
timestamp 1646674385
transform 1 0 25024 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_270
timestamp 1646674385
transform 1 0 25944 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1646674385
transform 1 0 24288 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _1308_
timestamp 1646674385
transform 1 0 25392 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1895_
timestamp 1646674385
transform -1 0 25024 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1643__A
timestamp 1646674385
transform 1 0 27600 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_277
timestamp 1646674385
transform 1 0 26588 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1646674385
transform 1 0 27232 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_290
timestamp 1646674385
transform 1 0 27784 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2396_
timestamp 1646674385
transform -1 0 26588 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2398_
timestamp 1646674385
transform 1 0 26956 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_297
timestamp 1646674385
transform 1 0 28428 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1646674385
transform 1 0 29072 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_309
timestamp 1646674385
transform 1 0 29532 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1646674385
transform 1 0 29440 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2399_
timestamp 1646674385
transform -1 0 29072 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2401_
timestamp 1646674385
transform -1 0 28428 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2726_
timestamp 1646674385
transform -1 0 31280 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_328
timestamp 1646674385
transform 1 0 31280 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_332
timestamp 1646674385
transform 1 0 31648 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1646674385
transform -1 0 32016 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__B2
timestamp 1646674385
transform 1 0 2760 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_14
timestamp 1646674385
transform 1 0 2392 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_20
timestamp 1646674385
transform 1 0 2944 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_3
timestamp 1646674385
transform 1 0 1380 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1646674385
transform 1 0 1748 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1646674385
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1931_
timestamp 1646674385
transform -1 0 2392 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2034_
timestamp 1646674385
transform 1 0 1472 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_33
timestamp 1646674385
transform 1 0 4140 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1466_
timestamp 1646674385
transform 1 0 3312 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1646674385
transform -1 0 5152 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_44
timestamp 1646674385
transform 1 0 5152 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1646674385
transform 1 0 5888 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_60
timestamp 1646674385
transform 1 0 6624 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1646674385
transform 1 0 6256 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1911_
timestamp 1646674385
transform -1 0 6624 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2099_
timestamp 1646674385
transform -1 0 5888 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_66
timestamp 1646674385
transform 1 0 7176 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_76
timestamp 1646674385
transform 1 0 8096 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1434_
timestamp 1646674385
transform 1 0 7268 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2843_
timestamp 1646674385
transform 1 0 8464 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__A1
timestamp 1646674385
transform -1 0 10488 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_102
timestamp 1646674385
transform 1 0 10488 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_96
timestamp 1646674385
transform 1 0 9936 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__B2
timestamp 1646674385
transform 1 0 10856 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1646674385
transform 1 0 11040 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1646674385
transform 1 0 11500 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1646674385
transform 1 0 11408 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2857_
timestamp 1646674385
transform 1 0 11868 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_49_133
timestamp 1646674385
transform 1 0 13340 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_141
timestamp 1646674385
transform 1 0 14076 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _2042_
timestamp 1646674385
transform 1 0 14168 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_49_149
timestamp 1646674385
transform 1 0 14812 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_157
timestamp 1646674385
transform 1 0 15548 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1646674385
transform 1 0 16192 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _2043_
timestamp 1646674385
transform 1 0 15640 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1646674385
transform 1 0 17480 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1646674385
transform 1 0 16560 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1351_
timestamp 1646674385
transform -1 0 17480 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1352_
timestamp 1646674385
transform 1 0 17848 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_191
timestamp 1646674385
transform 1 0 18676 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_204
timestamp 1646674385
transform 1 0 19872 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2117_
timestamp 1646674385
transform 1 0 19044 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1646674385
transform 1 0 21252 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1646674385
transform 1 0 21620 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1646674385
transform 1 0 21804 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_229
timestamp 1646674385
transform 1 0 22172 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1646674385
transform 1 0 21712 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2323_
timestamp 1646674385
transform 1 0 20424 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_234
timestamp 1646674385
transform 1 0 22632 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_244
timestamp 1646674385
transform 1 0 23552 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1295_
timestamp 1646674385
transform -1 0 24472 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1298_
timestamp 1646674385
transform -1 0 23552 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1617_
timestamp 1646674385
transform 1 0 22264 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_254
timestamp 1646674385
transform 1 0 24472 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_262
timestamp 1646674385
transform 1 0 25208 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1655_
timestamp 1646674385
transform -1 0 26220 0 -1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1646674385
transform -1 0 27140 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1646674385
transform 1 0 26220 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1646674385
transform 1 0 26772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_283
timestamp 1646674385
transform 1 0 27140 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_291
timestamp 1646674385
transform 1 0 27876 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1646674385
transform 1 0 26864 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1647_
timestamp 1646674385
transform 1 0 27508 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_305
timestamp 1646674385
transform 1 0 29164 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1643_
timestamp 1646674385
transform -1 0 29164 0 -1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1649_
timestamp 1646674385
transform 1 0 29532 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_49_318
timestamp 1646674385
transform 1 0 30360 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_329
timestamp 1646674385
transform 1 0 31372 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1646674385
transform -1 0 32016 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2572_
timestamp 1646674385
transform -1 0 31372 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_9
timestamp 1646674385
transform 1 0 1932 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1646674385
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _2036_
timestamp 1646674385
transform 1 0 2300 0 1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1646674385
transform 1 0 1380 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1646674385
transform 1 0 3220 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1646674385
transform 1 0 3588 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_32
timestamp 1646674385
transform 1 0 4048 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_40
timestamp 1646674385
transform 1 0 4784 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1646674385
transform 1 0 3680 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1914_
timestamp 1646674385
transform 1 0 4876 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2033_
timestamp 1646674385
transform 1 0 3772 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_44
timestamp 1646674385
transform 1 0 5152 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_56
timestamp 1646674385
transform 1 0 6256 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2098_
timestamp 1646674385
transform -1 0 6256 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__B2
timestamp 1646674385
transform 1 0 8280 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_64
timestamp 1646674385
transform 1 0 6992 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_74
timestamp 1646674385
transform 1 0 7912 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1646674385
transform 1 0 8464 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1437_
timestamp 1646674385
transform -1 0 7912 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1646674385
transform 1 0 8924 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 1646674385
transform 1 0 9292 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1646674385
transform 1 0 8832 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2860_
timestamp 1646674385
transform 1 0 9384 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_106
timestamp 1646674385
transform 1 0 10856 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_prog_clk
timestamp 1646674385
transform 1 0 11224 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2032__B2
timestamp 1646674385
transform 1 0 13432 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_130
timestamp 1646674385
transform 1 0 13064 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1646674385
transform 1 0 13616 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1646674385
transform 1 0 13984 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2032_
timestamp 1646674385
transform 1 0 14076 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_150
timestamp 1646674385
transform 1 0 14904 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_154
timestamp 1646674385
transform 1 0 15272 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_165
timestamp 1646674385
transform 1 0 16284 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1343_
timestamp 1646674385
transform -1 0 16284 0 1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_50_183
timestamp 1646674385
transform 1 0 17940 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1344_
timestamp 1646674385
transform 1 0 17020 0 1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1646674385
transform 1 0 18768 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1646674385
transform 1 0 19228 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1646674385
transform 1 0 19136 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2112_
timestamp 1646674385
transform 1 0 18492 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2119_
timestamp 1646674385
transform 1 0 19412 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_50_212
timestamp 1646674385
transform 1 0 20608 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2325_
timestamp 1646674385
transform 1 0 21160 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_231
timestamp 1646674385
transform 1 0 22356 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_235
timestamp 1646674385
transform 1 0 22724 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_240
timestamp 1646674385
transform 1 0 23184 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1646674385
transform 1 0 23920 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1288_
timestamp 1646674385
transform 1 0 23552 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1621_
timestamp 1646674385
transform 1 0 22816 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1646674385
transform 1 0 24380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_257
timestamp 1646674385
transform 1 0 24748 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1646674385
transform 1 0 24288 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2719_
timestamp 1646674385
transform 1 0 24840 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A
timestamp 1646674385
transform 1 0 26680 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_274
timestamp 1646674385
transform 1 0 26312 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_280
timestamp 1646674385
transform 1 0 26864 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1652_
timestamp 1646674385
transform 1 0 27232 0 1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_50_294
timestamp 1646674385
transform 1 0 28152 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1646674385
transform 1 0 28796 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1646674385
transform 1 0 29348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1646674385
transform 1 0 29440 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1651_
timestamp 1646674385
transform 1 0 29532 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2403_
timestamp 1646674385
transform 1 0 28520 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_318
timestamp 1646674385
transform 1 0 30360 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_329
timestamp 1646674385
transform 1 0 31372 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1646674385
transform -1 0 32016 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output49
timestamp 1646674385
transform -1 0 31372 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_10
timestamp 1646674385
transform 1 0 2024 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_3
timestamp 1646674385
transform 1 0 1380 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1646674385
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2040_
timestamp 1646674385
transform -1 0 2024 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _2041_
timestamp 1646674385
transform -1 0 3956 0 -1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_51_31
timestamp 1646674385
transform 1 0 3956 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_38
timestamp 1646674385
transform 1 0 4600 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1933_
timestamp 1646674385
transform 1 0 4324 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_46
timestamp 1646674385
transform 1 0 5336 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1646674385
transform 1 0 5796 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1646674385
transform 1 0 6164 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1646674385
transform 1 0 6256 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2100_
timestamp 1646674385
transform 1 0 6348 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2101_
timestamp 1646674385
transform 1 0 5428 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_65
timestamp 1646674385
transform 1 0 7084 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_71
timestamp 1646674385
transform 1 0 7636 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_82
timestamp 1646674385
transform 1 0 8648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1429_
timestamp 1646674385
transform 1 0 7728 0 -1 28832
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_51_95
timestamp 1646674385
transform 1 0 9844 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1392_
timestamp 1646674385
transform -1 0 11040 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1435_
timestamp 1646674385
transform -1 0 9844 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1646674385
transform 1 0 11040 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_122
timestamp 1646674385
transform 1 0 12328 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1646674385
transform 1 0 11408 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2252_
timestamp 1646674385
transform -1 0 12328 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_51_128
timestamp 1646674385
transform 1 0 12880 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_145
timestamp 1646674385
transform 1 0 14444 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2865_
timestamp 1646674385
transform 1 0 12972 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_156
timestamp 1646674385
transform 1 0 15456 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_163
timestamp 1646674385
transform 1 0 16100 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2019_
timestamp 1646674385
transform 1 0 15824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _2044_
timestamp 1646674385
transform 1 0 14812 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1646674385
transform 1 0 16468 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_178
timestamp 1646674385
transform 1 0 17480 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1646674385
transform 1 0 16560 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1350_
timestamp 1646674385
transform -1 0 17480 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2881_
timestamp 1646674385
transform 1 0 17848 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_51_198
timestamp 1646674385
transform 1 0 19320 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_204
timestamp 1646674385
transform 1 0 19872 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1369_
timestamp 1646674385
transform -1 0 20792 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1895__B
timestamp 1646674385
transform -1 0 21344 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_214
timestamp 1646674385
transform 1 0 20792 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1646674385
transform 1 0 21344 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1646674385
transform 1 0 21804 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1646674385
transform 1 0 21712 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2874_
timestamp 1646674385
transform -1 0 23460 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_243
timestamp 1646674385
transform 1 0 23460 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_250
timestamp 1646674385
transform 1 0 24104 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1646674385
transform -1 0 24104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_263
timestamp 1646674385
transform 1 0 25300 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1658_
timestamp 1646674385
transform 1 0 25668 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1659_
timestamp 1646674385
transform -1 0 25300 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1646674385
transform 1 0 26496 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1646674385
transform 1 0 26956 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_285
timestamp 1646674385
transform 1 0 27324 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1646674385
transform 1 0 26864 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1654_
timestamp 1646674385
transform 1 0 27416 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_295
timestamp 1646674385
transform 1 0 28244 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_308
timestamp 1646674385
transform 1 0 29440 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1650_
timestamp 1646674385
transform 1 0 28612 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2725_
timestamp 1646674385
transform -1 0 31280 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_328
timestamp 1646674385
transform 1 0 31280 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_332
timestamp 1646674385
transform 1 0 31648 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1646674385
transform -1 0 32016 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2037_
timestamp 1646674385
transform 1 0 1840 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2035_
timestamp 1646674385
transform 1 0 1564 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1646674385
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1646674385
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_7
timestamp 1646674385
transform 1 0 1748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1646674385
transform 1 0 1380 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1646674385
transform 1 0 1380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _2599_
timestamp 1646674385
transform -1 0 3220 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_16
timestamp 1646674385
transform 1 0 2576 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_10
timestamp 1646674385
transform 1 0 2024 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2038_
timestamp 1646674385
transform -1 0 3312 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1984_
timestamp 1646674385
transform 1 0 3772 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1928_
timestamp 1646674385
transform 1 0 3772 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1646674385
transform 1 0 3680 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_28
timestamp 1646674385
transform 1 0 3680 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_24
timestamp 1646674385
transform 1 0 3312 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1646674385
transform 1 0 3588 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 1646674385
transform 1 0 3220 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1929_
timestamp 1646674385
transform 1 0 4416 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_37
timestamp 1646674385
transform 1 0 4508 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_32
timestamp 1646674385
transform 1 0 4048 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_39
timestamp 1646674385
transform 1 0 4692 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1985__A2
timestamp 1646674385
transform 1 0 4876 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_46
timestamp 1646674385
transform 1 0 5336 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_60
timestamp 1646674385
transform 1 0 6624 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_43
timestamp 1646674385
transform 1 0 5060 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1646674385
transform 1 0 5888 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1646674385
transform 1 0 6256 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1934_
timestamp 1646674385
transform 1 0 5060 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _2097_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 5428 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _2102_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 5888 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 1646674385
transform -1 0 7176 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1646674385
transform 1 0 8464 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_66
timestamp 1646674385
transform 1 0 7176 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_79
timestamp 1646674385
transform 1 0 8372 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1525_
timestamp 1646674385
transform 1 0 7544 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2094_
timestamp 1646674385
transform 1 0 8740 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2841_
timestamp 1646674385
transform -1 0 8464 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__B1
timestamp 1646674385
transform -1 0 10028 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__B2
timestamp 1646674385
transform -1 0 9108 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_101
timestamp 1646674385
transform 1 0 10396 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_87
timestamp 1646674385
transform 1 0 9108 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 1646674385
transform 1 0 10028 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_86
timestamp 1646674385
transform 1 0 9016 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1646674385
transform 1 0 8832 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1393_
timestamp 1646674385
transform -1 0 11316 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2859_
timestamp 1646674385
transform 1 0 9384 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_2  _2254_
timestamp 1646674385
transform 1 0 11500 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1646674385
transform 1 0 11408 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_106
timestamp 1646674385
transform 1 0 10856 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_111
timestamp 1646674385
transform 1 0 11316 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _2253_
timestamp 1646674385
transform 1 0 11684 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_120
timestamp 1646674385
transform 1 0 12144 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_123
timestamp 1646674385
transform 1 0 12420 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_119
timestamp 1646674385
transform 1 0 12052 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1384_
timestamp 1646674385
transform -1 0 13340 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2042__C
timestamp 1646674385
transform 1 0 12512 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1646674385
transform 1 0 13340 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1646674385
transform 1 0 13892 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1646674385
transform 1 0 14076 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_126
timestamp 1646674385
transform 1 0 12696 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_139
timestamp 1646674385
transform 1 0 13892 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_145
timestamp 1646674385
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1646674385
transform 1 0 13984 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1379_
timestamp 1646674385
transform 1 0 14260 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1382_
timestamp 1646674385
transform 1 0 13064 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__A
timestamp 1646674385
transform 1 0 16284 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2016__A
timestamp 1646674385
transform 1 0 15456 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_152
timestamp 1646674385
transform 1 0 15088 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_158
timestamp 1646674385
transform 1 0 15640 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_164
timestamp 1646674385
transform 1 0 16192 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_156
timestamp 1646674385
transform 1 0 15456 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1646674385
transform 1 0 16192 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1370_
timestamp 1646674385
transform -1 0 16192 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1373_
timestamp 1646674385
transform 1 0 14536 0 -1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_52_167
timestamp 1646674385
transform 1 0 16468 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_173
timestamp 1646674385
transform 1 0 17020 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_184
timestamp 1646674385
transform 1 0 18032 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_185
timestamp 1646674385
transform 1 0 18124 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1646674385
transform 1 0 16560 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1347_
timestamp 1646674385
transform -1 0 18032 0 1 28832
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2884_
timestamp 1646674385
transform 1 0 16652 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1646674385
transform 1 0 19228 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1646674385
transform 1 0 18768 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_199
timestamp 1646674385
transform 1 0 19412 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_203
timestamp 1646674385
transform 1 0 19780 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1646674385
transform 1 0 19136 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1346_
timestamp 1646674385
transform 1 0 18860 0 -1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1353_
timestamp 1646674385
transform -1 0 18768 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1646674385
transform 1 0 20148 0 -1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2872_
timestamp 1646674385
transform -1 0 21252 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_52_219
timestamp 1646674385
transform 1 0 21252 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_227
timestamp 1646674385
transform 1 0 21988 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1646674385
transform 1 0 21068 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1646674385
transform 1 0 21620 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1646674385
transform 1 0 21712 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1367_
timestamp 1646674385
transform 1 0 21804 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2871_
timestamp 1646674385
transform -1 0 23552 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1617__A
timestamp 1646674385
transform -1 0 23184 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1646674385
transform 1 0 23552 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_234
timestamp 1646674385
transform 1 0 22632 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_240
timestamp 1646674385
transform 1 0 23184 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_prog_clk
timestamp 1646674385
transform 1 0 23736 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_52_269
timestamp 1646674385
transform 1 0 25852 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_266
timestamp 1646674385
transform 1 0 25576 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1646674385
transform 1 0 24288 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2421_
timestamp 1646674385
transform -1 0 26220 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2718_
timestamp 1646674385
transform 1 0 24380 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_52_289
timestamp 1646674385
transform 1 0 27692 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1646674385
transform 1 0 26220 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1646674385
transform 1 0 26772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1646674385
transform 1 0 26956 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_285
timestamp 1646674385
transform 1 0 27324 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1646674385
transform 1 0 26864 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2720_
timestamp 1646674385
transform 1 0 26220 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2722_
timestamp 1646674385
transform -1 0 28888 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_52_293
timestamp 1646674385
transform 1 0 28060 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1646674385
transform 1 0 29072 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_302
timestamp 1646674385
transform 1 0 28888 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1646674385
transform 1 0 29440 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1645_
timestamp 1646674385
transform 1 0 28152 0 1 28832
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2723_
timestamp 1646674385
transform -1 0 30728 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2724_
timestamp 1646674385
transform -1 0 31004 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_52_325
timestamp 1646674385
transform 1 0 31004 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_322
timestamp 1646674385
transform 1 0 30728 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_329
timestamp 1646674385
transform 1 0 31372 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1646674385
transform -1 0 32016 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1646674385
transform -1 0 32016 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1646674385
transform -1 0 31372 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_14
timestamp 1646674385
transform 1 0 2392 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_20
timestamp 1646674385
transform 1 0 2944 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1646674385
transform 1 0 1380 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1646674385
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2039_
timestamp 1646674385
transform 1 0 1656 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1981__A2
timestamp 1646674385
transform 1 0 3772 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1646674385
transform 1 0 3312 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_31
timestamp 1646674385
transform 1 0 3956 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1646674385
transform 1 0 3680 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1927_
timestamp 1646674385
transform -1 0 3312 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2598_
timestamp 1646674385
transform -1 0 5152 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2036__A2
timestamp 1646674385
transform 1 0 5520 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_44
timestamp 1646674385
transform 1 0 5152 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_50
timestamp 1646674385
transform 1 0 5704 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_59
timestamp 1646674385
transform 1 0 6532 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2096_
timestamp 1646674385
transform -1 0 6532 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_54_76
timestamp 1646674385
transform 1 0 8096 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1524_
timestamp 1646674385
transform 1 0 7268 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_54_101
timestamp 1646674385
transform 1 0 10396 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1646674385
transform 1 0 8832 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2797_
timestamp 1646674385
transform -1 0 10396 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2037__A2
timestamp 1646674385
transform -1 0 10948 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_107
timestamp 1646674385
transform 1 0 10948 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_114
timestamp 1646674385
transform 1 0 11592 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2251_
timestamp 1646674385
transform 1 0 11316 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2863_
timestamp 1646674385
transform 1 0 12144 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1646674385
transform 1 0 13616 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_141
timestamp 1646674385
transform 1 0 14076 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1646674385
transform 1 0 13984 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2866_
timestamp 1646674385
transform -1 0 15640 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_158
timestamp 1646674385
transform 1 0 15640 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1378_
timestamp 1646674385
transform 1 0 16008 0 1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_54_172
timestamp 1646674385
transform 1 0 16928 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2882_
timestamp 1646674385
transform 1 0 17296 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1646674385
transform 1 0 18768 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_197
timestamp 1646674385
transform 1 0 19228 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_201
timestamp 1646674385
transform 1 0 19596 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1646674385
transform 1 0 19136 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1364_
timestamp 1646674385
transform 1 0 19688 0 1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_54_212
timestamp 1646674385
transform 1 0 20608 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_226
timestamp 1646674385
transform 1 0 21896 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1365_
timestamp 1646674385
transform 1 0 20976 0 1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1621__A
timestamp 1646674385
transform -1 0 23644 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_239
timestamp 1646674385
transform 1 0 23092 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1646674385
transform 1 0 23644 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1371_
timestamp 1646674385
transform 1 0 22264 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1646674385
transform 1 0 24196 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_253
timestamp 1646674385
transform 1 0 24380 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_260
timestamp 1646674385
transform 1 0 25024 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1646674385
transform 1 0 24288 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1644_
timestamp 1646674385
transform 1 0 24656 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1653_
timestamp 1646674385
transform 1 0 25392 0 1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_54_274
timestamp 1646674385
transform 1 0 26312 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2721_
timestamp 1646674385
transform 1 0 26680 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_294
timestamp 1646674385
transform 1 0 28152 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1646674385
transform 1 0 28796 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1646674385
transform 1 0 29348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1646674385
transform 1 0 29440 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2422_
timestamp 1646674385
transform 1 0 28520 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_prog_clk
timestamp 1646674385
transform 1 0 29532 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_54_329
timestamp 1646674385
transform 1 0 31372 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1646674385
transform -1 0 32016 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_11
timestamp 1646674385
transform 1 0 2116 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_18
timestamp 1646674385
transform 1 0 2760 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1646674385
transform 1 0 1380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1646674385
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1920_
timestamp 1646674385
transform -1 0 2760 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1646674385
transform 1 0 1748 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_30
timestamp 1646674385
transform 1 0 3864 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _1981_
timestamp 1646674385
transform 1 0 4232 0 -1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1982_
timestamp 1646674385
transform -1 0 3864 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_44
timestamp 1646674385
transform 1 0 5152 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1646674385
transform 1 0 5796 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1646674385
transform 1 0 6164 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1646674385
transform 1 0 6348 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1646674385
transform 1 0 6256 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1436_
timestamp 1646674385
transform 1 0 6716 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1930_
timestamp 1646674385
transform 1 0 5520 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_65
timestamp 1646674385
transform 1 0 7084 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2798_
timestamp 1646674385
transform 1 0 7452 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__C1
timestamp 1646674385
transform 1 0 9292 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2001__A2
timestamp 1646674385
transform 1 0 9844 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_85
timestamp 1646674385
transform 1 0 8924 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_91
timestamp 1646674385
transform 1 0 9476 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_97
timestamp 1646674385
transform 1 0 10028 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2079__C
timestamp 1646674385
transform 1 0 10856 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_105
timestamp 1646674385
transform 1 0 10764 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1646674385
transform 1 0 11040 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1646674385
transform 1 0 11500 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1646674385
transform 1 0 11408 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1646674385
transform -1 0 12788 0 -1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_55_127
timestamp 1646674385
transform 1 0 12788 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_133
timestamp 1646674385
transform 1 0 13340 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_144
timestamp 1646674385
transform 1 0 14352 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1380_
timestamp 1646674385
transform -1 0 14352 0 -1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1646674385
transform 1 0 16192 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2869_
timestamp 1646674385
transform 1 0 14720 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1646674385
transform 1 0 16652 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_182
timestamp 1646674385
transform 1 0 17848 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1646674385
transform 1 0 16560 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1354_
timestamp 1646674385
transform 1 0 17020 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_prog_clk
timestamp 1646674385
transform 1 0 18216 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_55_206
timestamp 1646674385
transform 1 0 20056 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1646674385
transform 1 0 21344 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1646674385
transform 1 0 21712 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1357_
timestamp 1646674385
transform 1 0 20424 0 -1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1366_
timestamp 1646674385
transform 1 0 21804 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_234
timestamp 1646674385
transform 1 0 22632 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_245
timestamp 1646674385
transform 1 0 23644 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1897_
timestamp 1646674385
transform -1 0 24288 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2333_
timestamp 1646674385
transform 1 0 23000 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1644__A
timestamp 1646674385
transform -1 0 26128 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_252
timestamp 1646674385
transform 1 0 24288 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_266
timestamp 1646674385
transform 1 0 25576 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1662_
timestamp 1646674385
transform -1 0 25576 0 -1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1646674385
transform 1 0 26128 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_281
timestamp 1646674385
transform 1 0 26956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_291
timestamp 1646674385
transform 1 0 27876 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1646674385
transform 1 0 26864 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1656_
timestamp 1646674385
transform 1 0 27048 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2117__A2
timestamp 1646674385
transform -1 0 28428 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2117__B2
timestamp 1646674385
transform 1 0 28796 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2252__B2
timestamp 1646674385
transform 1 0 29348 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_297
timestamp 1646674385
transform 1 0 28428 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_303
timestamp 1646674385
transform 1 0 28980 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_309
timestamp 1646674385
transform 1 0 29532 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2254__B1
timestamp 1646674385
transform -1 0 30084 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2272__B2
timestamp 1646674385
transform 1 0 30452 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2274__B1
timestamp 1646674385
transform -1 0 31188 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_315
timestamp 1646674385
transform 1 0 30084 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_321
timestamp 1646674385
transform 1 0 30636 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_327
timestamp 1646674385
transform 1 0 31188 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1646674385
transform -1 0 32016 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_11
timestamp 1646674385
transform 1 0 2116 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_19
timestamp 1646674385
transform 1 0 2852 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1646674385
transform 1 0 1380 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1646674385
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1985_
timestamp 1646674385
transform 1 0 2944 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1646674385
transform 1 0 1748 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1949__A2
timestamp 1646674385
transform 1 0 3772 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1646674385
transform 1 0 3312 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_31
timestamp 1646674385
transform 1 0 3956 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1646674385
transform 1 0 3680 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_4  _1986_
timestamp 1646674385
transform -1 0 5888 0 1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_56_52
timestamp 1646674385
transform 1 0 5888 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_59
timestamp 1646674385
transform 1 0 6532 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2095_
timestamp 1646674385
transform -1 0 6532 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__C1
timestamp 1646674385
transform 1 0 8188 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1983__A2
timestamp 1646674385
transform 1 0 6900 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_65
timestamp 1646674385
transform 1 0 7084 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_69
timestamp 1646674385
transform 1 0 7452 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_73
timestamp 1646674385
transform 1 0 7820 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_79
timestamp 1646674385
transform 1 0 8372 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1646674385
transform 1 0 8740 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1937_
timestamp 1646674385
transform 1 0 7544 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1998__A2
timestamp 1646674385
transform 1 0 8924 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_87
timestamp 1646674385
transform 1 0 9108 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1646674385
transform 1 0 8832 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2862_
timestamp 1646674385
transform 1 0 9476 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2004__B2
timestamp 1646674385
transform 1 0 12512 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_107
timestamp 1646674385
transform 1 0 10948 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_120
timestamp 1646674385
transform 1 0 12144 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1385_
timestamp 1646674385
transform -1 0 12144 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1963__C
timestamp 1646674385
transform 1 0 14260 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2014__C
timestamp 1646674385
transform 1 0 13064 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_126
timestamp 1646674385
transform 1 0 12696 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_132
timestamp 1646674385
transform 1 0 13248 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1646674385
transform 1 0 14076 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_145
timestamp 1646674385
transform 1 0 14444 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1646674385
transform 1 0 13984 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_159
timestamp 1646674385
transform 1 0 15732 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1372_
timestamp 1646674385
transform 1 0 14812 0 1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_56_167
timestamp 1646674385
transform 1 0 16468 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_175
timestamp 1646674385
transform 1 0 17204 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2079_
timestamp 1646674385
transform 1 0 16560 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2081_
timestamp 1646674385
transform 1 0 17572 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1646674385
transform 1 0 18768 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1646674385
transform 1 0 19228 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_203
timestamp 1646674385
transform 1 0 19780 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1646674385
transform 1 0 19136 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2330_
timestamp 1646674385
transform -1 0 19780 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2876_
timestamp 1646674385
transform 1 0 20148 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1646674385
transform 1 0 21620 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2873_
timestamp 1646674385
transform 1 0 21988 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1646674385
transform 1 0 23460 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1663__B1
timestamp 1646674385
transform -1 0 25944 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1646674385
transform 1 0 24196 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1646674385
transform 1 0 24380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_264
timestamp 1646674385
transform 1 0 25392 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_270
timestamp 1646674385
transform 1 0 25944 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1646674385
transform 1 0 24288 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1663_
timestamp 1646674385
transform -1 0 25392 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1897__A
timestamp 1646674385
transform -1 0 27784 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_274
timestamp 1646674385
transform 1 0 26312 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_284
timestamp 1646674385
transform 1 0 27232 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_290
timestamp 1646674385
transform 1 0 27784 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1657_
timestamp 1646674385
transform 1 0 26404 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2196__B1
timestamp 1646674385
transform 1 0 28152 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2252__A2
timestamp 1646674385
transform -1 0 28888 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2272__A2
timestamp 1646674385
transform 1 0 29532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_296
timestamp 1646674385
transform 1 0 28336 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1646674385
transform 1 0 28888 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_311
timestamp 1646674385
transform 1 0 29716 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1646674385
transform 1 0 29440 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2273__C
timestamp 1646674385
transform 1 0 30084 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2286__A2
timestamp 1646674385
transform 1 0 30636 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2286__B2
timestamp 1646674385
transform -1 0 31372 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_317
timestamp 1646674385
transform 1 0 30268 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_323
timestamp 1646674385
transform 1 0 30820 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_329
timestamp 1646674385
transform 1 0 31372 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1646674385
transform -1 0 32016 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1946__A2
timestamp 1646674385
transform -1 0 1564 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_13
timestamp 1646674385
transform 1 0 2300 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_20
timestamp 1646674385
transform 1 0 2944 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_5
timestamp 1646674385
transform 1 0 1564 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1646674385
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1921_
timestamp 1646674385
transform 1 0 2668 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1950_
timestamp 1646674385
transform -1 0 2300 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_28
timestamp 1646674385
transform 1 0 3680 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_33
timestamp 1646674385
transform 1 0 4140 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1980_
timestamp 1646674385
transform 1 0 4508 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1983_
timestamp 1646674385
transform -1 0 4140 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1980__B
timestamp 1646674385
transform -1 0 6532 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_42
timestamp 1646674385
transform 1 0 4968 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1646674385
transform 1 0 5612 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1646674385
transform 1 0 6164 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_59
timestamp 1646674385
transform 1 0 6532 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1646674385
transform 1 0 6256 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1978_
timestamp 1646674385
transform 1 0 5336 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_71
timestamp 1646674385
transform 1 0 7636 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_78
timestamp 1646674385
transform 1 0 8280 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1936_
timestamp 1646674385
transform -1 0 8280 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1938_
timestamp 1646674385
transform -1 0 8924 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2000_
timestamp 1646674385
transform 1 0 7268 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_85
timestamp 1646674385
transform 1 0 8924 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_91
timestamp 1646674385
transform 1 0 9476 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2861_
timestamp 1646674385
transform 1 0 9568 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1646674385
transform 1 0 11040 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 1646674385
transform 1 0 11500 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1646674385
transform 1 0 11408 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1383_
timestamp 1646674385
transform -1 0 12696 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_126
timestamp 1646674385
transform 1 0 12696 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1646674385
transform 1 0 13708 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_144
timestamp 1646674385
transform 1 0 14352 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1991_
timestamp 1646674385
transform 1 0 14076 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2014_
timestamp 1646674385
transform 1 0 13064 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_57_150
timestamp 1646674385
transform 1 0 14904 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 1646674385
transform 1 0 15824 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1375_
timestamp 1646674385
transform -1 0 15824 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_57_169
timestamp 1646674385
transform 1 0 16652 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_181
timestamp 1646674385
transform 1 0 17756 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1646674385
transform 1 0 16560 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2077_
timestamp 1646674385
transform 1 0 18124 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2078_
timestamp 1646674385
transform 1 0 16928 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_57_188
timestamp 1646674385
transform 1 0 18400 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_206
timestamp 1646674385
transform 1 0 20056 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1355_
timestamp 1646674385
transform 1 0 19136 0 -1 32096
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1646674385
transform 1 0 21252 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1646674385
transform 1 0 21620 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1646674385
transform 1 0 21712 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1363_
timestamp 1646674385
transform -1 0 21252 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2875_
timestamp 1646674385
transform -1 0 23276 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1646674385
transform 1 0 23276 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2716_
timestamp 1646674385
transform -1 0 25208 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_57_262
timestamp 1646674385
transform 1 0 25208 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1667_
timestamp 1646674385
transform 1 0 25576 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1858__B
timestamp 1646674385
transform -1 0 27140 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2110__B1
timestamp 1646674385
transform 1 0 27508 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1646674385
transform 1 0 26404 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1646674385
transform 1 0 26772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_283
timestamp 1646674385
transform 1 0 27140 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_289
timestamp 1646674385
transform 1 0 27692 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1646674385
transform 1 0 26864 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2193__B1
timestamp 1646674385
transform -1 0 28244 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_295
timestamp 1646674385
transform 1 0 28244 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2712_
timestamp 1646674385
transform -1 0 30268 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_57_317
timestamp 1646674385
transform 1 0 30268 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_325
timestamp 1646674385
transform 1 0 31004 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_329
timestamp 1646674385
transform 1 0 31372 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1646674385
transform -1 0 32016 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output50
timestamp 1646674385
transform -1 0 31372 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_10
timestamp 1646674385
transform 1 0 2024 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp 1646674385
transform 1 0 1380 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1646674385
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _1946_
timestamp 1646674385
transform 1 0 2392 0 1 32096
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1948_
timestamp 1646674385
transform -1 0 2024 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1646674385
transform 1 0 3312 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_32
timestamp 1646674385
transform 1 0 4048 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_39
timestamp 1646674385
transform 1 0 4692 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1646674385
transform 1 0 3680 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1922_
timestamp 1646674385
transform 1 0 3772 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1932_
timestamp 1646674385
transform 1 0 4416 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_46
timestamp 1646674385
transform 1 0 5336 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_50
timestamp 1646674385
transform 1 0 5704 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1979_
timestamp 1646674385
transform 1 0 5060 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _2284_
timestamp 1646674385
transform -1 0 7360 0 1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_58_68
timestamp 1646674385
transform 1 0 7360 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1646674385
transform 1 0 8464 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2001_
timestamp 1646674385
transform 1 0 7728 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_88
timestamp 1646674385
transform 1 0 9200 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_95
timestamp 1646674385
transform 1 0 9844 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1646674385
transform 1 0 8832 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1388_
timestamp 1646674385
transform -1 0 11408 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1935_
timestamp 1646674385
transform -1 0 9200 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1995_
timestamp 1646674385
transform 1 0 9568 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_112
timestamp 1646674385
transform 1 0 11408 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2864_
timestamp 1646674385
transform 1 0 11776 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 1646674385
transform 1 0 13248 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1646674385
transform 1 0 13984 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _2017_
timestamp 1646674385
transform 1 0 14076 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_58_148
timestamp 1646674385
transform 1 0 14720 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_152
timestamp 1646674385
transform 1 0 15088 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_160
timestamp 1646674385
transform 1 0 15824 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1953_
timestamp 1646674385
transform -1 0 17020 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1963_
timestamp 1646674385
transform 1 0 15180 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1953__A2
timestamp 1646674385
transform 1 0 18308 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1646674385
transform 1 0 17020 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_183
timestamp 1646674385
transform 1 0 17940 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1898_
timestamp 1646674385
transform 1 0 17388 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1646674385
transform 1 0 18492 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1646674385
transform 1 0 19044 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_197
timestamp 1646674385
transform 1 0 19228 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_203
timestamp 1646674385
transform 1 0 19780 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1646674385
transform 1 0 19136 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2331_
timestamp 1646674385
transform -1 0 19780 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2332_
timestamp 1646674385
transform 1 0 20148 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_216
timestamp 1646674385
transform 1 0 20976 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_220
timestamp 1646674385
transform 1 0 21344 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1368_
timestamp 1646674385
transform 1 0 21436 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A
timestamp 1646674385
transform 1 0 22632 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_230
timestamp 1646674385
transform 1 0 22264 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_236
timestamp 1646674385
transform 1 0 22816 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1646674385
transform 1 0 23828 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1860_
timestamp 1646674385
transform 1 0 23552 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1646674385
transform 1 0 24196 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_253
timestamp 1646674385
transform 1 0 24380 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_261
timestamp 1646674385
transform 1 0 25116 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1646674385
transform 1 0 24288 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1858_
timestamp 1646674385
transform 1 0 24656 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2715_
timestamp 1646674385
transform 1 0 25484 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_281
timestamp 1646674385
transform 1 0 26956 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2713_
timestamp 1646674385
transform -1 0 28796 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1646674385
transform 1 0 28796 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1646674385
transform 1 0 29348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1646674385
transform 1 0 29440 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2711_
timestamp 1646674385
transform -1 0 31004 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_58_325
timestamp 1646674385
transform 1 0 31004 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1646674385
transform -1 0 32016 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1949_
timestamp 1646674385
transform 1 0 1748 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1947_
timestamp 1646674385
transform 1 0 1472 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1646674385
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1646674385
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1646674385
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_3
timestamp 1646674385
transform 1 0 1380 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1945_
timestamp 1646674385
transform 1 0 2852 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_60_15
timestamp 1646674385
transform 1 0 2484 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_12
timestamp 1646674385
transform 1 0 2208 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _1951_
timestamp 1646674385
transform -1 0 4140 0 -1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1945__B
timestamp 1646674385
transform 1 0 4416 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_33
timestamp 1646674385
transform 1 0 4140 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_37
timestamp 1646674385
transform 1 0 4508 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1646674385
transform 1 0 3312 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_32
timestamp 1646674385
transform 1 0 4048 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_38
timestamp 1646674385
transform 1 0 4600 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1646674385
transform 1 0 3680 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1943_
timestamp 1646674385
transform 1 0 3772 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2283_
timestamp 1646674385
transform 1 0 4600 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_42
timestamp 1646674385
transform 1 0 4968 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1646674385
transform 1 0 5704 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_52
timestamp 1646674385
transform 1 0 5888 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_61
timestamp 1646674385
transform 1 0 6716 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1646674385
transform 1 0 6256 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _2278_
timestamp 1646674385
transform 1 0 6256 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _2279_
timestamp 1646674385
transform 1 0 6348 0 -1 33184
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _2281_
timestamp 1646674385
transform 1 0 5336 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2282_
timestamp 1646674385
transform 1 0 5152 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1799__A
timestamp 1646674385
transform -1 0 7820 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_67
timestamp 1646674385
transform 1 0 7268 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_73
timestamp 1646674385
transform 1 0 7820 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_67
timestamp 1646674385
transform 1 0 7268 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_76
timestamp 1646674385
transform 1 0 8096 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1999_
timestamp 1646674385
transform 1 0 7360 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _2003_
timestamp 1646674385
transform -1 0 9752 0 -1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_59_100
timestamp 1646674385
transform 1 0 10304 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_94
timestamp 1646674385
transform 1 0 9752 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_101
timestamp 1646674385
transform 1 0 10396 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_95
timestamp 1646674385
transform 1 0 9844 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1646674385
transform 1 0 8832 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_2  _1998_
timestamp 1646674385
transform 1 0 8924 0 1 33184
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _2258_
timestamp 1646674385
transform -1 0 11040 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2259_
timestamp 1646674385
transform 1 0 10488 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2257_
timestamp 1646674385
transform -1 0 12328 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1646674385
transform 1 0 11408 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_109
timestamp 1646674385
transform 1 0 11132 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1646674385
transform 1 0 11040 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1997__B
timestamp 1646674385
transform -1 0 11684 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_122
timestamp 1646674385
transform 1 0 12328 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_121
timestamp 1646674385
transform 1 0 12236 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_115
timestamp 1646674385
transform 1 0 11684 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2004__A2
timestamp 1646674385
transform -1 0 12236 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _2004_
timestamp 1646674385
transform 1 0 12604 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1793__A
timestamp 1646674385
transform 1 0 13340 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_134
timestamp 1646674385
transform 1 0 13432 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_129
timestamp 1646674385
transform 1 0 12972 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_135
timestamp 1646674385
transform 1 0 13524 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1646674385
transform 1 0 13892 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1646674385
transform 1 0 13984 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1376_
timestamp 1646674385
transform -1 0 14628 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2256_
timestamp 1646674385
transform 1 0 12696 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2868_
timestamp 1646674385
transform 1 0 14076 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_59_147
timestamp 1646674385
transform 1 0 14628 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_160
timestamp 1646674385
transform 1 0 15824 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_157
timestamp 1646674385
transform 1 0 15548 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1374_
timestamp 1646674385
transform 1 0 14996 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2870_
timestamp 1646674385
transform 1 0 15916 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_59_176
timestamp 1646674385
transform 1 0 17296 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_177
timestamp 1646674385
transform 1 0 17388 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_184
timestamp 1646674385
transform 1 0 18032 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1646674385
transform 1 0 16560 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1952_
timestamp 1646674385
transform 1 0 17756 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1965_
timestamp 1646674385
transform 1 0 16652 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2879_
timestamp 1646674385
transform -1 0 19136 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_59_196
timestamp 1646674385
transform 1 0 19136 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_188
timestamp 1646674385
transform 1 0 18400 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1646674385
transform 1 0 18768 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_206
timestamp 1646674385
transform 1 0 20056 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1646674385
transform 1 0 19136 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1359_
timestamp 1646674385
transform -1 0 20332 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2107_
timestamp 1646674385
transform 1 0 18492 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2108_
timestamp 1646674385
transform 1 0 19228 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2110_
timestamp 1646674385
transform 1 0 20700 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2109_
timestamp 1646674385
transform 1 0 20424 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_60_217
timestamp 1646674385
transform 1 0 21068 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1646674385
transform 1 0 20332 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2339_
timestamp 1646674385
transform 1 0 21436 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1646674385
transform 1 0 21712 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1646674385
transform 1 0 21804 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1646674385
transform 1 0 21344 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1292_
timestamp 1646674385
transform 1 0 22172 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_228
timestamp 1646674385
transform 1 0 22080 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_233
timestamp 1646674385
transform 1 0 22540 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_236
timestamp 1646674385
transform 1 0 22816 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_243
timestamp 1646674385
transform 1 0 23460 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1289_
timestamp 1646674385
transform 1 0 22908 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2605_
timestamp 1646674385
transform 1 0 22908 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__o221a_1  _1669_
timestamp 1646674385
transform 1 0 24748 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1646674385
transform 1 0 24288 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1646674385
transform 1 0 24380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1646674385
transform 1 0 24196 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_259
timestamp 1646674385
transform 1 0 24932 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_253
timestamp 1646674385
transform 1 0 24380 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A
timestamp 1646674385
transform 1 0 24748 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1668_
timestamp 1646674385
transform 1 0 25392 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_266
timestamp 1646674385
transform 1 0 25576 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_263
timestamp 1646674385
transform 1 0 25300 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2714_
timestamp 1646674385
transform -1 0 27416 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1646674385
transform 1 0 26220 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1646674385
transform 1 0 26772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_286
timestamp 1646674385
transform 1 0 27416 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1646674385
transform 1 0 27416 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1646674385
transform 1 0 26864 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1672_
timestamp 1646674385
transform -1 0 28612 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1859_
timestamp 1646674385
transform -1 0 27416 0 -1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_59_292
timestamp 1646674385
transform 1 0 27968 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_303
timestamp 1646674385
transform 1 0 28980 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_299
timestamp 1646674385
transform 1 0 28612 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1646674385
transform 1 0 29348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1646674385
transform 1 0 29440 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1671_
timestamp 1646674385
transform 1 0 28060 0 -1 33184
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1674_
timestamp 1646674385
transform -1 0 30176 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1675_
timestamp 1646674385
transform 1 0 29532 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1646674385
transform 1 0 30360 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_316
timestamp 1646674385
transform 1 0 30176 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2287__C
timestamp 1646674385
transform -1 0 30728 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_324
timestamp 1646674385
transform 1 0 30912 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_328
timestamp 1646674385
transform 1 0 31280 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_322
timestamp 1646674385
transform 1 0 30728 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2288__B1
timestamp 1646674385
transform -1 0 31280 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2259__B1
timestamp 1646674385
transform -1 0 30912 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1646674385
transform -1 0 32016 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1646674385
transform -1 0 32016 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_332
timestamp 1646674385
transform 1 0 31648 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_332
timestamp 1646674385
transform 1 0 31648 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_7
timestamp 1646674385
transform 1 0 1748 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1646674385
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2597_
timestamp 1646674385
transform -1 0 3128 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1646674385
transform 1 0 1380 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_22
timestamp 1646674385
transform 1 0 3128 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_26
timestamp 1646674385
transform 1 0 3496 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_33
timestamp 1646674385
transform 1 0 4140 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_40
timestamp 1646674385
transform 1 0 4784 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1489_
timestamp 1646674385
transform -1 0 4140 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2246_
timestamp 1646674385
transform -1 0 4784 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1646674385
transform 1 0 5888 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1646674385
transform 1 0 6256 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _2280_
timestamp 1646674385
transform -1 0 5888 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2589_
timestamp 1646674385
transform 1 0 6348 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_61_66
timestamp 1646674385
transform 1 0 7176 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_78
timestamp 1646674385
transform 1 0 8280 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1799_
timestamp 1646674385
transform 1 0 7912 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2583_
timestamp 1646674385
transform -1 0 9476 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_61_104
timestamp 1646674385
transform 1 0 10672 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_91
timestamp 1646674385
transform 1 0 9476 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1997_
timestamp 1646674385
transform -1 0 10672 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_61_113
timestamp 1646674385
transform 1 0 11500 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_117
timestamp 1646674385
transform 1 0 11868 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_124
timestamp 1646674385
transform 1 0 12512 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1646674385
transform 1 0 11408 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _1793_
timestamp 1646674385
transform -1 0 12512 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1789__A
timestamp 1646674385
transform 1 0 12880 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_130
timestamp 1646674385
transform 1 0 13064 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_prog_clk
timestamp 1646674385
transform 1 0 13432 0 -1 34272
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_61_154
timestamp 1646674385
transform 1 0 15272 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1646674385
transform 1 0 15916 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2020_
timestamp 1646674385
transform -1 0 15916 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1965__B1
timestamp 1646674385
transform -1 0 16836 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1987__C
timestamp 1646674385
transform 1 0 17204 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2017__B1
timestamp 1646674385
transform -1 0 17940 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1646674385
transform 1 0 16468 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_171
timestamp 1646674385
transform 1 0 16836 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_177
timestamp 1646674385
transform 1 0 17388 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_183
timestamp 1646674385
transform 1 0 17940 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1646674385
transform 1 0 16560 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_200
timestamp 1646674385
transform 1 0 19504 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_204
timestamp 1646674385
transform 1 0 19872 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1358_
timestamp 1646674385
transform 1 0 18676 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1360_
timestamp 1646674385
transform 1 0 19964 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2078__B2
timestamp 1646674385
transform 1 0 21160 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_214
timestamp 1646674385
transform 1 0 20792 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1646674385
transform 1 0 21344 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1646674385
transform 1 0 21712 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2338_
timestamp 1646674385
transform -1 0 22632 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_61_234
timestamp 1646674385
transform 1 0 22632 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_240
timestamp 1646674385
transform 1 0 23184 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1646674385
transform 1 0 23920 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2192_
timestamp 1646674385
transform 1 0 23276 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_61_264
timestamp 1646674385
transform 1 0 25392 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _2191_
timestamp 1646674385
transform 1 0 25760 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _2193_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 24288 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1646674385
transform 1 0 26496 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1646674385
transform 1 0 26956 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_285
timestamp 1646674385
transform 1 0 27324 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_289
timestamp 1646674385
transform 1 0 27692 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1646674385
transform 1 0 26864 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2140_
timestamp 1646674385
transform 1 0 27416 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_296
timestamp 1646674385
transform 1 0 28336 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_302
timestamp 1646674385
transform 1 0 28888 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_312
timestamp 1646674385
transform 1 0 29808 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1677_
timestamp 1646674385
transform 1 0 28980 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2139_
timestamp 1646674385
transform -1 0 28336 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_319
timestamp 1646674385
transform 1 0 30452 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_325
timestamp 1646674385
transform 1 0 31004 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_329
timestamp 1646674385
transform 1 0 31372 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1646674385
transform -1 0 32016 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2142_
timestamp 1646674385
transform -1 0 30452 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output39
timestamp 1646674385
transform -1 0 31372 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1947__A2
timestamp 1646674385
transform -1 0 1656 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_13
timestamp 1646674385
transform 1 0 2300 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_3
timestamp 1646674385
transform 1 0 1380 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_6
timestamp 1646674385
transform 1 0 1656 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1646674385
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1491_
timestamp 1646674385
transform 1 0 2668 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1919_
timestamp 1646674385
transform -1 0 2300 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1646674385
transform 1 0 3036 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1646674385
transform 1 0 3588 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1646674385
transform 1 0 3772 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_41
timestamp 1646674385
transform 1 0 4876 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1646674385
transform 1 0 3680 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1499_
timestamp 1646674385
transform -1 0 4876 0 1 34272
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1999__A2
timestamp 1646674385
transform 1 0 5888 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_48
timestamp 1646674385
transform 1 0 5520 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_54
timestamp 1646674385
transform 1 0 6072 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_62
timestamp 1646674385
transform 1 0 6808 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2002_
timestamp 1646674385
transform 1 0 6440 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2243_
timestamp 1646674385
transform -1 0 5520 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_75
timestamp 1646674385
transform 1 0 8004 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1646674385
transform 1 0 8740 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1523_
timestamp 1646674385
transform 1 0 7176 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_62_103
timestamp 1646674385
transform 1 0 10580 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_95
timestamp 1646674385
transform 1 0 9844 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1646674385
transform 1 0 8832 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1521_
timestamp 1646674385
transform 1 0 8924 0 1 34272
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1794_
timestamp 1646674385
transform -1 0 10580 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_110
timestamp 1646674385
transform 1 0 11224 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_120
timestamp 1646674385
transform 1 0 12144 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1789_
timestamp 1646674385
transform -1 0 12144 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1996_
timestamp 1646674385
transform 1 0 10948 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_128
timestamp 1646674385
transform 1 0 12880 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1646674385
transform 1 0 13616 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_141
timestamp 1646674385
transform 1 0 14076 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1646674385
transform 1 0 13984 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1987_
timestamp 1646674385
transform 1 0 14352 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2021_
timestamp 1646674385
transform 1 0 12972 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_62_151
timestamp 1646674385
transform 1 0 14996 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_164
timestamp 1646674385
transform 1 0 16192 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1377_
timestamp 1646674385
transform -1 0 16192 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_62_172
timestamp 1646674385
transform 1 0 16928 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_178
timestamp 1646674385
transform 1 0 17480 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2115_
timestamp 1646674385
transform 1 0 17572 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_prog_clk
timestamp 1646674385
transform 1 0 16560 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2020__A
timestamp 1646674385
transform -1 0 19412 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1646674385
transform 1 0 18768 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_199
timestamp 1646674385
transform 1 0 19412 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1646674385
transform 1 0 19136 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2877_
timestamp 1646674385
transform 1 0 20148 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_62_223
timestamp 1646674385
transform 1 0 21620 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2878_
timestamp 1646674385
transform 1 0 21988 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_243
timestamp 1646674385
transform 1 0 23460 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1646674385
transform 1 0 24196 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1646674385
transform 1 0 24380 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_257
timestamp 1646674385
transform 1 0 24748 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_267
timestamp 1646674385
transform 1 0 25668 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1646674385
transform 1 0 24288 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1666_
timestamp 1646674385
transform 1 0 24840 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_62_274
timestamp 1646674385
transform 1 0 26312 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_286
timestamp 1646674385
transform 1 0 27416 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1665_
timestamp 1646674385
transform -1 0 27416 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2111_
timestamp 1646674385
transform 1 0 26036 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1646674385
transform 1 0 29072 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1646674385
transform 1 0 29440 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1673_
timestamp 1646674385
transform -1 0 29072 0 1 34272
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2710_
timestamp 1646674385
transform -1 0 31004 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_325
timestamp 1646674385
transform 1 0 31004 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1646674385
transform -1 0 32016 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_13
timestamp 1646674385
transform 1 0 2300 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_20
timestamp 1646674385
transform 1 0 2944 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1646674385
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1646674385
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1944_
timestamp 1646674385
transform 1 0 2668 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1646674385
transform -1 0 2300 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_40
timestamp 1646674385
transform 1 0 4784 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2807_
timestamp 1646674385
transform 1 0 3312 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1646674385
transform 1 0 5428 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1646674385
transform 1 0 6164 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_60
timestamp 1646674385
transform 1 0 6624 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1646674385
transform 1 0 6256 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2244_
timestamp 1646674385
transform -1 0 5428 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2245_
timestamp 1646674385
transform 1 0 6348 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1523__C1
timestamp 1646674385
transform -1 0 7176 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_66
timestamp 1646674385
transform 1 0 7176 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2799_
timestamp 1646674385
transform 1 0 7544 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_86
timestamp 1646674385
transform 1 0 9016 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_90
timestamp 1646674385
transform 1 0 9384 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2638_
timestamp 1646674385
transform -1 0 10948 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_107
timestamp 1646674385
transform 1 0 10948 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1646674385
transform 1 0 11316 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_113
timestamp 1646674385
transform 1 0 11500 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_117
timestamp 1646674385
transform 1 0 11868 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1646674385
transform 1 0 11408 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2602_
timestamp 1646674385
transform -1 0 13432 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_134
timestamp 1646674385
transform 1 0 13432 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_141
timestamp 1646674385
transform 1 0 14076 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1869_
timestamp 1646674385
transform 1 0 13800 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1977__A2
timestamp 1646674385
transform 1 0 15916 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_147
timestamp 1646674385
transform 1 0 14628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_157
timestamp 1646674385
transform 1 0 15548 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_163
timestamp 1646674385
transform 1 0 16100 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1977_
timestamp 1646674385
transform 1 0 14720 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1646674385
transform 1 0 16468 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_185
timestamp 1646674385
transform 1 0 18124 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1646674385
transform 1 0 16560 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2603_
timestamp 1646674385
transform 1 0 16652 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_196
timestamp 1646674385
transform 1 0 19136 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_200
timestamp 1646674385
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1361_
timestamp 1646674385
transform 1 0 19596 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _2113_
timestamp 1646674385
transform -1 0 19136 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_63_210
timestamp 1646674385
transform 1 0 20424 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_216
timestamp 1646674385
transform 1 0 20976 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1646674385
transform 1 0 21344 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_228
timestamp 1646674385
transform 1 0 22080 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1646674385
transform 1 0 21712 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2336_
timestamp 1646674385
transform -1 0 22080 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2337_
timestamp 1646674385
transform 1 0 21068 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_248
timestamp 1646674385
transform 1 0 23920 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2604_
timestamp 1646674385
transform 1 0 22448 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1664__A
timestamp 1646674385
transform 1 0 24288 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_254
timestamp 1646674385
transform 1 0 24472 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2717_
timestamp 1646674385
transform -1 0 26312 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1646674385
transform 1 0 26312 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_286
timestamp 1646674385
transform 1 0 27416 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1646674385
transform 1 0 26864 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _2138_
timestamp 1646674385
transform -1 0 27416 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_63_302
timestamp 1646674385
transform 1 0 28888 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_308
timestamp 1646674385
transform 1 0 29440 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1670_
timestamp 1646674385
transform 1 0 27968 0 -1 35360
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2709_
timestamp 1646674385
transform -1 0 31004 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_63_325
timestamp 1646674385
transform 1 0 31004 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1646674385
transform -1 0 32016 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2039__A2
timestamp 1646674385
transform -1 0 1656 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1646674385
transform 1 0 2944 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_3
timestamp 1646674385
transform 1 0 1380 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_6
timestamp 1646674385
transform 1 0 1656 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1646674385
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1493_
timestamp 1646674385
transform -1 0 2944 0 1 35360
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_64_38
timestamp 1646674385
transform 1 0 4600 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1646674385
transform 1 0 3680 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1506_
timestamp 1646674385
transform -1 0 4600 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_64_46
timestamp 1646674385
transform 1 0 5336 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_54
timestamp 1646674385
transform 1 0 6072 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_58
timestamp 1646674385
transform 1 0 6440 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1428_
timestamp 1646674385
transform 1 0 6808 0 1 35360
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1502_
timestamp 1646674385
transform -1 0 5336 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2276_
timestamp 1646674385
transform -1 0 6440 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_72
timestamp 1646674385
transform 1 0 7728 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 1646674385
transform 1 0 8372 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1646674385
transform 1 0 8740 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2277_
timestamp 1646674385
transform 1 0 8096 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1790__A
timestamp 1646674385
transform 1 0 9108 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_102
timestamp 1646674385
transform 1 0 10488 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1646674385
transform 1 0 8924 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_89
timestamp 1646674385
transform 1 0 9292 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1646674385
transform 1 0 8832 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1801_
timestamp 1646674385
transform 1 0 9660 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1794__A
timestamp 1646674385
transform -1 0 11040 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_108
timestamp 1646674385
transform 1 0 11040 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_121
timestamp 1646674385
transform 1 0 12236 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1868_
timestamp 1646674385
transform 1 0 11776 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_64_136
timestamp 1646674385
transform 1 0 13616 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_141
timestamp 1646674385
transform 1 0 14076 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_145
timestamp 1646674385
transform 1 0 14444 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1646674385
transform 1 0 13984 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1976_
timestamp 1646674385
transform -1 0 14444 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _2022_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform 1 0 12972 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_64_165
timestamp 1646674385
transform 1 0 16284 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2867_
timestamp 1646674385
transform -1 0 16284 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_64_169
timestamp 1646674385
transform 1 0 16652 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_173
timestamp 1646674385
transform 1 0 17020 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1646674385
transform 1 0 18124 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1866_
timestamp 1646674385
transform -1 0 17020 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _2114_
timestamp 1646674385
transform 1 0 17388 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2078__A2
timestamp 1646674385
transform 1 0 18492 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_191
timestamp 1646674385
transform 1 0 18676 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1646674385
transform 1 0 19044 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1646674385
transform 1 0 19136 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2880_
timestamp 1646674385
transform 1 0 19228 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_213
timestamp 1646674385
transform 1 0 20700 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_222
timestamp 1646674385
transform 1 0 21528 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_228
timestamp 1646674385
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1863_
timestamp 1646674385
transform -1 0 22448 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2340_
timestamp 1646674385
transform -1 0 21528 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_232
timestamp 1646674385
transform 1 0 22448 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1646674385
transform 1 0 23920 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1925_
timestamp 1646674385
transform 1 0 22816 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1646674385
transform 1 0 24380 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_261
timestamp 1646674385
transform 1 0 25116 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_269
timestamp 1646674385
transform 1 0 25852 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1646674385
transform 1 0 24288 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1660_
timestamp 1646674385
transform 1 0 24748 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1661_
timestamp 1646674385
transform -1 0 25852 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_277
timestamp 1646674385
transform 1 0 26588 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_283
timestamp 1646674385
transform 1 0 27140 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2121_
timestamp 1646674385
transform -1 0 27140 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2144_
timestamp 1646674385
transform -1 0 28336 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_296
timestamp 1646674385
transform 1 0 28336 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_303
timestamp 1646674385
transform 1 0 28980 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1646674385
transform 1 0 29348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1646674385
transform 1 0 29440 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1676_
timestamp 1646674385
transform 1 0 29532 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2133_
timestamp 1646674385
transform -1 0 28980 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2323__B2
timestamp 1646674385
transform -1 0 30912 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_318
timestamp 1646674385
transform 1 0 30360 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_324
timestamp 1646674385
transform 1 0 30912 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_332
timestamp 1646674385
transform 1 0 31648 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1646674385
transform -1 0 32016 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_19
timestamp 1646674385
transform 1 0 2852 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1646674385
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2814_
timestamp 1646674385
transform 1 0 1380 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_31
timestamp 1646674385
transform 1 0 3956 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1501_
timestamp 1646674385
transform -1 0 3956 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1505_
timestamp 1646674385
transform 1 0 4324 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__A
timestamp 1646674385
transform -1 0 5704 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_44
timestamp 1646674385
transform 1 0 5152 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_50
timestamp 1646674385
transform 1 0 5704 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_61
timestamp 1646674385
transform 1 0 6716 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1646674385
transform 1 0 6256 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1504_
timestamp 1646674385
transform -1 0 6716 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1526__C1
timestamp 1646674385
transform 1 0 8280 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_74
timestamp 1646674385
transform 1 0 7912 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_80
timestamp 1646674385
transform 1 0 8464 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1526_
timestamp 1646674385
transform -1 0 7912 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_65_84
timestamp 1646674385
transform 1 0 8832 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_95
timestamp 1646674385
transform 1 0 9844 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1790_
timestamp 1646674385
transform 1 0 8924 0 -1 36448
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2596_
timestamp 1646674385
transform -1 0 11040 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_65_108
timestamp 1646674385
transform 1 0 11040 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1646674385
transform 1 0 11500 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_120
timestamp 1646674385
transform 1 0 12144 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1646674385
transform 1 0 11408 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1867_
timestamp 1646674385
transform 1 0 11684 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_65_128
timestamp 1646674385
transform 1 0 12880 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _2657_
timestamp 1646674385
transform 1 0 12972 0 -1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_65_146
timestamp 1646674385
transform 1 0 14536 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_154
timestamp 1646674385
transform 1 0 15272 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_162
timestamp 1646674385
transform 1 0 16008 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1988_
timestamp 1646674385
transform 1 0 15364 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_65_174
timestamp 1646674385
transform 1 0 17112 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_187
timestamp 1646674385
transform 1 0 18308 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1646674385
transform 1 0 16560 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1735_
timestamp 1646674385
transform 1 0 17480 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1865_
timestamp 1646674385
transform -1 0 17112 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1988__B1
timestamp 1646674385
transform 1 0 18676 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2108__B2
timestamp 1646674385
transform -1 0 19412 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2109__C
timestamp 1646674385
transform 1 0 20240 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_193
timestamp 1646674385
transform 1 0 18860 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_199
timestamp 1646674385
transform 1 0 19412 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_207
timestamp 1646674385
transform 1 0 20148 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_210
timestamp 1646674385
transform 1 0 20424 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_216
timestamp 1646674385
transform 1 0 20976 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1646674385
transform 1 0 21344 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1646674385
transform 1 0 21712 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2334_
timestamp 1646674385
transform -1 0 21344 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2349_
timestamp 1646674385
transform 1 0 21804 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1861__B
timestamp 1646674385
transform 1 0 22632 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_230
timestamp 1646674385
transform 1 0 22264 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_236
timestamp 1646674385
transform 1 0 22816 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_247
timestamp 1646674385
transform 1 0 23828 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1924_
timestamp 1646674385
transform 1 0 23184 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1660__A
timestamp 1646674385
transform 1 0 25116 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_255
timestamp 1646674385
transform 1 0 24564 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_263
timestamp 1646674385
transform 1 0 25300 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1664_
timestamp 1646674385
transform 1 0 24196 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2588_
timestamp 1646674385
transform 1 0 25668 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1646674385
transform 1 0 26496 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_289
timestamp 1646674385
transform 1 0 27692 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1646674385
transform 1 0 26864 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _2149_
timestamp 1646674385
transform 1 0 26956 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2323__A2
timestamp 1646674385
transform -1 0 29900 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_300
timestamp 1646674385
transform 1 0 28704 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_307
timestamp 1646674385
transform 1 0 29348 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2141_
timestamp 1646674385
transform -1 0 29348 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2143_
timestamp 1646674385
transform 1 0 28060 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2324__C
timestamp 1646674385
transform -1 0 30452 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_313
timestamp 1646674385
transform 1 0 29900 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_319
timestamp 1646674385
transform 1 0 30452 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_325
timestamp 1646674385
transform 1 0 31004 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_329
timestamp 1646674385
transform 1 0 31372 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1646674385
transform -1 0 32016 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output51
timestamp 1646674385
transform -1 0 31372 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1494_
timestamp 1646674385
transform -1 0 2484 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1646674385
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1646674385
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_5
timestamp 1646674385
transform 1 0 1564 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_3
timestamp 1646674385
transform 1 0 1380 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2181__A2
timestamp 1646674385
transform -1 0 1564 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__B2
timestamp 1646674385
transform 1 0 1932 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_11
timestamp 1646674385
transform 1 0 2116 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_19
timestamp 1646674385
transform 1 0 2852 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_15
timestamp 1646674385
transform 1 0 2484 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__A
timestamp 1646674385
transform -1 0 3128 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2809_
timestamp 1646674385
transform -1 0 3956 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_66_22
timestamp 1646674385
transform 1 0 3128 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_39
timestamp 1646674385
transform 1 0 4692 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_31
timestamp 1646674385
transform 1 0 3956 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_35
timestamp 1646674385
transform 1 0 4324 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1646674385
transform 1 0 3680 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1492_
timestamp 1646674385
transform 1 0 3772 0 1 36448
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _2806_
timestamp 1646674385
transform 1 0 4416 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_66_61
timestamp 1646674385
transform 1 0 6716 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 1646674385
transform 1 0 5888 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_57
timestamp 1646674385
transform 1 0 6348 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1646674385
transform 1 0 6256 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2796_
timestamp 1646674385
transform 1 0 6624 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2808_
timestamp 1646674385
transform 1 0 5244 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1801__B2
timestamp 1646674385
transform -1 0 8464 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2097__A1
timestamp 1646674385
transform 1 0 7084 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2100__A2
timestamp 1646674385
transform -1 0 7820 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_67
timestamp 1646674385
transform 1 0 7268 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_73
timestamp 1646674385
transform 1 0 7820 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_77
timestamp 1646674385
transform 1 0 8188 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1646674385
transform 1 0 8464 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_76
timestamp 1646674385
transform 1 0 8096 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2639_
timestamp 1646674385
transform -1 0 9936 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_66_94
timestamp 1646674385
transform 1 0 9752 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_104
timestamp 1646674385
transform 1 0 10672 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_96
timestamp 1646674385
transform 1 0 9936 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1646674385
transform 1 0 8832 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1798_
timestamp 1646674385
transform 1 0 8924 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _2320_
timestamp 1646674385
transform 1 0 10304 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2655_
timestamp 1646674385
transform 1 0 10488 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1801__C1
timestamp 1646674385
transform -1 0 11684 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_118
timestamp 1646674385
transform 1 0 11960 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_122
timestamp 1646674385
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_115
timestamp 1646674385
transform 1 0 11684 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1646674385
transform 1 0 11408 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1768_
timestamp 1646674385
transform 1 0 12420 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _2656_
timestamp 1646674385
transform 1 0 12052 0 -1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1768__A1
timestamp 1646674385
transform 1 0 14076 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2021__B
timestamp 1646674385
transform -1 0 14168 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_132
timestamp 1646674385
transform 1 0 13248 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_143
timestamp 1646674385
transform 1 0 14260 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_136
timestamp 1646674385
transform 1 0 13616 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_142
timestamp 1646674385
transform 1 0 14168 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1646674385
transform 1 0 13984 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2046_
timestamp 1646674385
transform 1 0 15364 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_67_151
timestamp 1646674385
transform 1 0 14996 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_148
timestamp 1646674385
transform 1 0 14720 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_149
timestamp 1646674385
transform 1 0 14812 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2115__B1
timestamp 1646674385
transform -1 0 14996 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1867__B
timestamp 1646674385
transform -1 0 14812 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_160
timestamp 1646674385
transform 1 0 15824 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_159
timestamp 1646674385
transform 1 0 15732 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1977__B2
timestamp 1646674385
transform -1 0 15732 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2677_
timestamp 1646674385
transform 1 0 16284 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2081__B1
timestamp 1646674385
transform -1 0 18308 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_181
timestamp 1646674385
transform 1 0 17756 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_187
timestamp 1646674385
transform 1 0 18308 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_173
timestamp 1646674385
transform 1 0 17020 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_179
timestamp 1646674385
transform 1 0 17572 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1646674385
transform 1 0 16560 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _2076_
timestamp 1646674385
transform 1 0 16652 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2676_
timestamp 1646674385
transform 1 0 17664 0 -1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1646674385
transform 1 0 19044 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_206
timestamp 1646674385
transform 1 0 20056 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_197
timestamp 1646674385
transform 1 0 19228 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1646674385
transform 1 0 19136 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1732_
timestamp 1646674385
transform 1 0 19228 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2678_
timestamp 1646674385
transform 1 0 19596 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_66_214
timestamp 1646674385
transform 1 0 20792 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_220
timestamp 1646674385
transform 1 0 21344 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_229
timestamp 1646674385
transform 1 0 22172 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1646674385
transform 1 0 21068 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1646674385
transform 1 0 21620 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1646674385
transform 1 0 21712 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2335_
timestamp 1646674385
transform 1 0 21712 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2341_
timestamp 1646674385
transform -1 0 21344 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2342_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646674385
transform -1 0 22448 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1646674385
transform 1 0 23644 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_232
timestamp 1646674385
transform 1 0 22448 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_241
timestamp 1646674385
transform 1 0 23276 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_245
timestamp 1646674385
transform 1 0 23644 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_249
timestamp 1646674385
transform 1 0 24012 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1861_
timestamp 1646674385
transform 1 0 22816 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _1923_
timestamp 1646674385
transform 1 0 22908 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2369_
timestamp 1646674385
transform 1 0 23736 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1925__B1
timestamp 1646674385
transform -1 0 25392 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1646674385
transform 1 0 24196 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_258
timestamp 1646674385
transform 1 0 24840 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_264
timestamp 1646674385
transform 1 0 25392 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_270
timestamp 1646674385
transform 1 0 25944 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1646674385
transform 1 0 24288 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _1862_
timestamp 1646674385
transform -1 0 24840 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _2151_
timestamp 1646674385
transform -1 0 26128 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2696_
timestamp 1646674385
transform 1 0 24380 0 -1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__o311a_1  _2150_
timestamp 1646674385
transform 1 0 26496 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1646674385
transform 1 0 26864 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1646674385
transform 1 0 26496 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_272
timestamp 1646674385
transform 1 0 26128 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2105__A
timestamp 1646674385
transform 1 0 26312 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _2122_
timestamp 1646674385
transform 1 0 27600 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2120_
timestamp 1646674385
transform -1 0 27232 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_284
timestamp 1646674385
transform 1 0 27232 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_290
timestamp 1646674385
transform 1 0 27784 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_284
timestamp 1646674385
transform 1 0 27232 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2137_
timestamp 1646674385
transform 1 0 27876 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_67_291
timestamp 1646674385
transform 1 0 27876 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_300
timestamp 1646674385
transform 1 0 28704 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_312
timestamp 1646674385
transform 1 0 29808 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_295
timestamp 1646674385
transform 1 0 28244 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_306
timestamp 1646674385
transform 1 0 29256 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1646674385
transform 1 0 29440 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1679_
timestamp 1646674385
transform 1 0 28336 0 -1 37536
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2132_
timestamp 1646674385
transform -1 0 29808 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2135_
timestamp 1646674385
transform -1 0 29900 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_319
timestamp 1646674385
transform 1 0 30452 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_313
timestamp 1646674385
transform 1 0 29900 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_318
timestamp 1646674385
transform 1 0 30360 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2325__B1
timestamp 1646674385
transform -1 0 30360 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2129__B
timestamp 1646674385
transform 1 0 30268 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output40
timestamp 1646674385
transform -1 0 31372 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_329
timestamp 1646674385
transform 1 0 31372 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_325
timestamp 1646674385
transform 1 0 31004 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_324
timestamp 1646674385
transform 1 0 30912 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2327__A2
timestamp 1646674385
transform -1 0 30912 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1646674385
transform -1 0 32016 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1646674385
transform -1 0 32016 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_332
timestamp 1646674385
transform 1 0 31648 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__B1
timestamp 1646674385
transform 1 0 2668 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_13
timestamp 1646674385
transform 1 0 2300 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_19
timestamp 1646674385
transform 1 0 2852 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1646674385
transform 1 0 1380 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1646674385
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1646674385
transform 1 0 1748 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1646674385
transform 1 0 3588 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_38
timestamp 1646674385
transform 1 0 4600 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1646674385
transform 1 0 3680 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1503_
timestamp 1646674385
transform -1 0 4600 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1969__B
timestamp 1646674385
transform 1 0 6256 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1970__A2
timestamp 1646674385
transform 1 0 4968 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1972__A2
timestamp 1646674385
transform 1 0 5520 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_44
timestamp 1646674385
transform 1 0 5152 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_50
timestamp 1646674385
transform 1 0 5704 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_58
timestamp 1646674385
transform 1 0 6440 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1974_
timestamp 1646674385
transform 1 0 6808 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1974__A2
timestamp 1646674385
transform 1 0 7544 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2101__A1
timestamp 1646674385
transform -1 0 8280 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_66
timestamp 1646674385
transform 1 0 7176 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_72
timestamp 1646674385
transform 1 0 7728 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_78
timestamp 1646674385
transform 1 0 8280 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_88
timestamp 1646674385
transform 1 0 9200 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_92
timestamp 1646674385
transform 1 0 9568 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_98
timestamp 1646674385
transform 1 0 10120 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1646674385
transform 1 0 8832 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1770_
timestamp 1646674385
transform -1 0 11316 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2295_
timestamp 1646674385
transform -1 0 10120 0 1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2315_
timestamp 1646674385
transform 1 0 8924 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_111
timestamp 1646674385
transform 1 0 11316 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_124
timestamp 1646674385
transform 1 0 12512 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1769_
timestamp 1646674385
transform 1 0 11684 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1730__A
timestamp 1646674385
transform 1 0 14076 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1746__A
timestamp 1646674385
transform 1 0 12880 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2180__A2
timestamp 1646674385
transform -1 0 13616 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_130
timestamp 1646674385
transform 1 0 13064 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1646674385
transform 1 0 13616 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_143
timestamp 1646674385
transform 1 0 14260 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1646674385
transform 1 0 13984 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1864__B
timestamp 1646674385
transform -1 0 16560 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_150
timestamp 1646674385
transform 1 0 14904 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_162
timestamp 1646674385
transform 1 0 16008 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2018_
timestamp 1646674385
transform 1 0 14628 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2074_
timestamp 1646674385
transform 1 0 15272 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_168
timestamp 1646674385
transform 1 0 16560 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_181
timestamp 1646674385
transform 1 0 17756 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1734_
timestamp 1646674385
transform -1 0 17756 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1646674385
transform 1 0 18768 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_197
timestamp 1646674385
transform 1 0 19228 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_207
timestamp 1646674385
transform 1 0 20148 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1646674385
transform 1 0 19136 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1728_
timestamp 1646674385
transform 1 0 19320 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2370_
timestamp 1646674385
transform 1 0 18492 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1703__A
timestamp 1646674385
transform 1 0 20516 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_213
timestamp 1646674385
transform 1 0 20700 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_220
timestamp 1646674385
transform 1 0 21344 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2343_
timestamp 1646674385
transform -1 0 21344 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2593_
timestamp 1646674385
transform -1 0 22540 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_68_233
timestamp 1646674385
transform 1 0 22540 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1646674385
transform 1 0 23920 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1700_
timestamp 1646674385
transform 1 0 23092 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1646674385
transform 1 0 24380 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1646674385
transform 1 0 24288 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2697_
timestamp 1646674385
transform -1 0 26220 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_273
timestamp 1646674385
transform 1 0 26220 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_280
timestamp 1646674385
transform 1 0 26864 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_291
timestamp 1646674385
transform 1 0 27876 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2105_
timestamp 1646674385
transform -1 0 26864 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2136_
timestamp 1646674385
transform -1 0 27876 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_68_304
timestamp 1646674385
transform 1 0 29072 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1646674385
transform 1 0 29440 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1680_
timestamp 1646674385
transform 1 0 28244 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2708_
timestamp 1646674385
transform 1 0 29532 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_68_325
timestamp 1646674385
transform 1 0 31004 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1646674385
transform -1 0 32016 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_16
timestamp 1646674385
transform 1 0 2576 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1646674385
transform 1 0 1380 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1646674385
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1496_
timestamp 1646674385
transform -1 0 2576 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_69_22
timestamp 1646674385
transform 1 0 3128 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_26
timestamp 1646674385
transform 1 0 3496 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_39
timestamp 1646674385
transform 1 0 4692 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1507_
timestamp 1646674385
transform 1 0 3864 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1888_
timestamp 1646674385
transform 1 0 3220 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_49
timestamp 1646674385
transform 1 0 5612 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1646674385
transform 1 0 6164 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_57
timestamp 1646674385
transform 1 0 6348 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1646674385
transform 1 0 6256 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1972_
timestamp 1646674385
transform -1 0 5612 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2640_
timestamp 1646674385
transform 1 0 6716 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_77
timestamp 1646674385
transform 1 0 8188 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1797_
timestamp 1646674385
transform -1 0 9384 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_69_101
timestamp 1646674385
transform 1 0 10396 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_90
timestamp 1646674385
transform 1 0 9384 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _2316_
timestamp 1646674385
transform -1 0 10396 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_69_108
timestamp 1646674385
transform 1 0 11040 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_116
timestamp 1646674385
transform 1 0 11776 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1646674385
transform 1 0 11408 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1766_
timestamp 1646674385
transform 1 0 12144 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2255_
timestamp 1646674385
transform -1 0 11040 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2260_
timestamp 1646674385
transform 1 0 11500 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_129
timestamp 1646674385
transform 1 0 12972 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2658_
timestamp 1646674385
transform 1 0 13340 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_149
timestamp 1646674385
transform 1 0 14812 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_153
timestamp 1646674385
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_163
timestamp 1646674385
transform 1 0 16100 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2585_
timestamp 1646674385
transform -1 0 16100 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1646674385
transform 1 0 16468 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_174
timestamp 1646674385
transform 1 0 17112 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_187
timestamp 1646674385
transform 1 0 18308 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1646674385
transform 1 0 16560 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1736_
timestamp 1646674385
transform 1 0 17480 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1864_
timestamp 1646674385
transform -1 0 17112 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_69_194
timestamp 1646674385
transform 1 0 18952 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_202
timestamp 1646674385
transform 1 0 19688 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _2047_
timestamp 1646674385
transform 1 0 18676 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2679_
timestamp 1646674385
transform 1 0 19780 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_219
timestamp 1646674385
transform 1 0 21252 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1646674385
transform 1 0 21620 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_225
timestamp 1646674385
transform 1 0 21804 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1646674385
transform 1 0 21712 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _2375_
timestamp 1646674385
transform 1 0 21988 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_231
timestamp 1646674385
transform 1 0 22356 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_235
timestamp 1646674385
transform 1 0 22724 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2695_
timestamp 1646674385
transform -1 0 24288 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_252
timestamp 1646674385
transform 1 0 24288 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_265
timestamp 1646674385
transform 1 0 25484 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1699_
timestamp 1646674385
transform 1 0 24656 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 1646674385
transform 1 0 26496 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_281
timestamp 1646674385
transform 1 0 26956 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_290
timestamp 1646674385
transform 1 0 27784 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1646674385
transform 1 0 26864 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _2106_
timestamp 1646674385
transform 1 0 27324 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2124_
timestamp 1646674385
transform -1 0 26496 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_69_303
timestamp 1646674385
transform 1 0 28980 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1682_
timestamp 1646674385
transform 1 0 28152 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2707_
timestamp 1646674385
transform 1 0 29348 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2124__A
timestamp 1646674385
transform -1 0 31372 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_323
timestamp 1646674385
transform 1 0 30820 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_329
timestamp 1646674385
transform 1 0 31372 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1646674385
transform -1 0 32016 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1646674385
transform 1 0 2852 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1646674385
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2812_
timestamp 1646674385
transform 1 0 1380 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__B2
timestamp 1646674385
transform 1 0 3772 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1646674385
transform 1 0 3588 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_31
timestamp 1646674385
transform 1 0 3956 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1646674385
transform 1 0 3680 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_prog_clk
timestamp 1646674385
transform 1 0 4508 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_70_57
timestamp 1646674385
transform 1 0 6348 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1969_
timestamp 1646674385
transform -1 0 7176 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_70_66
timestamp 1646674385
transform 1 0 7176 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_70
timestamp 1646674385
transform 1 0 7544 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_80
timestamp 1646674385
transform 1 0 8464 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1796_
timestamp 1646674385
transform 1 0 7636 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_70_100
timestamp 1646674385
transform 1 0 10304 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_85
timestamp 1646674385
transform 1 0 8924 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_91
timestamp 1646674385
transform 1 0 9476 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1646674385
transform 1 0 8832 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _2261_
timestamp 1646674385
transform -1 0 10304 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2298_
timestamp 1646674385
transform -1 0 9476 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_70_106
timestamp 1646674385
transform 1 0 10856 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_123
timestamp 1646674385
transform 1 0 12420 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2654_
timestamp 1646674385
transform -1 0 12420 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_136
timestamp 1646674385
transform 1 0 13616 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_70_141
timestamp 1646674385
transform 1 0 14076 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1646674385
transform 1 0 13984 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1771_
timestamp 1646674385
transform -1 0 13616 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2045_
timestamp 1646674385
transform -1 0 14628 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_147
timestamp 1646674385
transform 1 0 14628 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_159
timestamp 1646674385
transform 1 0 15732 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _2075_
timestamp 1646674385
transform -1 0 15732 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_177
timestamp 1646674385
transform 1 0 17388 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1726_
timestamp 1646674385
transform -1 0 18768 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1731_
timestamp 1646674385
transform 1 0 16468 0 1 38624
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1646674385
transform 1 0 18768 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_207
timestamp 1646674385
transform 1 0 20148 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1646674385
transform 1 0 19136 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1703_
timestamp 1646674385
transform -1 0 20148 0 1 38624
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_70_220
timestamp 1646674385
transform 1 0 21344 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_228
timestamp 1646674385
transform 1 0 22080 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1727_
timestamp 1646674385
transform -1 0 21344 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2344_
timestamp 1646674385
transform -1 0 22448 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_232
timestamp 1646674385
transform 1 0 22448 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_238
timestamp 1646674385
transform 1 0 23000 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1646674385
transform 1 0 23920 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1701_
timestamp 1646674385
transform 1 0 23092 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_70_253
timestamp 1646674385
transform 1 0 24380 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_261
timestamp 1646674385
transform 1 0 25116 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_267
timestamp 1646674385
transform 1 0 25668 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1646674385
transform 1 0 24288 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1698_
timestamp 1646674385
transform 1 0 24748 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2126_
timestamp 1646674385
transform 1 0 25760 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_70_273
timestamp 1646674385
transform 1 0 26220 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_284
timestamp 1646674385
transform 1 0 27232 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_288
timestamp 1646674385
transform 1 0 27600 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2131_
timestamp 1646674385
transform 1 0 27692 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2147_
timestamp 1646674385
transform 1 0 26588 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2082__A
timestamp 1646674385
transform 1 0 28888 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_298
timestamp 1646674385
transform 1 0 28520 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1646674385
transform 1 0 29072 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1646674385
transform 1 0 29440 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1681_
timestamp 1646674385
transform 1 0 29532 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_313
timestamp 1646674385
transform 1 0 29900 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_320
timestamp 1646674385
transform 1 0 30544 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_329
timestamp 1646674385
transform 1 0 31372 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1646674385
transform -1 0 32016 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2134_
timestamp 1646674385
transform -1 0 30544 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2573_
timestamp 1646674385
transform -1 0 31372 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_19
timestamp 1646674385
transform 1 0 2852 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1646674385
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2813_
timestamp 1646674385
transform 1 0 1380 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__B2
timestamp 1646674385
transform -1 0 4600 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_32
timestamp 1646674385
transform 1 0 4048 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_38
timestamp 1646674385
transform 1 0 4600 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1500_
timestamp 1646674385
transform -1 0 4048 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_71_52
timestamp 1646674385
transform 1 0 5888 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1646674385
transform 1 0 6256 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_2  _1970_
timestamp 1646674385
transform 1 0 4968 0 -1 39712
box -38 -48 958 592
use sky130_fd_sc_hd__o211ai_4  _1975_
timestamp 1646674385
transform 1 0 6348 0 -1 39712
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_71_74
timestamp 1646674385
transform 1 0 7912 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2641_
timestamp 1646674385
transform 1 0 8280 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_71_103
timestamp 1646674385
transform 1 0 10580 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_94
timestamp 1646674385
transform 1 0 9752 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2293_
timestamp 1646674385
transform -1 0 10580 0 -1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1646674385
transform 1 0 11316 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_113
timestamp 1646674385
transform 1 0 11500 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1646674385
transform 1 0 11408 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1764_
timestamp 1646674385
transform 1 0 11776 0 -1 39712
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_71_126
timestamp 1646674385
transform 1 0 12696 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_140
timestamp 1646674385
transform 1 0 13984 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1765_
timestamp 1646674385
transform -1 0 13984 0 -1 39712
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2071_
timestamp 1646674385
transform 1 0 14352 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_147
timestamp 1646674385
transform 1 0 14628 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_155
timestamp 1646674385
transform 1 0 15364 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1646674385
transform 1 0 15916 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2063_
timestamp 1646674385
transform -1 0 15916 0 -1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1646674385
transform 1 0 16468 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_169
timestamp 1646674385
transform 1 0 16652 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_173
timestamp 1646674385
transform 1 0 17020 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1646674385
transform 1 0 16560 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2675_
timestamp 1646674385
transform -1 0 18584 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_71_190
timestamp 1646674385
transform 1 0 18584 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_198
timestamp 1646674385
transform 1 0 19320 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2680_
timestamp 1646674385
transform -1 0 20884 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_71_215
timestamp 1646674385
transform 1 0 20884 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1646674385
transform 1 0 21620 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_225
timestamp 1646674385
transform 1 0 21804 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1646674385
transform 1 0 21712 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _2373_
timestamp 1646674385
transform 1 0 22080 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_236
timestamp 1646674385
transform 1 0 22816 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_246
timestamp 1646674385
transform 1 0 23736 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_250
timestamp 1646674385
transform 1 0 24104 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1687_
timestamp 1646674385
transform -1 0 23736 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_254
timestamp 1646674385
transform 1 0 24472 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_268
timestamp 1646674385
transform 1 0 25760 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1695_
timestamp 1646674385
transform -1 0 25760 0 -1 39712
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2354_
timestamp 1646674385
transform 1 0 24196 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_276
timestamp 1646674385
transform 1 0 26496 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_290
timestamp 1646674385
transform 1 0 27784 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1646674385
transform 1 0 26864 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1690_
timestamp 1646674385
transform -1 0 26496 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2148_
timestamp 1646674385
transform -1 0 27784 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_71_294
timestamp 1646674385
transform 1 0 28152 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_304
timestamp 1646674385
transform 1 0 29072 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1685_
timestamp 1646674385
transform 1 0 28244 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2129_
timestamp 1646674385
transform -1 0 29900 0 -1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2126__A
timestamp 1646674385
transform 1 0 30268 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2126__B
timestamp 1646674385
transform -1 0 31004 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_313
timestamp 1646674385
transform 1 0 29900 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_319
timestamp 1646674385
transform 1 0 30452 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_325
timestamp 1646674385
transform 1 0 31004 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1646674385
transform -1 0 32016 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_15
timestamp 1646674385
transform 1 0 2484 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_72_3
timestamp 1646674385
transform 1 0 1380 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_13
timestamp 1646674385
transform 1 0 2300 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1646674385
transform 1 0 1380 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1646674385
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1646674385
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1495_
timestamp 1646674385
transform -1 0 2484 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2810_
timestamp 1646674385
transform 1 0 2668 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1646674385
transform 1 0 1748 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1646674385
transform 1 0 3312 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_38
timestamp 1646674385
transform 1 0 4600 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_33
timestamp 1646674385
transform 1 0 4140 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1646674385
transform 1 0 3680 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1498_
timestamp 1646674385
transform 1 0 3772 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1887_
timestamp 1646674385
transform -1 0 3312 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1971_
timestamp 1646674385
transform -1 0 5244 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2582_
timestamp 1646674385
transform -1 0 6072 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1968_
timestamp 1646674385
transform -1 0 5888 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_52
timestamp 1646674385
transform 1 0 5888 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_45
timestamp 1646674385
transform 1 0 5244 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_44
timestamp 1646674385
transform 1 0 5152 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1497_
timestamp 1646674385
transform -1 0 6808 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1646674385
transform 1 0 6256 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_57
timestamp 1646674385
transform 1 0 6348 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_62
timestamp 1646674385
transform 1 0 6808 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_54
timestamp 1646674385
transform 1 0 6072 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2642_
timestamp 1646674385
transform 1 0 6440 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_72_69
timestamp 1646674385
transform 1 0 7452 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_80
timestamp 1646674385
transform 1 0 8464 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_74
timestamp 1646674385
transform 1 0 7912 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1795_
timestamp 1646674385
transform -1 0 9108 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1967_
timestamp 1646674385
transform 1 0 7176 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2314_
timestamp 1646674385
transform 1 0 8188 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_85
timestamp 1646674385
transform 1 0 8924 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_97
timestamp 1646674385
transform 1 0 10028 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_87
timestamp 1646674385
transform 1 0 9108 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_94
timestamp 1646674385
transform 1 0 9752 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1646674385
transform 1 0 8832 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _2290_
timestamp 1646674385
transform -1 0 10856 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2291_
timestamp 1646674385
transform -1 0 9752 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2317_
timestamp 1646674385
transform 1 0 9200 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _2318_
timestamp 1646674385
transform -1 0 10856 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2289_
timestamp 1646674385
transform -1 0 11500 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2275_
timestamp 1646674385
transform -1 0 11776 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1646674385
transform 1 0 11408 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_106
timestamp 1646674385
transform 1 0 10856 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_113
timestamp 1646674385
transform 1 0 11500 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_106
timestamp 1646674385
transform 1 0 10856 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1761_
timestamp 1646674385
transform -1 0 13064 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_73_120
timestamp 1646674385
transform 1 0 12144 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_116
timestamp 1646674385
transform 1 0 11776 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1746_
timestamp 1646674385
transform -1 0 12788 0 1 39712
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_72_127
timestamp 1646674385
transform 1 0 12788 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_135
timestamp 1646674385
transform 1 0 13524 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1646674385
transform 1 0 13892 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_130
timestamp 1646674385
transform 1 0 13064 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1646674385
transform 1 0 13984 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1730_
timestamp 1646674385
transform 1 0 13156 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1762_
timestamp 1646674385
transform -1 0 14904 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2659_
timestamp 1646674385
transform 1 0 13432 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_72_150
timestamp 1646674385
transform 1 0 14904 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_158
timestamp 1646674385
transform 1 0 15640 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_164
timestamp 1646674385
transform 1 0 16192 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_150
timestamp 1646674385
transform 1 0 14904 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_158
timestamp 1646674385
transform 1 0 15640 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1646674385
transform 1 0 16192 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1990_
timestamp 1646674385
transform -1 0 16192 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2051_
timestamp 1646674385
transform -1 0 16192 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_72_170
timestamp 1646674385
transform 1 0 16744 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_187
timestamp 1646674385
transform 1 0 18308 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 1646674385
transform 1 0 16652 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_180
timestamp 1646674385
transform 1 0 17664 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1646674385
transform 1 0 16560 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1729_
timestamp 1646674385
transform -1 0 18952 0 -1 40800
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1737_
timestamp 1646674385
transform 1 0 16836 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2674_
timestamp 1646674385
transform -1 0 18308 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1646674385
transform 1 0 19044 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_197
timestamp 1646674385
transform 1 0 19228 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_194
timestamp 1646674385
transform 1 0 18952 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1646674385
transform 1 0 19136 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2681_
timestamp 1646674385
transform 1 0 19320 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_prog_clk
timestamp 1646674385
transform 1 0 19596 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1687__A
timestamp 1646674385
transform -1 0 21344 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_221
timestamp 1646674385
transform 1 0 21436 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_214
timestamp 1646674385
transform 1 0 20792 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_220
timestamp 1646674385
transform 1 0 21344 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1646674385
transform 1 0 21712 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2372_
timestamp 1646674385
transform 1 0 21804 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _2374_
timestamp 1646674385
transform 1 0 21804 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_234
timestamp 1646674385
transform 1 0 22632 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_238
timestamp 1646674385
transform 1 0 23000 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1646674385
transform 1 0 23920 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_233
timestamp 1646674385
transform 1 0 22540 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_239
timestamp 1646674385
transform 1 0 23092 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1702_
timestamp 1646674385
transform -1 0 23920 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2694_
timestamp 1646674385
transform -1 0 24656 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_72_256
timestamp 1646674385
transform 1 0 24656 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_256
timestamp 1646674385
transform 1 0 24656 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_269
timestamp 1646674385
transform 1 0 25852 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1646674385
transform 1 0 24288 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1697_
timestamp 1646674385
transform 1 0 25024 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2346_
timestamp 1646674385
transform -1 0 24656 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2698_
timestamp 1646674385
transform 1 0 25024 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_72_276
timestamp 1646674385
transform 1 0 26496 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1646674385
transform 1 0 26496 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_288
timestamp 1646674385
transform 1 0 27600 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1646674385
transform 1 0 26864 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1686_
timestamp 1646674385
transform -1 0 27968 0 1 39712
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _2130_
timestamp 1646674385
transform 1 0 26956 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2363_
timestamp 1646674385
transform 1 0 26220 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2082_
timestamp 1646674385
transform -1 0 28612 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_299
timestamp 1646674385
transform 1 0 28612 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_292
timestamp 1646674385
transform 1 0 27968 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1683_
timestamp 1646674385
transform 1 0 29532 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1646674385
transform 1 0 29440 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_308
timestamp 1646674385
transform 1 0 29440 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_304
timestamp 1646674385
transform 1 0 29072 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1646674385
transform 1 0 29348 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2706_
timestamp 1646674385
transform 1 0 29532 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1678_
timestamp 1646674385
transform 1 0 28152 0 -1 40800
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_72_318
timestamp 1646674385
transform 1 0 30360 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_329
timestamp 1646674385
transform 1 0 31372 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_325
timestamp 1646674385
transform 1 0 31004 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1646674385
transform -1 0 32016 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1646674385
transform -1 0 32016 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output52
timestamp 1646674385
transform -1 0 31372 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__B2
timestamp 1646674385
transform -1 0 2668 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2319__A2
timestamp 1646674385
transform -1 0 2116 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_prog_clk_A
timestamp 1646674385
transform -1 0 1564 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_11
timestamp 1646674385
transform 1 0 2116 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_17
timestamp 1646674385
transform 1 0 2668 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_5
timestamp 1646674385
transform 1 0 1564 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1646674385
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1973__A2
timestamp 1646674385
transform -1 0 3312 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_21
timestamp 1646674385
transform 1 0 3036 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_24
timestamp 1646674385
transform 1 0 3312 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_29
timestamp 1646674385
transform 1 0 3772 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_33
timestamp 1646674385
transform 1 0 4140 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1646674385
transform 1 0 3680 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1886_
timestamp 1646674385
transform -1 0 4140 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1973_
timestamp 1646674385
transform -1 0 5244 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2183__A2
timestamp 1646674385
transform -1 0 6716 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_45
timestamp 1646674385
transform 1 0 5244 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_52
timestamp 1646674385
transform 1 0 5888 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_58
timestamp 1646674385
transform 1 0 6440 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_61
timestamp 1646674385
transform 1 0 6716 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1889_
timestamp 1646674385
transform -1 0 5888 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1791__A
timestamp 1646674385
transform 1 0 7636 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2182__A2
timestamp 1646674385
transform -1 0 7268 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_67
timestamp 1646674385
transform 1 0 7268 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_73
timestamp 1646674385
transform 1 0 7820 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1646674385
transform 1 0 8464 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2296_
timestamp 1646674385
transform 1 0 8188 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_95
timestamp 1646674385
transform 1 0 9844 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1646674385
transform 1 0 8832 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1791_
timestamp 1646674385
transform 1 0 8924 0 1 40800
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_1  _2319_
timestamp 1646674385
transform -1 0 10948 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_107
timestamp 1646674385
transform 1 0 10948 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2661_
timestamp 1646674385
transform 1 0 11684 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_74_131
timestamp 1646674385
transform 1 0 13156 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1646674385
transform 1 0 13892 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1646674385
transform 1 0 13984 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2660_
timestamp 1646674385
transform -1 0 15548 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_74_157
timestamp 1646674385
transform 1 0 15548 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _2072_
timestamp 1646674385
transform 1 0 15916 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_74_168
timestamp 1646674385
transform 1 0 16560 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_177
timestamp 1646674385
transform 1 0 17388 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_186
timestamp 1646674385
transform 1 0 18216 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2049_
timestamp 1646674385
transform -1 0 17388 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2054_
timestamp 1646674385
transform -1 0 18216 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1707__A
timestamp 1646674385
transform 1 0 18584 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1646674385
transform 1 0 18768 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_206
timestamp 1646674385
transform 1 0 20056 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1646674385
transform 1 0 19136 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1725_
timestamp 1646674385
transform -1 0 20056 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_74_224
timestamp 1646674385
transform 1 0 21712 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1721_
timestamp 1646674385
transform 1 0 20792 0 1 40800
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _2371_
timestamp 1646674385
transform -1 0 22724 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_74_235
timestamp 1646674385
transform 1 0 22724 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_244
timestamp 1646674385
transform 1 0 23552 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2361_
timestamp 1646674385
transform 1 0 23092 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_74_263
timestamp 1646674385
transform 1 0 25300 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_267
timestamp 1646674385
transform 1 0 25668 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1646674385
transform 1 0 24288 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1694_
timestamp 1646674385
transform -1 0 26588 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1696_
timestamp 1646674385
transform 1 0 24380 0 1 40800
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_74_277
timestamp 1646674385
transform 1 0 26588 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_prog_clk
timestamp 1646674385
transform 1 0 26956 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1646674385
transform 1 0 28796 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1646674385
transform 1 0 29348 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_309
timestamp 1646674385
transform 1 0 29532 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1646674385
transform 1 0 29440 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2705_
timestamp 1646674385
transform 1 0 29624 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_74_326
timestamp 1646674385
transform 1 0 31096 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_332
timestamp 1646674385
transform 1 0 31648 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1646674385
transform -1 0 32016 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2492__B2
timestamp 1646674385
transform -1 0 2760 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1646674385
transform -1 0 2208 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1646674385
transform -1 0 1656 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_12
timestamp 1646674385
transform 1 0 2208 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_18
timestamp 1646674385
transform 1 0 2760 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_3
timestamp 1646674385
transform 1 0 1380 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_6
timestamp 1646674385
transform 1 0 1656 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1646674385
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2318__A2
timestamp 1646674385
transform 1 0 3128 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_24
timestamp 1646674385
transform 1 0 3312 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2811_
timestamp 1646674385
transform 1 0 3680 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2258__C
timestamp 1646674385
transform -1 0 5888 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_44
timestamp 1646674385
transform 1 0 5152 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_52
timestamp 1646674385
transform 1 0 5888 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1646674385
transform 1 0 6256 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2643_
timestamp 1646674385
transform -1 0 7820 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_73
timestamp 1646674385
transform 1 0 7820 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1792_
timestamp 1646674385
transform -1 0 9016 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_75_86
timestamp 1646674385
transform 1 0 9016 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_97
timestamp 1646674385
transform 1 0 10028 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2299_
timestamp 1646674385
transform 1 0 9384 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2307_
timestamp 1646674385
transform -1 0 10856 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_75_106
timestamp 1646674385
transform 1 0 10856 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_113
timestamp 1646674385
transform 1 0 11500 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_120
timestamp 1646674385
transform 1 0 12144 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1646674385
transform 1 0 11408 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1759_
timestamp 1646674385
transform -1 0 13432 0 -1 41888
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2070_
timestamp 1646674385
transform -1 0 12144 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_134
timestamp 1646674385
transform 1 0 13432 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_prog_clk
timestamp 1646674385
transform 1 0 14168 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_75_162
timestamp 1646674385
transform 1 0 16008 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2275__A
timestamp 1646674385
transform -1 0 18032 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_178
timestamp 1646674385
transform 1 0 17480 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_184
timestamp 1646674385
transform 1 0 18032 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1646674385
transform 1 0 16560 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2073_
timestamp 1646674385
transform 1 0 16652 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_75_198
timestamp 1646674385
transform 1 0 19320 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1707_
timestamp 1646674385
transform -1 0 19320 0 -1 41888
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1722_
timestamp 1646674385
transform -1 0 20608 0 -1 41888
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_75_212
timestamp 1646674385
transform 1 0 20608 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_219
timestamp 1646674385
transform 1 0 21252 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1646674385
transform 1 0 21620 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1646674385
transform 1 0 21712 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1989_
timestamp 1646674385
transform 1 0 20976 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2351_
timestamp 1646674385
transform 1 0 21804 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_75_230
timestamp 1646674385
transform 1 0 22264 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_243
timestamp 1646674385
transform 1 0 23460 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_250
timestamp 1646674385
transform 1 0 24104 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2345_
timestamp 1646674385
transform 1 0 23828 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2368_
timestamp 1646674385
transform -1 0 23460 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1697__B1
timestamp 1646674385
transform -1 0 24656 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_256
timestamp 1646674385
transform 1 0 24656 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2699_
timestamp 1646674385
transform 1 0 25024 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1646674385
transform 1 0 26496 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_281
timestamp 1646674385
transform 1 0 26956 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_285
timestamp 1646674385
transform 1 0 27324 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_291
timestamp 1646674385
transform 1 0 27876 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1646674385
transform 1 0 26864 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2145_
timestamp 1646674385
transform 1 0 27048 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_295
timestamp 1646674385
transform 1 0 28244 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2125_
timestamp 1646674385
transform -1 0 28244 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2704_
timestamp 1646674385
transform 1 0 28612 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2338__A2
timestamp 1646674385
transform -1 0 30636 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2338__B2
timestamp 1646674385
transform 1 0 31004 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_315
timestamp 1646674385
transform 1 0 30084 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_321
timestamp 1646674385
transform 1 0 30636 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_327
timestamp 1646674385
transform 1 0 31188 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1646674385
transform -1 0 32016 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_13
timestamp 1646674385
transform 1 0 2300 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1646674385
transform 1 0 1380 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1646674385
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1646674385
transform 1 0 1748 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1971__A2
timestamp 1646674385
transform -1 0 4508 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2318__A1
timestamp 1646674385
transform -1 0 3956 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2571__A
timestamp 1646674385
transform -1 0 3312 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_21
timestamp 1646674385
transform 1 0 3036 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1646674385
transform 1 0 3312 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_31
timestamp 1646674385
transform 1 0 3956 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_37
timestamp 1646674385
transform 1 0 4508 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_41
timestamp 1646674385
transform 1 0 4876 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1646674385
transform 1 0 3680 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2278__B
timestamp 1646674385
transform -1 0 6256 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2279__A2
timestamp 1646674385
transform -1 0 5704 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2280__A2
timestamp 1646674385
transform 1 0 4968 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_44
timestamp 1646674385
transform 1 0 5152 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_50
timestamp 1646674385
transform 1 0 5704 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_56
timestamp 1646674385
transform 1 0 6256 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2297_
timestamp 1646674385
transform 1 0 6624 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_63
timestamp 1646674385
transform 1 0 6900 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_76
timestamp 1646674385
transform 1 0 8096 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1788_
timestamp 1646674385
transform -1 0 8096 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_94
timestamp 1646674385
transform 1 0 9752 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1646674385
transform 1 0 8832 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _2300_
timestamp 1646674385
transform 1 0 8924 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2313_
timestamp 1646674385
transform 1 0 10120 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_107
timestamp 1646674385
transform 1 0 10948 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_111
timestamp 1646674385
transform 1 0 11316 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_116
timestamp 1646674385
transform 1 0 11776 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1750_
timestamp 1646674385
transform 1 0 12144 0 1 41888
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1767_
timestamp 1646674385
transform 1 0 11408 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1750__A
timestamp 1646674385
transform -1 0 13616 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_130
timestamp 1646674385
transform 1 0 13064 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1646674385
transform 1 0 13616 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1646674385
transform 1 0 13984 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1763_
timestamp 1646674385
transform -1 0 14904 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2257__B2
timestamp 1646674385
transform 1 0 15272 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_150
timestamp 1646674385
transform 1 0 14904 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_156
timestamp 1646674385
transform 1 0 15456 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2069_
timestamp 1646674385
transform -1 0 16652 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_169
timestamp 1646674385
transform 1 0 16652 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2673_
timestamp 1646674385
transform -1 0 18492 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1646674385
transform 1 0 18492 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1646674385
transform 1 0 19044 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_200
timestamp 1646674385
transform 1 0 19504 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1646674385
transform 1 0 19136 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1966_
timestamp 1646674385
transform 1 0 19228 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2683_
timestamp 1646674385
transform 1 0 19872 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_220
timestamp 1646674385
transform 1 0 21344 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2353_
timestamp 1646674385
transform 1 0 21712 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_233
timestamp 1646674385
transform 1 0 22540 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_244
timestamp 1646674385
transform 1 0 23552 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2366_
timestamp 1646674385
transform 1 0 22908 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_76_269
timestamp 1646674385
transform 1 0 25852 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1646674385
transform 1 0 24288 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2693_
timestamp 1646674385
transform 1 0 24380 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_282
timestamp 1646674385
transform 1 0 27048 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_289
timestamp 1646674385
transform 1 0 27692 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1693_
timestamp 1646674385
transform 1 0 26220 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2146_
timestamp 1646674385
transform 1 0 27416 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_296
timestamp 1646674385
transform 1 0 28336 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_300
timestamp 1646674385
transform 1 0 28704 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1646674385
transform 1 0 29072 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1646674385
transform 1 0 29440 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1684_
timestamp 1646674385
transform 1 0 29532 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2123_
timestamp 1646674385
transform -1 0 29072 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2128_
timestamp 1646674385
transform -1 0 28336 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_318
timestamp 1646674385
transform 1 0 30360 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_329
timestamp 1646674385
transform 1 0 31372 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1646674385
transform -1 0 32016 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output30
timestamp 1646674385
transform -1 0 31372 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1646674385
transform -1 0 1564 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1646674385
transform -1 0 2116 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1646674385
transform -1 0 2668 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_11
timestamp 1646674385
transform 1 0 2116 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_17
timestamp 1646674385
transform 1 0 2668 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_5
timestamp 1646674385
transform 1 0 1564 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1646674385
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2283__A2
timestamp 1646674385
transform -1 0 4600 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_prog_clk_A
timestamp 1646674385
transform -1 0 4048 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1646674385
transform -1 0 3220 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_23
timestamp 1646674385
transform 1 0 3220 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_29
timestamp 1646674385
transform 1 0 3772 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_32
timestamp 1646674385
transform 1 0 4048 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_38
timestamp 1646674385
transform 1 0 4600 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1782__A
timestamp 1646674385
transform -1 0 6900 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2281__A2
timestamp 1646674385
transform -1 0 5336 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2282__A2
timestamp 1646674385
transform 1 0 5704 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_46
timestamp 1646674385
transform 1 0 5336 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_52
timestamp 1646674385
transform 1 0 5888 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_57
timestamp 1646674385
transform 1 0 6348 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1646674385
transform 1 0 6256 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_63
timestamp 1646674385
transform 1 0 6900 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_70
timestamp 1646674385
transform 1 0 7544 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1782_
timestamp 1646674385
transform 1 0 7912 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2294_
timestamp 1646674385
transform 1 0 7268 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_84
timestamp 1646674385
transform 1 0 8832 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_97
timestamp 1646674385
transform 1 0 10028 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2306_
timestamp 1646674385
transform 1 0 9200 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2312_
timestamp 1646674385
transform 1 0 10396 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_77_108
timestamp 1646674385
transform 1 0 11040 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1646674385
transform 1 0 11408 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2653_
timestamp 1646674385
transform 1 0 11500 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_129
timestamp 1646674385
transform 1 0 12972 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_143
timestamp 1646674385
transform 1 0 14260 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1757_
timestamp 1646674385
transform 1 0 13340 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_77_156
timestamp 1646674385
transform 1 0 15456 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_163
timestamp 1646674385
transform 1 0 16100 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1760_
timestamp 1646674385
transform 1 0 14628 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2052_
timestamp 1646674385
transform 1 0 15824 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1646674385
transform 1 0 16468 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_169
timestamp 1646674385
transform 1 0 16652 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_181
timestamp 1646674385
transform 1 0 17756 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1646674385
transform 1 0 16560 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1740_
timestamp 1646674385
transform 1 0 16928 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_77_189
timestamp 1646674385
transform 1 0 18492 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_206
timestamp 1646674385
transform 1 0 20056 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2682_
timestamp 1646674385
transform 1 0 18584 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2327__B2
timestamp 1646674385
transform 1 0 21804 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_220
timestamp 1646674385
transform 1 0 21344 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_227
timestamp 1646674385
transform 1 0 21988 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1646674385
transform 1 0 21712 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1724_
timestamp 1646674385
transform 1 0 20424 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_77_240
timestamp 1646674385
transform 1 0 23184 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1706_
timestamp 1646674385
transform 1 0 23552 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1709_
timestamp 1646674385
transform -1 0 23184 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_77_253
timestamp 1646674385
transform 1 0 24380 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_269
timestamp 1646674385
transform 1 0 25852 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1688_
timestamp 1646674385
transform 1 0 24932 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2147__B
timestamp 1646674385
transform -1 0 27140 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_276
timestamp 1646674385
transform 1 0 26496 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_283
timestamp 1646674385
transform 1 0 27140 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1646674385
transform 1 0 26864 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1689_
timestamp 1646674385
transform 1 0 27508 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2364_
timestamp 1646674385
transform 1 0 26220 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_296
timestamp 1646674385
transform 1 0 28336 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_303
timestamp 1646674385
transform 1 0 28980 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_310
timestamp 1646674385
transform 1 0 29624 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2127_
timestamp 1646674385
transform 1 0 28704 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2365_
timestamp 1646674385
transform 1 0 29348 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2389__C
timestamp 1646674385
transform 1 0 29992 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2572__A
timestamp 1646674385
transform 1 0 30912 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_316
timestamp 1646674385
transform 1 0 30176 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_77_326
timestamp 1646674385
transform 1 0 31096 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_332
timestamp 1646674385
transform 1 0 31648 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1646674385
transform -1 0 32016 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1646674385
transform -1 0 1564 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1646674385
transform -1 0 2116 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1646674385
transform -1 0 2668 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_11
timestamp 1646674385
transform 1 0 2116 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_17
timestamp 1646674385
transform 1 0 2668 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_5
timestamp 1646674385
transform 1 0 1564 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1646674385
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_prog_clk_A
timestamp 1646674385
transform 1 0 4876 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1646674385
transform -1 0 3220 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1646674385
transform 1 0 3220 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1646674385
transform 1 0 3588 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1646674385
transform 1 0 3772 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1646674385
transform 1 0 3680 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2307__A
timestamp 1646674385
transform -1 0 5612 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_43
timestamp 1646674385
transform 1 0 5060 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_49
timestamp 1646674385
transform 1 0 5612 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2644_
timestamp 1646674385
transform 1 0 5980 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_78_69
timestamp 1646674385
transform 1 0 7452 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1646674385
transform 1 0 8464 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2292_
timestamp 1646674385
transform 1 0 8188 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_100
timestamp 1646674385
transform 1 0 10304 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_85
timestamp 1646674385
transform 1 0 8924 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_89
timestamp 1646674385
transform 1 0 9292 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1646674385
transform 1 0 8832 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1774_
timestamp 1646674385
transform 1 0 9384 0 1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1775_
timestamp 1646674385
transform 1 0 10672 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2257__A2
timestamp 1646674385
transform -1 0 12052 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_113
timestamp 1646674385
transform 1 0 11500 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_119
timestamp 1646674385
transform 1 0 12052 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1756_
timestamp 1646674385
transform 1 0 12420 0 1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1646674385
transform 1 0 13340 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1646674385
transform 1 0 13892 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1646674385
transform 1 0 13984 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2662_
timestamp 1646674385
transform -1 0 15548 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_78_157
timestamp 1646674385
transform 1 0 15548 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1739_
timestamp 1646674385
transform 1 0 16284 0 1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_78_175
timestamp 1646674385
transform 1 0 17204 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_181
timestamp 1646674385
transform 1 0 17756 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1741_
timestamp 1646674385
transform -1 0 18768 0 1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_78_192
timestamp 1646674385
transform 1 0 18768 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_197
timestamp 1646674385
transform 1 0 19228 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_202
timestamp 1646674385
transform 1 0 19688 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1646674385
transform 1 0 19136 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1716_
timestamp 1646674385
transform -1 0 20976 0 1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1733_
timestamp 1646674385
transform -1 0 19688 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_216
timestamp 1646674385
transform 1 0 20976 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_224
timestamp 1646674385
transform 1 0 21712 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1708_
timestamp 1646674385
transform 1 0 21344 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2328__C
timestamp 1646674385
transform -1 0 23920 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_242
timestamp 1646674385
transform 1 0 23368 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1646674385
transform 1 0 23920 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1704_
timestamp 1646674385
transform 1 0 22448 0 1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_78_269
timestamp 1646674385
transform 1 0 25852 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1646674385
transform 1 0 24288 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2692_
timestamp 1646674385
transform 1 0 24380 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_284
timestamp 1646674385
transform 1 0 27232 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1691_
timestamp 1646674385
transform 1 0 26404 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2703_
timestamp 1646674385
transform 1 0 27600 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1646674385
transform -1 0 29716 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1646674385
transform 1 0 29072 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_311
timestamp 1646674385
transform 1 0 29716 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1646674385
transform 1 0 29440 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2573__A
timestamp 1646674385
transform 1 0 30544 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_319
timestamp 1646674385
transform 1 0 30452 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_322
timestamp 1646674385
transform 1 0 30728 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_329
timestamp 1646674385
transform 1 0 31372 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1646674385
transform -1 0 32016 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2574_
timestamp 1646674385
transform -1 0 31372 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1646674385
transform 1 0 1748 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1646674385
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1646674385
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1646674385
transform 1 0 1380 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_7
timestamp 1646674385
transform 1 0 1748 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1646674385
transform 1 0 1380 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1646674385
transform -1 0 1748 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1646674385
transform -1 0 2300 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_13
timestamp 1646674385
transform 1 0 2300 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_13
timestamp 1646674385
transform 1 0 2300 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_25
timestamp 1646674385
transform 1 0 3404 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_37
timestamp 1646674385
transform 1 0 4508 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_25
timestamp 1646674385
transform 1 0 3404 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1646674385
transform 1 0 3772 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_41
timestamp 1646674385
transform 1 0 4876 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1646674385
transform 1 0 3680 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2493__C
timestamp 1646674385
transform -1 0 5888 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_49
timestamp 1646674385
transform 1 0 5612 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1646674385
transform 1 0 5888 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_57
timestamp 1646674385
transform 1 0 6348 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_61
timestamp 1646674385
transform 1 0 6716 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_49
timestamp 1646674385
transform 1 0 5612 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1646674385
transform 1 0 6256 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1787_
timestamp 1646674385
transform -1 0 7636 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2645_
timestamp 1646674385
transform 1 0 5796 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_79_71
timestamp 1646674385
transform 1 0 7636 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_67
timestamp 1646674385
transform 1 0 7268 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1646674385
transform 1 0 8464 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1784_
timestamp 1646674385
transform -1 0 8924 0 -1 44064
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _2305_
timestamp 1646674385
transform 1 0 7820 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1646674385
transform 1 0 8832 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_90
timestamp 1646674385
transform 1 0 9384 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_85
timestamp 1646674385
transform 1 0 8924 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_85
timestamp 1646674385
transform 1 0 8924 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1774__A
timestamp 1646674385
transform -1 0 9384 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _2308_
timestamp 1646674385
transform -1 0 10948 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_94
timestamp 1646674385
transform 1 0 9752 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_99
timestamp 1646674385
transform 1 0 10212 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_103
timestamp 1646674385
transform 1 0 10580 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_prog_clk
timestamp 1646674385
transform 1 0 9844 0 1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1772_
timestamp 1646674385
transform 1 0 9292 0 -1 44064
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_79_107
timestamp 1646674385
transform 1 0 10948 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1646674385
transform 1 0 11316 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1646674385
transform 1 0 11500 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_118
timestamp 1646674385
transform 1 0 11960 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_115
timestamp 1646674385
transform 1 0 11684 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1646674385
transform 1 0 11408 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2053_
timestamp 1646674385
transform -1 0 11960 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2652_
timestamp 1646674385
transform 1 0 12052 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2663_
timestamp 1646674385
transform 1 0 12328 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_79_138
timestamp 1646674385
transform 1 0 13800 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1646674385
transform 1 0 13524 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1646674385
transform 1 0 13892 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1646674385
transform 1 0 13984 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1751_
timestamp 1646674385
transform 1 0 14076 0 1 44064
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1758_
timestamp 1646674385
transform -1 0 14996 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_79_151
timestamp 1646674385
transform 1 0 14996 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1646674385
transform 1 0 16192 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_151
timestamp 1646674385
transform 1 0 14996 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_155
timestamp 1646674385
transform 1 0 15364 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_165
timestamp 1646674385
transform 1 0 16284 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2056_
timestamp 1646674385
transform -1 0 16192 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _2062_
timestamp 1646674385
transform 1 0 15456 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2332__A2
timestamp 1646674385
transform -1 0 16836 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_171
timestamp 1646674385
transform 1 0 16836 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_180
timestamp 1646674385
transform 1 0 17664 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_187
timestamp 1646674385
transform 1 0 18308 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1646674385
transform 1 0 16560 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1742_
timestamp 1646674385
transform 1 0 16836 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2064_
timestamp 1646674385
transform -1 0 18308 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2672_
timestamp 1646674385
transform 1 0 17204 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_79_191
timestamp 1646674385
transform 1 0 18676 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_205
timestamp 1646674385
transform 1 0 19964 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1646674385
transform 1 0 19044 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_200
timestamp 1646674385
transform 1 0 19504 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_206
timestamp 1646674385
transform 1 0 20056 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1646674385
transform 1 0 19136 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1714_
timestamp 1646674385
transform -1 0 21068 0 1 44064
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1738_
timestamp 1646674385
transform 1 0 19044 0 -1 44064
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2065_
timestamp 1646674385
transform 1 0 19228 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_218
timestamp 1646674385
transform 1 0 21160 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_217
timestamp 1646674385
transform 1 0 21068 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_224
timestamp 1646674385
transform 1 0 21712 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1646674385
transform 1 0 21712 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1723_
timestamp 1646674385
transform 1 0 20332 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2347_
timestamp 1646674385
transform 1 0 21436 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2360_
timestamp 1646674385
transform -1 0 22632 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_79_234
timestamp 1646674385
transform 1 0 22632 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_250
timestamp 1646674385
transform 1 0 24104 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_239
timestamp 1646674385
transform 1 0 23092 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_246
timestamp 1646674385
transform 1 0 23736 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1705_
timestamp 1646674385
transform 1 0 23184 0 -1 44064
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2356_
timestamp 1646674385
transform -1 0 23736 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2367_
timestamp 1646674385
transform -1 0 23092 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2362_
timestamp 1646674385
transform -1 0 24748 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2357_
timestamp 1646674385
transform 1 0 24380 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1646674385
transform 1 0 24288 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_256
timestamp 1646674385
transform 1 0 24656 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_257
timestamp 1646674385
transform 1 0 24748 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2333__A3
timestamp 1646674385
transform -1 0 25208 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1692_
timestamp 1646674385
transform 1 0 25668 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_80_262
timestamp 1646674385
transform 1 0 25208 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_263
timestamp 1646674385
transform 1 0 25300 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2329__B1
timestamp 1646674385
transform -1 0 25300 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2700_
timestamp 1646674385
transform -1 0 27048 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2604__CLK
timestamp 1646674385
transform -1 0 27600 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_276
timestamp 1646674385
transform 1 0 26496 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_281
timestamp 1646674385
transform 1 0 26956 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_285
timestamp 1646674385
transform 1 0 27324 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_282
timestamp 1646674385
transform 1 0 27048 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_288
timestamp 1646674385
transform 1 0 27600 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1646674385
transform 1 0 26864 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2702_
timestamp 1646674385
transform 1 0 27416 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_80_300
timestamp 1646674385
transform 1 0 28704 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_294
timestamp 1646674385
transform 1 0 28152 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_prog_clk_A
timestamp 1646674385
transform 1 0 28520 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2606__CLK
timestamp 1646674385
transform -1 0 28152 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1646674385
transform 1 0 29440 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_309
timestamp 1646674385
transform 1 0 29532 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_309
timestamp 1646674385
transform 1 0 29532 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_306
timestamp 1646674385
transform 1 0 29256 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_302
timestamp 1646674385
transform 1 0 28888 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_prog_clk_A
timestamp 1646674385
transform 1 0 29348 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_317
timestamp 1646674385
transform 1 0 30268 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_79_317
timestamp 1646674385
transform 1 0 30268 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1646674385
transform 1 0 30360 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output42
timestamp 1646674385
transform -1 0 31372 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_322
timestamp 1646674385
transform 1 0 30728 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_326
timestamp 1646674385
transform 1 0 31096 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_320
timestamp 1646674385
transform 1 0 30544 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output37_A
timestamp 1646674385
transform -1 0 30728 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2574__A
timestamp 1646674385
transform 1 0 30912 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1646674385
transform -1 0 32016 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1646674385
transform -1 0 32016 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_329
timestamp 1646674385
transform 1 0 31372 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_332
timestamp 1646674385
transform 1 0 31648 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1646674385
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1646674385
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1646674385
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1646674385
transform 1 0 3588 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1646674385
transform 1 0 4692 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1646674385
transform 1 0 5796 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1646674385
transform 1 0 6164 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_57
timestamp 1646674385
transform 1 0 6348 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1646674385
transform 1 0 6256 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_65
timestamp 1646674385
transform 1 0 7084 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_75
timestamp 1646674385
transform 1 0 8004 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1781_
timestamp 1646674385
transform -1 0 9476 0 -1 45152
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1786_
timestamp 1646674385
transform -1 0 8004 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_81_91
timestamp 1646674385
transform 1 0 9476 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1777_
timestamp 1646674385
transform 1 0 10212 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1646674385
transform 1 0 11040 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_116
timestamp 1646674385
transform 1 0 11776 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_123
timestamp 1646674385
transform 1 0 12420 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1646674385
transform 1 0 11408 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2309_
timestamp 1646674385
transform -1 0 11776 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2311_
timestamp 1646674385
transform 1 0 12144 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_139
timestamp 1646674385
transform 1 0 13892 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1748_
timestamp 1646674385
transform -1 0 13892 0 -1 45152
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _2055_
timestamp 1646674385
transform 1 0 14444 0 -1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_81_152
timestamp 1646674385
transform 1 0 15088 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_163
timestamp 1646674385
transform 1 0 16100 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2061_
timestamp 1646674385
transform 1 0 15456 0 -1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2388__A2
timestamp 1646674385
transform -1 0 16836 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1646674385
transform 1 0 16468 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_171
timestamp 1646674385
transform 1 0 16836 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_184
timestamp 1646674385
transform 1 0 18032 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1646674385
transform 1 0 16560 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1743_
timestamp 1646674385
transform 1 0 17204 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1646674385
transform 1 0 18676 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_198
timestamp 1646674385
transform 1 0 19320 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_202
timestamp 1646674385
transform 1 0 19688 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_206
timestamp 1646674385
transform 1 0 20056 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2066_
timestamp 1646674385
transform -1 0 18676 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2067_
timestamp 1646674385
transform 1 0 19044 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2348_
timestamp 1646674385
transform 1 0 19780 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1646674385
transform 1 0 21344 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1646674385
transform 1 0 21712 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1713_
timestamp 1646674385
transform -1 0 21344 0 -1 45152
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1720_
timestamp 1646674385
transform 1 0 21804 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_81_234
timestamp 1646674385
transform 1 0 22632 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1711_
timestamp 1646674385
transform 1 0 23368 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2335__A
timestamp 1646674385
transform -1 0 25760 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_251
timestamp 1646674385
transform 1 0 24196 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_262
timestamp 1646674385
transform 1 0 25208 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_268
timestamp 1646674385
transform 1 0 25760 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2359_
timestamp 1646674385
transform -1 0 25208 0 -1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2388__B2
timestamp 1646674385
transform -1 0 26312 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_274
timestamp 1646674385
transform 1 0 26312 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1646674385
transform 1 0 26864 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2701_
timestamp 1646674385
transform -1 0 28428 0 -1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_81_297
timestamp 1646674385
transform 1 0 28428 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_309
timestamp 1646674385
transform 1 0 29532 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output40_A
timestamp 1646674385
transform -1 0 31096 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_321
timestamp 1646674385
transform 1 0 30636 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_326
timestamp 1646674385
transform 1 0 31096 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_332
timestamp 1646674385
transform 1 0 31648 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1646674385
transform -1 0 32016 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1646674385
transform -1 0 1564 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_17
timestamp 1646674385
transform 1 0 2668 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_5
timestamp 1646674385
transform 1 0 1564 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1646674385
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_25
timestamp 1646674385
transform 1 0 3404 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1646674385
transform 1 0 3772 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1646674385
transform 1 0 4876 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1646674385
transform 1 0 3680 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_53
timestamp 1646674385
transform 1 0 5980 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_59
timestamp 1646674385
transform 1 0 6532 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2304_
timestamp 1646674385
transform -1 0 6900 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1646674385
transform 1 0 6900 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_76
timestamp 1646674385
transform 1 0 8096 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1785_
timestamp 1646674385
transform 1 0 7268 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_82_100
timestamp 1646674385
transform 1 0 10304 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1646674385
transform 1 0 8924 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_93
timestamp 1646674385
transform 1 0 9660 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1646674385
transform 1 0 8832 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1776_
timestamp 1646674385
transform -1 0 9660 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2301_
timestamp 1646674385
transform 1 0 10028 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2302_
timestamp 1646674385
transform -1 0 10948 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2289__A
timestamp 1646674385
transform -1 0 11500 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_107
timestamp 1646674385
transform 1 0 10948 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_113
timestamp 1646674385
transform 1 0 11500 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_120
timestamp 1646674385
transform 1 0 12144 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1747_
timestamp 1646674385
transform 1 0 12512 0 1 45152
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2060_
timestamp 1646674385
transform -1 0 12144 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_134
timestamp 1646674385
transform 1 0 13432 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1646674385
transform 1 0 13984 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1755_
timestamp 1646674385
transform -1 0 14904 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_82_150
timestamp 1646674385
transform 1 0 14904 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_157
timestamp 1646674385
transform 1 0 15548 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2048_
timestamp 1646674385
transform 1 0 15272 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2068_
timestamp 1646674385
transform 1 0 15916 0 1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_82_168
timestamp 1646674385
transform 1 0 16560 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2671_
timestamp 1646674385
transform 1 0 17296 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_82_192
timestamp 1646674385
transform 1 0 18768 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1646674385
transform 1 0 19136 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2684_
timestamp 1646674385
transform -1 0 20700 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_82_213
timestamp 1646674385
transform 1 0 20700 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_226
timestamp 1646674385
transform 1 0 21896 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1718_
timestamp 1646674385
transform -1 0 21896 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_82_233
timestamp 1646674385
transform 1 0 22540 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1646674385
transform 1 0 23920 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1710_
timestamp 1646674385
transform 1 0 23092 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2350_
timestamp 1646674385
transform 1 0 22264 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_269
timestamp 1646674385
transform 1 0 25852 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1646674385
transform 1 0 24288 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2691_
timestamp 1646674385
transform 1 0 24380 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2605__CLK
timestamp 1646674385
transform 1 0 26220 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_prog_clk_A
timestamp 1646674385
transform 1 0 26772 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_275
timestamp 1646674385
transform 1 0 26404 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1646674385
transform 1 0 26956 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_293
timestamp 1646674385
transform 1 0 28060 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1646674385
transform 1 0 29164 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1646674385
transform 1 0 29532 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1646674385
transform 1 0 29440 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1646674385
transform 1 0 30636 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1646674385
transform -1 0 32016 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_19
timestamp 1646674385
transform 1 0 2852 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_7
timestamp 1646674385
transform 1 0 1748 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1646674385
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1646674385
transform 1 0 1380 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_31
timestamp 1646674385
transform 1 0 3956 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_43
timestamp 1646674385
transform 1 0 5060 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1646674385
transform 1 0 6164 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1646674385
transform 1 0 6256 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2646_
timestamp 1646674385
transform 1 0 6348 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_83_73
timestamp 1646674385
transform 1 0 7820 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_82
timestamp 1646674385
transform 1 0 8648 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2303_
timestamp 1646674385
transform 1 0 8372 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_95
timestamp 1646674385
transform 1 0 9844 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1778_
timestamp 1646674385
transform 1 0 10212 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1780_
timestamp 1646674385
transform 1 0 9016 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_83_108
timestamp 1646674385
transform 1 0 11040 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_116
timestamp 1646674385
transform 1 0 11776 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_124
timestamp 1646674385
transform 1 0 12512 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1646674385
transform 1 0 11408 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1753_
timestamp 1646674385
transform 1 0 12604 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2310_
timestamp 1646674385
transform -1 0 11776 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_134
timestamp 1646674385
transform 1 0 13432 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1752_
timestamp 1646674385
transform 1 0 13800 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_83_147
timestamp 1646674385
transform 1 0 14628 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_160
timestamp 1646674385
transform 1 0 15824 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1749_
timestamp 1646674385
transform 1 0 14996 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_83_178
timestamp 1646674385
transform 1 0 17480 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_185
timestamp 1646674385
transform 1 0 18124 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1646674385
transform 1 0 16560 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1745_
timestamp 1646674385
transform 1 0 16652 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2058_
timestamp 1646674385
transform 1 0 17848 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_83_191
timestamp 1646674385
transform 1 0 18676 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_201
timestamp 1646674385
transform 1 0 19596 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1717_
timestamp 1646674385
transform 1 0 19964 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1719_
timestamp 1646674385
transform -1 0 19596 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2332__B2
timestamp 1646674385
transform -1 0 21344 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_214
timestamp 1646674385
transform 1 0 20792 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_220
timestamp 1646674385
transform 1 0 21344 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1646674385
transform 1 0 21712 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _2352_
timestamp 1646674385
transform 1 0 21804 0 -1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_83_232
timestamp 1646674385
transform 1 0 22448 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_236
timestamp 1646674385
transform 1 0 22816 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2689_
timestamp 1646674385
transform 1 0 22908 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_83_253
timestamp 1646674385
transform 1 0 24380 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2690_
timestamp 1646674385
transform -1 0 26220 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1646674385
transform 1 0 26220 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1646674385
transform 1 0 26772 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_281
timestamp 1646674385
transform 1 0 26956 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1646674385
transform 1 0 26864 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_293
timestamp 1646674385
transform 1 0 28060 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_305
timestamp 1646674385
transform 1 0 29164 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1646674385
transform 1 0 30544 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_83_317
timestamp 1646674385
transform 1 0 30268 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_322
timestamp 1646674385
transform 1 0 30728 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_329
timestamp 1646674385
transform 1 0 31372 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1646674385
transform -1 0 32016 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output31
timestamp 1646674385
transform -1 0 31372 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1646674385
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1646674385
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1646674385
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1646674385
transform 1 0 3588 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1646674385
transform 1 0 3772 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1646674385
transform 1 0 4876 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1646674385
transform 1 0 3680 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1646674385
transform 1 0 5980 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_65
timestamp 1646674385
transform 1 0 7084 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_80
timestamp 1646674385
transform 1 0 8464 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1783_
timestamp 1646674385
transform 1 0 7636 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_84_85
timestamp 1646674385
transform 1 0 8924 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_96
timestamp 1646674385
transform 1 0 9936 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1646674385
transform 1 0 8832 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1779_
timestamp 1646674385
transform 1 0 9108 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2650_
timestamp 1646674385
transform 1 0 10304 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_84_116
timestamp 1646674385
transform 1 0 11776 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2664_
timestamp 1646674385
transform 1 0 12144 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_84_136
timestamp 1646674385
transform 1 0 13616 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_84_141
timestamp 1646674385
transform 1 0 14076 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1646674385
transform 1 0 13984 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2667_
timestamp 1646674385
transform 1 0 14352 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_84_160
timestamp 1646674385
transform 1 0 15824 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2050_
timestamp 1646674385
transform 1 0 16192 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2603__CLK
timestamp 1646674385
transform 1 0 18308 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_167
timestamp 1646674385
transform 1 0 16468 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_173
timestamp 1646674385
transform 1 0 17020 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_183
timestamp 1646674385
transform 1 0 17940 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1744_
timestamp 1646674385
transform 1 0 17112 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2340__A
timestamp 1646674385
transform -1 0 19872 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1646674385
transform 1 0 18492 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1646674385
transform 1 0 19044 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_197
timestamp 1646674385
transform 1 0 19228 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_201
timestamp 1646674385
transform 1 0 19596 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_204
timestamp 1646674385
transform 1 0 19872 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1646674385
transform 1 0 19136 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_prog_clk
timestamp 1646674385
transform 1 0 20240 0 1 46240
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_84_228
timestamp 1646674385
transform 1 0 22080 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_248
timestamp 1646674385
transform 1 0 23920 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2687_
timestamp 1646674385
transform 1 0 22448 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_84_262
timestamp 1646674385
transform 1 0 25208 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_269
timestamp 1646674385
transform 1 0 25852 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1646674385
transform 1 0 24288 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1712_
timestamp 1646674385
transform 1 0 24380 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2358_
timestamp 1646674385
transform 1 0 25576 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_281
timestamp 1646674385
transform 1 0 26956 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_293
timestamp 1646674385
transform 1 0 28060 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_305
timestamp 1646674385
transform 1 0 29164 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_309
timestamp 1646674385
transform 1 0 29532 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1646674385
transform 1 0 29440 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_321
timestamp 1646674385
transform 1 0 30636 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1646674385
transform -1 0 32016 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1646674385
transform -1 0 1564 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1646674385
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1646674385
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_17
timestamp 1646674385
transform 1 0 2668 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_5
timestamp 1646674385
transform 1 0 1564 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1646674385
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1646674385
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1646674385
transform 1 0 3588 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1646674385
transform 1 0 4692 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_25
timestamp 1646674385
transform 1 0 3404 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1646674385
transform 1 0 3772 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1646674385
transform 1 0 4876 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1646674385
transform 1 0 3680 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1646674385
transform 1 0 5796 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1646674385
transform 1 0 6164 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1646674385
transform 1 0 6348 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_53
timestamp 1646674385
transform 1 0 5980 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_61
timestamp 1646674385
transform 1 0 6716 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1646674385
transform 1 0 6256 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_69
timestamp 1646674385
transform 1 0 7452 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_79
timestamp 1646674385
transform 1 0 8372 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1646674385
transform 1 0 8740 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2647_
timestamp 1646674385
transform -1 0 8372 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2648_
timestamp 1646674385
transform 1 0 7728 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_85_88
timestamp 1646674385
transform 1 0 9200 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_101
timestamp 1646674385
transform 1 0 10396 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1646674385
transform 1 0 8924 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_97
timestamp 1646674385
transform 1 0 10028 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1646674385
transform 1 0 8832 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2649_
timestamp 1646674385
transform 1 0 9568 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2651_
timestamp 1646674385
transform 1 0 10488 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_prog_clk_A
timestamp 1646674385
transform 1 0 11592 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_108
timestamp 1646674385
transform 1 0 11040 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_113
timestamp 1646674385
transform 1 0 11500 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_116
timestamp 1646674385
transform 1 0 11776 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_118
timestamp 1646674385
transform 1 0 11960 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1646674385
transform 1 0 11408 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2665_
timestamp 1646674385
transform 1 0 12144 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2602__CLK
timestamp 1646674385
transform -1 0 14260 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_136
timestamp 1646674385
transform 1 0 13616 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_126
timestamp 1646674385
transform 1 0 12696 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_136
timestamp 1646674385
transform 1 0 13616 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_143
timestamp 1646674385
transform 1 0 14260 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1646674385
transform 1 0 13984 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1754_
timestamp 1646674385
transform -1 0 13616 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2666_
timestamp 1646674385
transform 1 0 13984 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_prog_clk_A
timestamp 1646674385
transform 1 0 14812 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_156
timestamp 1646674385
transform 1 0 15456 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_160
timestamp 1646674385
transform 1 0 15824 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_164
timestamp 1646674385
transform 1 0 16192 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_151
timestamp 1646674385
transform 1 0 14996 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2057_
timestamp 1646674385
transform -1 0 16192 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2668_
timestamp 1646674385
transform 1 0 15364 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_85_185
timestamp 1646674385
transform 1 0 18124 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_171
timestamp 1646674385
transform 1 0 16836 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_175
timestamp 1646674385
transform 1 0 17204 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1646674385
transform 1 0 16560 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2669_
timestamp 1646674385
transform -1 0 18124 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2670_
timestamp 1646674385
transform 1 0 17296 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_85_207
timestamp 1646674385
transform 1 0 20148 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_192
timestamp 1646674385
transform 1 0 18768 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_197
timestamp 1646674385
transform 1 0 19228 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_201
timestamp 1646674385
transform 1 0 19596 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1646674385
transform 1 0 19136 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2685_
timestamp 1646674385
transform 1 0 18676 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2686_
timestamp 1646674385
transform -1 0 21160 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2339__A3
timestamp 1646674385
transform -1 0 20700 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_213
timestamp 1646674385
transform 1 0 20700 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_220
timestamp 1646674385
transform 1 0 21344 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_218
timestamp 1646674385
transform 1 0 21160 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_224
timestamp 1646674385
transform 1 0 21712 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1646674385
transform 1 0 21712 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1715_
timestamp 1646674385
transform 1 0 21804 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2355_
timestamp 1646674385
transform 1 0 21068 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2688_
timestamp 1646674385
transform 1 0 21804 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_85_234
timestamp 1646674385
transform 1 0 22632 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_86_241
timestamp 1646674385
transform 1 0 23276 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_249
timestamp 1646674385
transform 1 0 24012 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2613_
timestamp 1646674385
transform 1 0 23368 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2613__D
timestamp 1646674385
transform -1 0 25392 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_258
timestamp 1646674385
transform 1 0 24840 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_264
timestamp 1646674385
transform 1 0 25392 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_253
timestamp 1646674385
transform 1 0 24380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_265
timestamp 1646674385
transform 1 0 25484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1646674385
transform 1 0 24288 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_276
timestamp 1646674385
transform 1 0 26496 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1646674385
transform 1 0 26956 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_277
timestamp 1646674385
transform 1 0 26588 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_289
timestamp 1646674385
transform 1 0 27692 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1646674385
transform 1 0 26864 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_293
timestamp 1646674385
transform 1 0 28060 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_305
timestamp 1646674385
transform 1 0 29164 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1646674385
transform 1 0 28796 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1646674385
transform 1 0 29348 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_309
timestamp 1646674385
transform 1 0 29532 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1646674385
transform 1 0 29440 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2575__A
timestamp 1646674385
transform 1 0 30544 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_85_317
timestamp 1646674385
transform 1 0 30268 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_322
timestamp 1646674385
transform 1 0 30728 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_329
timestamp 1646674385
transform 1 0 31372 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_321
timestamp 1646674385
transform 1 0 30636 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1646674385
transform -1 0 32016 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1646674385
transform -1 0 32016 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2575_
timestamp 1646674385
transform -1 0 31372 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_87_19
timestamp 1646674385
transform 1 0 2852 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_7
timestamp 1646674385
transform 1 0 1748 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1646674385
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1646674385
transform 1 0 1380 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_27
timestamp 1646674385
transform 1 0 3588 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_29
timestamp 1646674385
transform 1 0 3772 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_41
timestamp 1646674385
transform 1 0 4876 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1646674385
transform 1 0 3680 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1646674385
transform 1 0 5980 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1646674385
transform 1 0 6348 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1646674385
transform 1 0 6256 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1646674385
transform 1 0 7452 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_81
timestamp 1646674385
transform 1 0 8556 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_100
timestamp 1646674385
transform 1 0 10304 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_88
timestamp 1646674385
transform 1 0 9200 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1646674385
transform 1 0 8832 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  output53
timestamp 1646674385
transform 1 0 8924 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_prog_clk_A
timestamp 1646674385
transform -1 0 11868 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_113
timestamp 1646674385
transform 1 0 11500 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_117
timestamp 1646674385
transform 1 0 11868 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1646674385
transform 1 0 11408 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_129
timestamp 1646674385
transform 1 0 12972 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_137
timestamp 1646674385
transform 1 0 13708 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_141
timestamp 1646674385
transform 1 0 14076 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1646674385
transform 1 0 13984 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_prog_clk_A
timestamp 1646674385
transform -1 0 15456 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_153
timestamp 1646674385
transform 1 0 15180 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_156
timestamp 1646674385
transform 1 0 15456 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_163
timestamp 1646674385
transform 1 0 16100 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2059_
timestamp 1646674385
transform 1 0 15824 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1646674385
transform -1 0 17112 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_prog_clk_A
timestamp 1646674385
transform -1 0 18216 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1646674385
transform 1 0 16468 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_87_169
timestamp 1646674385
transform 1 0 16652 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_87_174
timestamp 1646674385
transform 1 0 17112 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_182
timestamp 1646674385
transform 1 0 17848 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_87_186
timestamp 1646674385
transform 1 0 18216 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1646674385
transform 1 0 16560 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_prog_clk_A
timestamp 1646674385
transform -1 0 20240 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_prog_clk_A
timestamp 1646674385
transform -1 0 19596 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_194
timestamp 1646674385
transform 1 0 18952 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_197
timestamp 1646674385
transform 1 0 19228 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_201
timestamp 1646674385
transform 1 0 19596 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_205
timestamp 1646674385
transform 1 0 19964 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_208
timestamp 1646674385
transform 1 0 20240 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1646674385
transform 1 0 19136 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_220
timestamp 1646674385
transform 1 0 21344 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_225
timestamp 1646674385
transform 1 0 21804 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1646674385
transform 1 0 21712 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_237
timestamp 1646674385
transform 1 0 22908 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_249
timestamp 1646674385
transform 1 0 24012 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_87_253
timestamp 1646674385
transform 1 0 24380 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_262
timestamp 1646674385
transform 1 0 25208 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1646674385
transform 1 0 24288 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  output54
timestamp 1646674385
transform 1 0 24932 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_87_274
timestamp 1646674385
transform 1 0 26312 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1646674385
transform 1 0 26956 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1646674385
transform 1 0 26864 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_293
timestamp 1646674385
transform 1 0 28060 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_305
timestamp 1646674385
transform 1 0 29164 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_309
timestamp 1646674385
transform 1 0 29532 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1646674385
transform 1 0 29440 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_321
timestamp 1646674385
transform 1 0 30636 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_325
timestamp 1646674385
transform 1 0 31004 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_329
timestamp 1646674385
transform 1 0 31372 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1646674385
transform -1 0 32016 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output43
timestamp 1646674385
transform -1 0 31372 0 -1 48416
box -38 -48 314 592
<< labels >>
rlabel metal1 s 0 1026 800 1082 6 bi_u1y0n_L1[0]
port 0 nsew signal input
rlabel metal1 s 0 41826 800 41882 6 bi_u1y0n_L1[10]
port 1 nsew signal input
rlabel metal1 s 0 45906 800 45962 6 bi_u1y0n_L1[11]
port 2 nsew signal input
rlabel metal1 s 0 5106 800 5162 6 bi_u1y0n_L1[1]
port 3 nsew signal input
rlabel metal1 s 0 9186 800 9242 6 bi_u1y0n_L1[2]
port 4 nsew signal input
rlabel metal1 s 0 13266 800 13322 6 bi_u1y0n_L1[3]
port 5 nsew signal input
rlabel metal1 s 0 17346 800 17402 6 bi_u1y0n_L1[4]
port 6 nsew signal input
rlabel metal1 s 0 21426 800 21482 6 bi_u1y0n_L1[5]
port 7 nsew signal input
rlabel metal1 s 0 25506 800 25562 6 bi_u1y0n_L1[6]
port 8 nsew signal input
rlabel metal1 s 0 29586 800 29642 6 bi_u1y0n_L1[7]
port 9 nsew signal input
rlabel metal1 s 0 33666 800 33722 6 bi_u1y0n_L1[8]
port 10 nsew signal input
rlabel metal1 s 0 37746 800 37802 6 bi_u1y0n_L1[9]
port 11 nsew signal input
rlabel metal1 s 0 3066 800 3122 6 bi_u1y0s_L1[0]
port 12 nsew signal input
rlabel metal1 s 0 43866 800 43922 6 bi_u1y0s_L1[10]
port 13 nsew signal input
rlabel metal1 s 0 47946 800 48002 6 bi_u1y0s_L1[11]
port 14 nsew signal input
rlabel metal1 s 0 7146 800 7202 6 bi_u1y0s_L1[1]
port 15 nsew signal input
rlabel metal1 s 0 11226 800 11282 6 bi_u1y0s_L1[2]
port 16 nsew signal input
rlabel metal1 s 0 15306 800 15362 6 bi_u1y0s_L1[3]
port 17 nsew signal input
rlabel metal1 s 0 19386 800 19442 6 bi_u1y0s_L1[4]
port 18 nsew signal input
rlabel metal1 s 0 23466 800 23522 6 bi_u1y0s_L1[5]
port 19 nsew signal input
rlabel metal1 s 0 27546 800 27602 6 bi_u1y0s_L1[6]
port 20 nsew signal input
rlabel metal1 s 0 31626 800 31682 6 bi_u1y0s_L1[7]
port 21 nsew signal input
rlabel metal1 s 0 35706 800 35762 6 bi_u1y0s_L1[8]
port 22 nsew signal input
rlabel metal1 s 0 39786 800 39842 6 bi_u1y0s_L1[9]
port 23 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 clk
port 24 nsew signal input
rlabel metal1 s 32320 1026 33120 1082 6 cu_x0y0n_L1[0]
port 25 nsew signal tristate
rlabel metal1 s 32320 41826 33120 41882 6 cu_x0y0n_L1[10]
port 26 nsew signal tristate
rlabel metal1 s 32320 45906 33120 45962 6 cu_x0y0n_L1[11]
port 27 nsew signal tristate
rlabel metal1 s 32320 5106 33120 5162 6 cu_x0y0n_L1[1]
port 28 nsew signal tristate
rlabel metal1 s 32320 9186 33120 9242 6 cu_x0y0n_L1[2]
port 29 nsew signal tristate
rlabel metal1 s 32320 13266 33120 13322 6 cu_x0y0n_L1[3]
port 30 nsew signal tristate
rlabel metal1 s 32320 17346 33120 17402 6 cu_x0y0n_L1[4]
port 31 nsew signal tristate
rlabel metal1 s 32320 21426 33120 21482 6 cu_x0y0n_L1[5]
port 32 nsew signal tristate
rlabel metal1 s 32320 25506 33120 25562 6 cu_x0y0n_L1[6]
port 33 nsew signal tristate
rlabel metal1 s 32320 29586 33120 29642 6 cu_x0y0n_L1[7]
port 34 nsew signal tristate
rlabel metal1 s 32320 33666 33120 33722 6 cu_x0y0n_L1[8]
port 35 nsew signal tristate
rlabel metal1 s 32320 37746 33120 37802 6 cu_x0y0n_L1[9]
port 36 nsew signal tristate
rlabel metal1 s 32320 3066 33120 3122 6 cu_x0y0s_L1[0]
port 37 nsew signal tristate
rlabel metal1 s 32320 43866 33120 43922 6 cu_x0y0s_L1[10]
port 38 nsew signal tristate
rlabel metal1 s 32320 47946 33120 48002 6 cu_x0y0s_L1[11]
port 39 nsew signal tristate
rlabel metal1 s 32320 7146 33120 7202 6 cu_x0y0s_L1[1]
port 40 nsew signal tristate
rlabel metal1 s 32320 11226 33120 11282 6 cu_x0y0s_L1[2]
port 41 nsew signal tristate
rlabel metal1 s 32320 15306 33120 15362 6 cu_x0y0s_L1[3]
port 42 nsew signal tristate
rlabel metal1 s 32320 19386 33120 19442 6 cu_x0y0s_L1[4]
port 43 nsew signal tristate
rlabel metal1 s 32320 23466 33120 23522 6 cu_x0y0s_L1[5]
port 44 nsew signal tristate
rlabel metal1 s 32320 27546 33120 27602 6 cu_x0y0s_L1[6]
port 45 nsew signal tristate
rlabel metal1 s 32320 31626 33120 31682 6 cu_x0y0s_L1[7]
port 46 nsew signal tristate
rlabel metal1 s 32320 35706 33120 35762 6 cu_x0y0s_L1[8]
port 47 nsew signal tristate
rlabel metal1 s 32320 39786 33120 39842 6 cu_x0y0s_L1[9]
port 48 nsew signal tristate
rlabel metal2 s 30378 0 30434 800 6 prog_clk
port 49 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 prog_din
port 50 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 prog_done
port 51 nsew signal input
rlabel metal2 s 8298 48160 8354 48960 6 prog_dout
port 52 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 prog_rst
port 53 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 prog_we
port 54 nsew signal input
rlabel metal2 s 24858 48160 24914 48960 6 prog_we_o
port 55 nsew signal tristate
rlabel metal4 s 6095 496 6415 48464 6 vccd1
port 56 nsew power input
rlabel metal4 s 16399 496 16719 48464 6 vccd1
port 56 nsew power input
rlabel metal4 s 26703 496 27023 48464 6 vccd1
port 56 nsew power input
rlabel metal4 s 11247 496 11567 48464 6 vssd1
port 57 nsew ground input
rlabel metal4 s 21551 496 21871 48464 6 vssd1
port 57 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 33120 48960
<< end >>
