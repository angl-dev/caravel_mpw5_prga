magic
tech sky130A
magscale 1 2
timestamp 1654095952
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 273254 700748 273260 700800
rect 273312 700788 273318 700800
rect 348786 700788 348792 700800
rect 273312 700760 348792 700788
rect 273312 700748 273318 700760
rect 348786 700748 348792 700760
rect 348844 700748 348850 700800
rect 52454 700680 52460 700732
rect 52512 700720 52518 700732
rect 170306 700720 170312 700732
rect 52512 700692 170312 700720
rect 52512 700680 52518 700692
rect 170306 700680 170312 700692
rect 170364 700680 170370 700732
rect 292574 700680 292580 700732
rect 292632 700720 292638 700732
rect 413646 700720 413652 700732
rect 292632 700692 413652 700720
rect 292632 700680 292638 700692
rect 413646 700680 413652 700692
rect 413704 700680 413710 700732
rect 62114 700612 62120 700664
rect 62172 700652 62178 700664
rect 235166 700652 235172 700664
rect 62172 700624 235172 700652
rect 62172 700612 62178 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 253934 700612 253940 700664
rect 253992 700652 253998 700664
rect 283834 700652 283840 700664
rect 253992 700624 283840 700652
rect 253992 700612 253998 700624
rect 283834 700612 283840 700624
rect 283892 700612 283898 700664
rect 311894 700612 311900 700664
rect 311952 700652 311958 700664
rect 478506 700652 478512 700664
rect 311952 700624 478512 700652
rect 311952 700612 311958 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 81434 700544 81440 700596
rect 81492 700584 81498 700596
rect 300118 700584 300124 700596
rect 81492 700556 300124 700584
rect 81492 700544 81498 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 340874 700544 340880 700596
rect 340932 700584 340938 700596
rect 543458 700584 543464 700596
rect 340932 700556 543464 700584
rect 340932 700544 340938 700556
rect 543458 700544 543464 700556
rect 543516 700544 543522 700596
rect 100754 700476 100760 700528
rect 100812 700516 100818 700528
rect 364978 700516 364984 700528
rect 100812 700488 364984 700516
rect 100812 700476 100818 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 120074 700408 120080 700460
rect 120132 700448 120138 700460
rect 429838 700448 429844 700460
rect 120132 700420 429844 700448
rect 120132 700408 120138 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 139394 700340 139400 700392
rect 139452 700380 139458 700392
rect 494790 700380 494796 700392
rect 139452 700352 494796 700380
rect 139452 700340 139458 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 514754 700340 514760 700392
rect 514812 700380 514818 700392
rect 527174 700380 527180 700392
rect 514812 700352 527180 700380
rect 514812 700340 514818 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 23566 700272 23572 700324
rect 23624 700312 23630 700324
rect 40494 700312 40500 700324
rect 23624 700284 40500 700312
rect 23624 700272 23630 700284
rect 40494 700272 40500 700284
rect 40552 700272 40558 700324
rect 166994 700272 167000 700324
rect 167052 700312 167058 700324
rect 559650 700312 559656 700324
rect 167052 700284 559656 700312
rect 167052 700272 167058 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 541618 696940 541624 696992
rect 541676 696980 541682 696992
rect 580166 696980 580172 696992
rect 541676 696952 580172 696980
rect 541676 696940 541682 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 558178 683136 558184 683188
rect 558236 683176 558242 683188
rect 580166 683176 580172 683188
rect 558236 683148 580172 683176
rect 558236 683136 558242 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 556798 670692 556804 670744
rect 556856 670732 556862 670744
rect 580166 670732 580172 670744
rect 556856 670704 580172 670732
rect 556856 670692 556862 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 153194 657840 153200 657892
rect 153252 657880 153258 657892
rect 225782 657880 225788 657892
rect 153252 657852 225788 657880
rect 153252 657840 153258 657852
rect 225782 657840 225788 657852
rect 225840 657840 225846 657892
rect 331214 657840 331220 657892
rect 331272 657880 331278 657892
rect 447226 657880 447232 657892
rect 331272 657852 447232 657880
rect 331272 657840 331278 657852
rect 447226 657840 447232 657852
rect 447284 657840 447290 657892
rect 88334 657772 88340 657824
rect 88392 657812 88398 657824
rect 216122 657812 216128 657824
rect 88392 657784 216128 657812
rect 88392 657772 88398 657784
rect 216122 657772 216128 657784
rect 216180 657772 216186 657824
rect 218054 657772 218060 657824
rect 218112 657812 218118 657824
rect 235350 657812 235356 657824
rect 218112 657784 235356 657812
rect 218112 657772 218118 657784
rect 235350 657772 235356 657784
rect 235408 657772 235414 657824
rect 266354 657772 266360 657824
rect 266412 657812 266418 657824
rect 427998 657812 428004 657824
rect 266412 657784 428004 657812
rect 266412 657772 266418 657784
rect 427998 657772 428004 657784
rect 428056 657772 428062 657824
rect 23474 657704 23480 657756
rect 23532 657744 23538 657756
rect 196894 657744 196900 657756
rect 23532 657716 196900 657744
rect 23532 657704 23538 657716
rect 196894 657704 196900 657716
rect 196952 657704 196958 657756
rect 201494 657704 201500 657756
rect 201552 657744 201558 657756
rect 408678 657744 408684 657756
rect 201552 657716 408684 657744
rect 201552 657704 201558 657716
rect 408678 657704 408684 657716
rect 408736 657704 408742 657756
rect 43438 657636 43444 657688
rect 43496 657676 43502 657688
rect 104894 657676 104900 657688
rect 43496 657648 104900 657676
rect 43496 657636 43502 657648
rect 104894 657636 104900 657648
rect 104952 657636 104958 657688
rect 136634 657636 136640 657688
rect 136692 657676 136698 657688
rect 399110 657676 399116 657688
rect 136692 657648 399116 657676
rect 136692 657636 136698 657648
rect 399110 657636 399116 657648
rect 399168 657636 399174 657688
rect 71774 657568 71780 657620
rect 71832 657608 71838 657620
rect 389450 657608 389456 657620
rect 71832 657580 389456 657608
rect 71832 657568 71838 657580
rect 389450 657568 389456 657580
rect 389508 657568 389514 657620
rect 462314 657568 462320 657620
rect 462372 657608 462378 657620
rect 485774 657608 485780 657620
rect 462372 657580 485780 657608
rect 462372 657568 462378 657580
rect 485774 657568 485780 657580
rect 485832 657568 485838 657620
rect 6914 657500 6920 657552
rect 6972 657540 6978 657552
rect 370222 657540 370228 657552
rect 6972 657512 370228 657540
rect 6972 657500 6978 657512
rect 370222 657500 370228 657512
rect 370280 657500 370286 657552
rect 397454 657500 397460 657552
rect 397512 657540 397518 657552
rect 466454 657540 466460 657552
rect 397512 657512 466460 657540
rect 397512 657500 397518 657512
rect 466454 657500 466460 657512
rect 466512 657500 466518 657552
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4890 632108 4896 632120
rect 2832 632080 4896 632108
rect 2832 632068 2838 632080
rect 4890 632068 4896 632080
rect 4948 632068 4954 632120
rect 573450 630640 573456 630692
rect 573508 630680 573514 630692
rect 579982 630680 579988 630692
rect 573508 630652 579988 630680
rect 573508 630640 573514 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 573358 616836 573364 616888
rect 573416 616876 573422 616888
rect 580166 616876 580172 616888
rect 573416 616848 580172 616876
rect 573416 616836 573422 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 614048 3424 614100
rect 3476 614088 3482 614100
rect 17034 614088 17040 614100
rect 3476 614060 17040 614088
rect 3476 614048 3482 614060
rect 17034 614048 17040 614060
rect 17092 614048 17098 614100
rect 542262 601604 542268 601656
rect 542320 601644 542326 601656
rect 580258 601644 580264 601656
rect 542320 601616 580264 601644
rect 542320 601604 542326 601616
rect 580258 601604 580264 601616
rect 580316 601604 580322 601656
rect 541802 590656 541808 590708
rect 541860 590696 541866 590708
rect 579798 590696 579804 590708
rect 541860 590668 579804 590696
rect 541860 590656 541866 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3418 590588 3424 590640
rect 3476 590628 3482 590640
rect 17862 590628 17868 590640
rect 3476 590600 17868 590628
rect 3476 590588 3482 590600
rect 17862 590588 17868 590600
rect 17920 590588 17926 590640
rect 3142 579776 3148 579828
rect 3200 579816 3206 579828
rect 8938 579816 8944 579828
rect 3200 579788 8944 579816
rect 3200 579776 3206 579788
rect 8938 579776 8944 579788
rect 8996 579776 9002 579828
rect 572070 576852 572076 576904
rect 572128 576892 572134 576904
rect 580166 576892 580172 576904
rect 572128 576864 580172 576892
rect 572128 576852 572134 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 15838 565904 15844 565956
rect 15896 565944 15902 565956
rect 17862 565944 17868 565956
rect 15896 565916 17868 565944
rect 15896 565904 15902 565916
rect 17862 565904 17868 565916
rect 17920 565904 17926 565956
rect 571978 563048 571984 563100
rect 572036 563088 572042 563100
rect 579798 563088 579804 563100
rect 572036 563060 579804 563088
rect 572036 563048 572042 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 2958 554684 2964 554736
rect 3016 554724 3022 554736
rect 15838 554724 15844 554736
rect 3016 554696 15844 554724
rect 3016 554684 3022 554696
rect 15838 554684 15844 554696
rect 15896 554684 15902 554736
rect 541710 538160 541716 538212
rect 541768 538200 541774 538212
rect 580166 538200 580172 538212
rect 541768 538172 580172 538200
rect 541768 538160 541774 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 558270 524424 558276 524476
rect 558328 524464 558334 524476
rect 580166 524464 580172 524476
rect 558328 524436 580172 524464
rect 558328 524424 558334 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 502256 3332 502308
rect 3384 502296 3390 502308
rect 17218 502296 17224 502308
rect 3384 502268 17224 502296
rect 3384 502256 3390 502268
rect 17218 502256 17224 502268
rect 17276 502256 17282 502308
rect 542262 494096 542268 494148
rect 542320 494136 542326 494148
rect 548518 494136 548524 494148
rect 542320 494108 548524 494136
rect 542320 494096 542326 494108
rect 548518 494096 548524 494108
rect 548576 494096 548582 494148
rect 541618 485732 541624 485784
rect 541676 485772 541682 485784
rect 580166 485772 580172 485784
rect 541676 485744 580172 485772
rect 541676 485732 541682 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 2774 474920 2780 474972
rect 2832 474960 2838 474972
rect 4982 474960 4988 474972
rect 2832 474932 4988 474960
rect 2832 474920 2838 474932
rect 4982 474920 4988 474932
rect 5040 474920 5046 474972
rect 542262 471112 542268 471164
rect 542320 471152 542326 471164
rect 547138 471152 547144 471164
rect 542320 471124 547144 471152
rect 542320 471112 542326 471124
rect 547138 471112 547144 471124
rect 547196 471112 547202 471164
rect 7558 470568 7564 470620
rect 7616 470608 7622 470620
rect 17862 470608 17868 470620
rect 7616 470580 17868 470608
rect 7616 470568 7622 470580
rect 17862 470568 17868 470580
rect 17920 470568 17926 470620
rect 542170 458192 542176 458244
rect 542228 458232 542234 458244
rect 545758 458232 545764 458244
rect 542228 458204 545764 458232
rect 542228 458192 542234 458204
rect 545758 458192 545764 458204
rect 545816 458192 545822 458244
rect 556890 456764 556896 456816
rect 556948 456804 556954 456816
rect 580166 456804 580172 456816
rect 556948 456776 580172 456804
rect 556948 456764 556954 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 17402 449868 17408 449880
rect 3384 449840 17408 449868
rect 3384 449828 3390 449840
rect 17402 449828 17408 449840
rect 17460 449828 17466 449880
rect 541434 447312 541440 447364
rect 541492 447352 541498 447364
rect 544378 447352 544384 447364
rect 541492 447324 544384 447352
rect 541492 447312 541498 447324
rect 544378 447312 544384 447324
rect 544436 447312 544442 447364
rect 541894 431876 541900 431928
rect 541952 431916 541958 431928
rect 579614 431916 579620 431928
rect 541952 431888 579620 431916
rect 541952 431876 541958 431888
rect 579614 431876 579620 431888
rect 579672 431876 579678 431928
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 9030 422328 9036 422340
rect 3016 422300 9036 422328
rect 3016 422288 3022 422300
rect 9030 422288 9036 422300
rect 9088 422288 9094 422340
rect 542998 404336 543004 404388
rect 543056 404376 543062 404388
rect 580166 404376 580172 404388
rect 543056 404348 580172 404376
rect 543056 404336 543062 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 400120 3516 400172
rect 3568 400160 3574 400172
rect 17862 400160 17868 400172
rect 3568 400132 17868 400160
rect 3568 400120 3574 400132
rect 17862 400120 17868 400132
rect 17920 400120 17926 400172
rect 542262 400120 542268 400172
rect 542320 400160 542326 400172
rect 558178 400160 558184 400172
rect 542320 400132 558184 400160
rect 542320 400120 542326 400132
rect 558178 400120 558184 400132
rect 558236 400120 558242 400172
rect 3510 398760 3516 398812
rect 3568 398800 3574 398812
rect 17218 398800 17224 398812
rect 3568 398772 17224 398800
rect 3568 398760 3574 398772
rect 17218 398760 17224 398772
rect 17276 398760 17282 398812
rect 542262 389104 542268 389156
rect 542320 389144 542326 389156
rect 573450 389144 573456 389156
rect 542320 389116 573456 389144
rect 542320 389104 542326 389116
rect 573450 389104 573456 389116
rect 573508 389104 573514 389156
rect 541802 379448 541808 379500
rect 541860 379488 541866 379500
rect 579798 379488 579804 379500
rect 541860 379460 579804 379488
rect 541860 379448 541866 379460
rect 579798 379448 579804 379460
rect 579856 379448 579862 379500
rect 3602 376660 3608 376712
rect 3660 376700 3666 376712
rect 16758 376700 16764 376712
rect 3660 376672 16764 376700
rect 3660 376660 3666 376672
rect 16758 376660 16764 376672
rect 16816 376660 16822 376712
rect 541894 376660 541900 376712
rect 541952 376700 541958 376712
rect 572070 376700 572076 376712
rect 541952 376672 572076 376700
rect 541952 376660 541958 376672
rect 572070 376660 572076 376672
rect 572128 376660 572134 376712
rect 3142 371288 3148 371340
rect 3200 371328 3206 371340
rect 6178 371328 6184 371340
rect 3200 371300 6184 371328
rect 3200 371288 3206 371300
rect 6178 371288 6184 371300
rect 6236 371288 6242 371340
rect 3694 353200 3700 353252
rect 3752 353240 3758 353252
rect 17862 353240 17868 353252
rect 3752 353212 17868 353240
rect 3752 353200 3758 353212
rect 17862 353200 17868 353212
rect 17920 353200 17926 353252
rect 541250 353200 541256 353252
rect 541308 353240 541314 353252
rect 558270 353240 558276 353252
rect 541308 353212 558276 353240
rect 541308 353200 541314 353212
rect 558270 353200 558276 353212
rect 558328 353200 558334 353252
rect 558178 351908 558184 351960
rect 558236 351948 558242 351960
rect 580166 351948 580172 351960
rect 558236 351920 580172 351948
rect 558236 351908 558242 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3510 346196 3516 346248
rect 3568 346236 3574 346248
rect 7558 346236 7564 346248
rect 3568 346208 7564 346236
rect 3568 346196 3574 346208
rect 7558 346196 7564 346208
rect 7616 346196 7622 346248
rect 541986 342184 541992 342236
rect 542044 342224 542050 342236
rect 580350 342224 580356 342236
rect 542044 342196 580356 342224
rect 542044 342184 542050 342196
rect 580350 342184 580356 342196
rect 580408 342184 580414 342236
rect 3786 329740 3792 329792
rect 3844 329780 3850 329792
rect 17862 329780 17868 329792
rect 3844 329752 17868 329780
rect 3844 329740 3850 329752
rect 17862 329740 17868 329752
rect 17920 329740 17926 329792
rect 542262 329740 542268 329792
rect 542320 329780 542326 329792
rect 580442 329780 580448 329792
rect 542320 329752 580448 329780
rect 542320 329740 542326 329752
rect 580442 329740 580448 329752
rect 580500 329740 580506 329792
rect 541710 325592 541716 325644
rect 541768 325632 541774 325644
rect 580166 325632 580172 325644
rect 541768 325604 580172 325632
rect 541768 325592 541774 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 17218 318832 17224 318844
rect 3384 318804 17224 318832
rect 3384 318792 3390 318804
rect 17218 318792 17224 318804
rect 17276 318792 17282 318844
rect 3878 306280 3884 306332
rect 3936 306320 3942 306332
rect 17862 306320 17868 306332
rect 3936 306292 17868 306320
rect 3936 306280 3942 306292
rect 17862 306280 17868 306292
rect 17920 306280 17926 306332
rect 541894 306280 541900 306332
rect 541952 306320 541958 306332
rect 580534 306320 580540 306332
rect 541952 306292 580540 306320
rect 541952 306280 541958 306292
rect 580534 306280 580540 306292
rect 580592 306280 580598 306332
rect 572070 298120 572076 298172
rect 572128 298160 572134 298172
rect 579982 298160 579988 298172
rect 572128 298132 579988 298160
rect 572128 298120 572134 298132
rect 579982 298120 579988 298132
rect 580040 298120 580046 298172
rect 3510 293904 3516 293956
rect 3568 293944 3574 293956
rect 17310 293944 17316 293956
rect 3568 293916 17316 293944
rect 3568 293904 3574 293916
rect 17310 293904 17316 293916
rect 17368 293904 17374 293956
rect 541342 293904 541348 293956
rect 541400 293944 541406 293956
rect 580350 293944 580356 293956
rect 541400 293916 580356 293944
rect 541400 293904 541406 293916
rect 580350 293904 580356 293916
rect 580408 293904 580414 293956
rect 3970 282820 3976 282872
rect 4028 282860 4034 282872
rect 16942 282860 16948 282872
rect 4028 282832 16948 282860
rect 4028 282820 4034 282832
rect 16942 282820 16948 282832
rect 17000 282820 17006 282872
rect 548518 273164 548524 273216
rect 548576 273204 548582 273216
rect 579890 273204 579896 273216
rect 548576 273176 579896 273204
rect 548576 273164 548582 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 541710 259360 541716 259412
rect 541768 259400 541774 259412
rect 579798 259400 579804 259412
rect 541768 259372 579804 259400
rect 541768 259360 541774 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3602 258000 3608 258052
rect 3660 258040 3666 258052
rect 17862 258040 17868 258052
rect 3660 258012 17868 258040
rect 3660 258000 3666 258012
rect 17862 258000 17868 258012
rect 17920 258000 17926 258052
rect 3694 246984 3700 247036
rect 3752 247024 3758 247036
rect 16758 247024 16764 247036
rect 3752 246996 16764 247024
rect 3752 246984 3758 246996
rect 16758 246984 16764 246996
rect 16816 246984 16822 247036
rect 573450 244264 573456 244316
rect 573508 244304 573514 244316
rect 580166 244304 580172 244316
rect 573508 244276 580172 244304
rect 573508 244264 573514 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 541618 233180 541624 233232
rect 541676 233220 541682 233232
rect 580166 233220 580172 233232
rect 541676 233192 580172 233220
rect 541676 233180 541682 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 541986 219376 541992 219428
rect 542044 219416 542050 219428
rect 579890 219416 579896 219428
rect 542044 219388 579896 219416
rect 542044 219376 542050 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 547138 193128 547144 193180
rect 547196 193168 547202 193180
rect 580166 193168 580172 193180
rect 547196 193140 580172 193168
rect 547196 193128 547202 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 4798 187620 4804 187672
rect 4856 187660 4862 187672
rect 17862 187660 17868 187672
rect 4856 187632 17868 187660
rect 4856 187620 4862 187632
rect 17862 187620 17868 187632
rect 17920 187620 17926 187672
rect 542262 187620 542268 187672
rect 542320 187660 542326 187672
rect 556798 187660 556804 187672
rect 542320 187632 556804 187660
rect 542320 187620 542326 187632
rect 556798 187620 556804 187632
rect 556856 187620 556862 187672
rect 541894 179324 541900 179376
rect 541952 179364 541958 179376
rect 580166 179364 580172 179376
rect 541952 179336 580172 179364
rect 541952 179324 541958 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 542262 175176 542268 175228
rect 542320 175216 542326 175228
rect 573358 175216 573364 175228
rect 542320 175188 573364 175216
rect 542320 175176 542326 175188
rect 573358 175176 573364 175188
rect 573416 175176 573422 175228
rect 4890 164160 4896 164212
rect 4948 164200 4954 164212
rect 17862 164200 17868 164212
rect 4948 164172 17868 164200
rect 4948 164160 4954 164172
rect 17862 164160 17868 164172
rect 17920 164160 17926 164212
rect 541986 164160 541992 164212
rect 542044 164200 542050 164212
rect 571978 164200 571984 164212
rect 542044 164172 571984 164200
rect 542044 164160 542050 164172
rect 571978 164160 571984 164172
rect 572036 164160 572042 164212
rect 545758 153144 545764 153196
rect 545816 153184 545822 153196
rect 580166 153184 580172 153196
rect 545816 153156 580172 153184
rect 545816 153144 545822 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 8938 139340 8944 139392
rect 8996 139380 9002 139392
rect 16942 139380 16948 139392
rect 8996 139352 16948 139380
rect 8996 139340 9002 139352
rect 16942 139340 16948 139352
rect 17000 139340 17006 139392
rect 541802 139340 541808 139392
rect 541860 139380 541866 139392
rect 580166 139380 580172 139392
rect 541860 139352 580172 139380
rect 541860 139340 541866 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 542262 139272 542268 139324
rect 542320 139312 542326 139324
rect 580258 139312 580264 139324
rect 542320 139284 580264 139312
rect 542320 139272 542326 139284
rect 580258 139272 580264 139284
rect 580316 139272 580322 139324
rect 542262 128256 542268 128308
rect 542320 128296 542326 128308
rect 556890 128296 556896 128308
rect 542320 128268 556896 128296
rect 542320 128256 542326 128268
rect 556890 128256 556896 128268
rect 556948 128256 556954 128308
rect 3418 115880 3424 115932
rect 3476 115920 3482 115932
rect 17862 115920 17868 115932
rect 3476 115892 17868 115920
rect 3476 115880 3482 115892
rect 17862 115880 17868 115892
rect 17920 115880 17926 115932
rect 540974 115676 540980 115728
rect 541032 115716 541038 115728
rect 542998 115716 543004 115728
rect 541032 115688 543004 115716
rect 541032 115676 541038 115688
rect 542998 115676 543004 115688
rect 543056 115676 543062 115728
rect 544378 113092 544384 113144
rect 544436 113132 544442 113144
rect 580166 113132 580172 113144
rect 544436 113104 580172 113132
rect 544436 113092 544442 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 541710 100648 541716 100700
rect 541768 100688 541774 100700
rect 579706 100688 579712 100700
rect 541768 100660 579712 100688
rect 541768 100648 541774 100660
rect 579706 100648 579712 100660
rect 579764 100648 579770 100700
rect 4982 92420 4988 92472
rect 5040 92460 5046 92472
rect 17862 92460 17868 92472
rect 5040 92432 17868 92460
rect 5040 92420 5046 92432
rect 17862 92420 17868 92432
rect 17920 92420 17926 92472
rect 542262 92420 542268 92472
rect 542320 92460 542326 92472
rect 558178 92460 558184 92472
rect 542320 92432 558184 92460
rect 542320 92420 542326 92432
rect 558178 92420 558184 92432
rect 558236 92420 558242 92472
rect 542262 79976 542268 80028
rect 542320 80016 542326 80028
rect 572070 80016 572076 80028
rect 542320 79988 572076 80016
rect 542320 79976 542326 79988
rect 572070 79976 572076 79988
rect 572128 79976 572134 80028
rect 9030 68960 9036 69012
rect 9088 69000 9094 69012
rect 17862 69000 17868 69012
rect 9088 68972 17868 69000
rect 9088 68960 9094 68972
rect 17862 68960 17868 68972
rect 17920 68960 17926 69012
rect 542262 68960 542268 69012
rect 542320 69000 542326 69012
rect 573450 69000 573456 69012
rect 542320 68972 573456 69000
rect 542320 68960 542326 68972
rect 573450 68960 573456 68972
rect 573508 68960 573514 69012
rect 542262 56516 542268 56568
rect 542320 56556 542326 56568
rect 580350 56556 580356 56568
rect 542320 56528 580356 56556
rect 542320 56516 542326 56528
rect 580350 56516 580356 56528
rect 580408 56516 580414 56568
rect 6178 45500 6184 45552
rect 6236 45540 6242 45552
rect 16758 45540 16764 45552
rect 6236 45512 16764 45540
rect 6236 45500 6242 45512
rect 16758 45500 16764 45512
rect 16816 45500 16822 45552
rect 541894 45500 541900 45552
rect 541952 45540 541958 45552
rect 580442 45540 580448 45552
rect 541952 45512 580448 45540
rect 541952 45500 541958 45512
rect 580442 45500 580448 45512
rect 580500 45500 580506 45552
rect 542262 33056 542268 33108
rect 542320 33096 542326 33108
rect 580258 33096 580264 33108
rect 542320 33068 580264 33096
rect 542320 33056 542326 33068
rect 580258 33056 580264 33068
rect 580316 33056 580322 33108
rect 3878 22040 3884 22092
rect 3936 22080 3942 22092
rect 17862 22080 17868 22092
rect 3936 22052 17868 22080
rect 3936 22040 3942 22052
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 541986 22040 541992 22092
rect 542044 22080 542050 22092
rect 580534 22080 580540 22092
rect 542044 22052 580540 22080
rect 542044 22040 542050 22052
rect 580534 22040 580540 22052
rect 580592 22040 580598 22092
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 55858 13784 55864 13796
rect 3476 13756 55864 13784
rect 3476 13744 3482 13756
rect 55858 13744 55864 13756
rect 55916 13744 55922 13796
rect 279326 13744 279332 13796
rect 279384 13784 279390 13796
rect 580626 13784 580632 13796
rect 279384 13756 580632 13784
rect 279384 13744 279390 13756
rect 580626 13744 580632 13756
rect 580684 13744 580690 13796
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 427262 13716 427268 13728
rect 3568 13688 427268 13716
rect 3568 13676 3574 13688
rect 427262 13676 427268 13688
rect 427320 13676 427326 13728
rect 502150 13676 502156 13728
rect 502208 13716 502214 13728
rect 580258 13716 580264 13728
rect 502208 13688 580264 13716
rect 502208 13676 502214 13688
rect 580258 13676 580264 13688
rect 580316 13676 580322 13728
rect 3602 13608 3608 13660
rect 3660 13648 3666 13660
rect 352926 13648 352932 13660
rect 3660 13620 352932 13648
rect 3660 13608 3666 13620
rect 352926 13608 352932 13620
rect 352984 13608 352990 13660
rect 3694 13540 3700 13592
rect 3752 13580 3758 13592
rect 204346 13580 204352 13592
rect 3752 13552 204352 13580
rect 3752 13540 3758 13552
rect 204346 13540 204352 13552
rect 204404 13540 204410 13592
rect 3786 13472 3792 13524
rect 3844 13512 3850 13524
rect 130102 13512 130108 13524
rect 3844 13484 130108 13512
rect 3844 13472 3850 13484
rect 130102 13472 130108 13484
rect 130160 13472 130166 13524
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 273260 700748 273312 700800
rect 348792 700748 348844 700800
rect 52460 700680 52512 700732
rect 170312 700680 170364 700732
rect 292580 700680 292632 700732
rect 413652 700680 413704 700732
rect 62120 700612 62172 700664
rect 235172 700612 235224 700664
rect 253940 700612 253992 700664
rect 283840 700612 283892 700664
rect 311900 700612 311952 700664
rect 478512 700612 478564 700664
rect 81440 700544 81492 700596
rect 300124 700544 300176 700596
rect 340880 700544 340932 700596
rect 543464 700544 543516 700596
rect 100760 700476 100812 700528
rect 364984 700476 365036 700528
rect 120080 700408 120132 700460
rect 429844 700408 429896 700460
rect 139400 700340 139452 700392
rect 494796 700340 494848 700392
rect 514760 700340 514812 700392
rect 527180 700340 527232 700392
rect 23572 700272 23624 700324
rect 40500 700272 40552 700324
rect 167000 700272 167052 700324
rect 559656 700272 559708 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 541624 696940 541676 696992
rect 580172 696940 580224 696992
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 558184 683136 558236 683188
rect 580172 683136 580224 683188
rect 556804 670692 556856 670744
rect 580172 670692 580224 670744
rect 153200 657840 153252 657892
rect 225788 657840 225840 657892
rect 331220 657840 331272 657892
rect 447232 657840 447284 657892
rect 88340 657772 88392 657824
rect 216128 657772 216180 657824
rect 218060 657772 218112 657824
rect 235356 657772 235408 657824
rect 266360 657772 266412 657824
rect 428004 657772 428056 657824
rect 23480 657704 23532 657756
rect 196900 657704 196952 657756
rect 201500 657704 201552 657756
rect 408684 657704 408736 657756
rect 43444 657636 43496 657688
rect 104900 657636 104952 657688
rect 136640 657636 136692 657688
rect 399116 657636 399168 657688
rect 71780 657568 71832 657620
rect 389456 657568 389508 657620
rect 462320 657568 462372 657620
rect 485780 657568 485832 657620
rect 6920 657500 6972 657552
rect 370228 657500 370280 657552
rect 397460 657500 397512 657552
rect 466460 657500 466512 657552
rect 2780 632068 2832 632120
rect 4896 632068 4948 632120
rect 573456 630640 573508 630692
rect 579988 630640 580040 630692
rect 573364 616836 573416 616888
rect 580172 616836 580224 616888
rect 3424 614048 3476 614100
rect 17040 614048 17092 614100
rect 542268 601604 542320 601656
rect 580264 601604 580316 601656
rect 541808 590656 541860 590708
rect 579804 590656 579856 590708
rect 3424 590588 3476 590640
rect 17868 590588 17920 590640
rect 3148 579776 3200 579828
rect 8944 579776 8996 579828
rect 572076 576852 572128 576904
rect 580172 576852 580224 576904
rect 15844 565904 15896 565956
rect 17868 565904 17920 565956
rect 571984 563048 572036 563100
rect 579804 563048 579856 563100
rect 2964 554684 3016 554736
rect 15844 554684 15896 554736
rect 541716 538160 541768 538212
rect 580172 538160 580224 538212
rect 558276 524424 558328 524476
rect 580172 524424 580224 524476
rect 3332 502256 3384 502308
rect 17224 502256 17276 502308
rect 542268 494096 542320 494148
rect 548524 494096 548576 494148
rect 541624 485732 541676 485784
rect 580172 485732 580224 485784
rect 2780 474920 2832 474972
rect 4988 474920 5040 474972
rect 542268 471112 542320 471164
rect 547144 471112 547196 471164
rect 7564 470568 7616 470620
rect 17868 470568 17920 470620
rect 542176 458192 542228 458244
rect 545764 458192 545816 458244
rect 556896 456764 556948 456816
rect 580172 456764 580224 456816
rect 3332 449828 3384 449880
rect 17408 449828 17460 449880
rect 541440 447312 541492 447364
rect 544384 447312 544436 447364
rect 541900 431876 541952 431928
rect 579620 431876 579672 431928
rect 2964 422288 3016 422340
rect 9036 422288 9088 422340
rect 543004 404336 543056 404388
rect 580172 404336 580224 404388
rect 3516 400120 3568 400172
rect 17868 400120 17920 400172
rect 542268 400120 542320 400172
rect 558184 400120 558236 400172
rect 3516 398760 3568 398812
rect 17224 398760 17276 398812
rect 542268 389104 542320 389156
rect 573456 389104 573508 389156
rect 541808 379448 541860 379500
rect 579804 379448 579856 379500
rect 3608 376660 3660 376712
rect 16764 376660 16816 376712
rect 541900 376660 541952 376712
rect 572076 376660 572128 376712
rect 3148 371288 3200 371340
rect 6184 371288 6236 371340
rect 3700 353200 3752 353252
rect 17868 353200 17920 353252
rect 541256 353200 541308 353252
rect 558276 353200 558328 353252
rect 558184 351908 558236 351960
rect 580172 351908 580224 351960
rect 3516 346196 3568 346248
rect 7564 346196 7616 346248
rect 541992 342184 542044 342236
rect 580356 342184 580408 342236
rect 3792 329740 3844 329792
rect 17868 329740 17920 329792
rect 542268 329740 542320 329792
rect 580448 329740 580500 329792
rect 541716 325592 541768 325644
rect 580172 325592 580224 325644
rect 3332 318792 3384 318844
rect 17224 318792 17276 318844
rect 3884 306280 3936 306332
rect 17868 306280 17920 306332
rect 541900 306280 541952 306332
rect 580540 306280 580592 306332
rect 572076 298120 572128 298172
rect 579988 298120 580040 298172
rect 3516 293904 3568 293956
rect 17316 293904 17368 293956
rect 541348 293904 541400 293956
rect 580356 293904 580408 293956
rect 3976 282820 4028 282872
rect 16948 282820 17000 282872
rect 548524 273164 548576 273216
rect 579896 273164 579948 273216
rect 541716 259360 541768 259412
rect 579804 259360 579856 259412
rect 3608 258000 3660 258052
rect 17868 258000 17920 258052
rect 3700 246984 3752 247036
rect 16764 246984 16816 247036
rect 573456 244264 573508 244316
rect 580172 244264 580224 244316
rect 541624 233180 541676 233232
rect 580172 233180 580224 233232
rect 541992 219376 542044 219428
rect 579896 219376 579948 219428
rect 547144 193128 547196 193180
rect 580172 193128 580224 193180
rect 4804 187620 4856 187672
rect 17868 187620 17920 187672
rect 542268 187620 542320 187672
rect 556804 187620 556856 187672
rect 541900 179324 541952 179376
rect 580172 179324 580224 179376
rect 542268 175176 542320 175228
rect 573364 175176 573416 175228
rect 4896 164160 4948 164212
rect 17868 164160 17920 164212
rect 541992 164160 542044 164212
rect 571984 164160 572036 164212
rect 545764 153144 545816 153196
rect 580172 153144 580224 153196
rect 8944 139340 8996 139392
rect 16948 139340 17000 139392
rect 541808 139340 541860 139392
rect 580172 139340 580224 139392
rect 542268 139272 542320 139324
rect 580264 139272 580316 139324
rect 542268 128256 542320 128308
rect 556896 128256 556948 128308
rect 3424 115880 3476 115932
rect 17868 115880 17920 115932
rect 540980 115676 541032 115728
rect 543004 115676 543056 115728
rect 544384 113092 544436 113144
rect 580172 113092 580224 113144
rect 541716 100648 541768 100700
rect 579712 100648 579764 100700
rect 4988 92420 5040 92472
rect 17868 92420 17920 92472
rect 542268 92420 542320 92472
rect 558184 92420 558236 92472
rect 542268 79976 542320 80028
rect 572076 79976 572128 80028
rect 9036 68960 9088 69012
rect 17868 68960 17920 69012
rect 542268 68960 542320 69012
rect 573456 68960 573508 69012
rect 542268 56516 542320 56568
rect 580356 56516 580408 56568
rect 6184 45500 6236 45552
rect 16764 45500 16816 45552
rect 541900 45500 541952 45552
rect 580448 45500 580500 45552
rect 542268 33056 542320 33108
rect 580264 33056 580316 33108
rect 3884 22040 3936 22092
rect 17868 22040 17920 22092
rect 541992 22040 542044 22092
rect 580540 22040 580592 22092
rect 3424 13744 3476 13796
rect 55864 13744 55916 13796
rect 279332 13744 279384 13796
rect 580632 13744 580684 13796
rect 3516 13676 3568 13728
rect 427268 13676 427320 13728
rect 502156 13676 502208 13728
rect 580264 13676 580316 13728
rect 3608 13608 3660 13660
rect 352932 13608 352984 13660
rect 3700 13540 3752 13592
rect 204352 13540 204404 13592
rect 3792 13472 3844 13524
rect 130108 13472 130160 13524
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3436 614106 3464 658135
rect 3424 614100 3476 614106
rect 3424 614042 3476 614048
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 3436 590646 3464 606047
rect 3424 590640 3476 590646
rect 3424 590582 3476 590588
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3160 579834 3188 579935
rect 3148 579828 3200 579834
rect 3148 579770 3200 579776
rect 2964 554736 3016 554742
rect 2964 554678 3016 554684
rect 2976 553897 3004 554678
rect 2962 553888 3018 553897
rect 2962 553823 3018 553832
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3332 502308 3384 502314
rect 3332 502250 3384 502256
rect 3344 501809 3372 502250
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 2792 474978 2820 475623
rect 2780 474972 2832 474978
rect 2780 474914 2832 474920
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 2962 423600 3018 423609
rect 2962 423535 3018 423544
rect 2976 422346 3004 423535
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3146 371376 3202 371385
rect 3146 371311 3148 371320
rect 3200 371311 3202 371320
rect 3148 371282 3200 371288
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3436 115938 3464 527847
rect 3528 400178 3556 671191
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3516 400172 3568 400178
rect 3516 400114 3568 400120
rect 3516 398812 3568 398818
rect 3516 398754 3568 398760
rect 3528 397497 3556 398754
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3620 376718 3648 619103
rect 3698 566944 3754 566953
rect 3698 566879 3754 566888
rect 3608 376712 3660 376718
rect 3608 376654 3660 376660
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 3516 346248 3568 346254
rect 3516 346190 3568 346196
rect 3528 345409 3556 346190
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3516 293956 3568 293962
rect 3516 293898 3568 293904
rect 3528 293185 3556 293898
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3424 115932 3476 115938
rect 3424 115874 3476 115880
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3436 13802 3464 32399
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3528 13734 3556 267135
rect 3620 258058 3648 358391
rect 3712 353258 3740 566879
rect 3790 514856 3846 514865
rect 3790 514791 3846 514800
rect 3700 353252 3752 353258
rect 3700 353194 3752 353200
rect 3804 329798 3832 514791
rect 3882 462632 3938 462641
rect 3882 462567 3938 462576
rect 3792 329792 3844 329798
rect 3792 329734 3844 329740
rect 3896 306338 3924 462567
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 3884 306332 3936 306338
rect 3884 306274 3936 306280
rect 3698 306232 3754 306241
rect 3698 306167 3754 306176
rect 3608 258052 3660 258058
rect 3608 257994 3660 258000
rect 3712 247042 3740 306167
rect 3988 282878 4016 410479
rect 3976 282872 4028 282878
rect 3976 282814 4028 282820
rect 3700 247036 3752 247042
rect 3700 246978 3752 246984
rect 3606 214976 3662 214985
rect 3606 214911 3662 214920
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3620 13666 3648 214911
rect 4816 187678 4844 683674
rect 6932 657558 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 23492 657762 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40512 700330 40540 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 52460 700732 52512 700738
rect 52460 700674 52512 700680
rect 23572 700324 23624 700330
rect 23572 700266 23624 700272
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 23480 657756 23532 657762
rect 23480 657698 23532 657704
rect 6920 657552 6972 657558
rect 6920 657494 6972 657500
rect 23584 654922 23612 700266
rect 43444 657688 43496 657694
rect 43444 657630 43496 657636
rect 43456 654922 43484 657630
rect 23584 654894 23920 654922
rect 43148 654894 43484 654922
rect 52472 654922 52500 700674
rect 62120 700664 62172 700670
rect 62120 700606 62172 700612
rect 62132 654922 62160 700606
rect 71792 657626 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 81440 700596 81492 700602
rect 81440 700538 81492 700544
rect 71780 657620 71832 657626
rect 71780 657562 71832 657568
rect 81452 654922 81480 700538
rect 88352 657830 88380 702406
rect 100760 700528 100812 700534
rect 100760 700470 100812 700476
rect 88340 657824 88392 657830
rect 88340 657766 88392 657772
rect 100772 654922 100800 700470
rect 104912 657694 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 120080 700460 120132 700466
rect 120080 700402 120132 700408
rect 104900 657688 104952 657694
rect 104900 657630 104952 657636
rect 120092 654922 120120 700402
rect 136652 657694 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 139400 700392 139452 700398
rect 139400 700334 139452 700340
rect 136640 657688 136692 657694
rect 136640 657630 136692 657636
rect 139412 654922 139440 700334
rect 153212 657898 153240 702406
rect 170324 700738 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170312 700732 170364 700738
rect 170312 700674 170364 700680
rect 167000 700324 167052 700330
rect 167000 700266 167052 700272
rect 167012 673454 167040 700266
rect 167012 673426 167960 673454
rect 153200 657892 153252 657898
rect 153200 657834 153252 657840
rect 167932 654922 167960 673426
rect 201512 657762 201540 702986
rect 218072 657830 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 253940 700664 253992 700670
rect 253940 700606 253992 700612
rect 253952 673454 253980 700606
rect 267660 697610 267688 703520
rect 273260 700800 273312 700806
rect 273260 700742 273312 700748
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 253952 673426 254624 673454
rect 225788 657892 225840 657898
rect 225788 657834 225840 657840
rect 216128 657824 216180 657830
rect 216128 657766 216180 657772
rect 218060 657824 218112 657830
rect 218060 657766 218112 657772
rect 196900 657756 196952 657762
rect 196900 657698 196952 657704
rect 201500 657756 201552 657762
rect 201500 657698 201552 657704
rect 196912 654922 196940 657698
rect 216140 654922 216168 657766
rect 225800 654922 225828 657834
rect 235356 657824 235408 657830
rect 235356 657766 235408 657772
rect 235368 654922 235396 657766
rect 254596 654922 254624 673426
rect 266372 657830 266400 697546
rect 273272 673454 273300 700742
rect 283852 700670 283880 703520
rect 292580 700732 292632 700738
rect 292580 700674 292632 700680
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 292592 673454 292620 700674
rect 300136 700602 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 311900 700664 311952 700670
rect 311900 700606 311952 700612
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 311912 673454 311940 700606
rect 273272 673426 273852 673454
rect 292592 673426 293080 673454
rect 311912 673426 312400 673454
rect 266360 657824 266412 657830
rect 266360 657766 266412 657772
rect 273824 654922 273852 673426
rect 293052 654922 293080 673426
rect 312372 654922 312400 673426
rect 331232 657898 331260 702986
rect 348804 700806 348832 703520
rect 348792 700800 348844 700806
rect 348792 700742 348844 700748
rect 340880 700596 340932 700602
rect 340880 700538 340932 700544
rect 340892 673454 340920 700538
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 340892 673426 341288 673454
rect 331220 657892 331272 657898
rect 331220 657834 331272 657840
rect 341260 654922 341288 673426
rect 389456 657620 389508 657626
rect 389456 657562 389508 657568
rect 370228 657552 370280 657558
rect 370228 657494 370280 657500
rect 370240 654922 370268 657494
rect 389468 654922 389496 657562
rect 397472 657558 397500 703520
rect 413664 700738 413692 703520
rect 413652 700732 413704 700738
rect 413652 700674 413704 700680
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 447232 657892 447284 657898
rect 447232 657834 447284 657840
rect 428004 657824 428056 657830
rect 428004 657766 428056 657772
rect 408684 657756 408736 657762
rect 408684 657698 408736 657704
rect 399116 657688 399168 657694
rect 399116 657630 399168 657636
rect 397460 657552 397512 657558
rect 397460 657494 397512 657500
rect 399128 654922 399156 657630
rect 408696 654922 408724 657698
rect 428016 654922 428044 657766
rect 447244 654922 447272 657834
rect 462332 657626 462360 703520
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 494808 700398 494836 703520
rect 527192 700398 527220 703520
rect 543476 700602 543504 703520
rect 543464 700596 543516 700602
rect 543464 700538 543516 700544
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 514760 700392 514812 700398
rect 514760 700334 514812 700340
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 462320 657620 462372 657626
rect 462320 657562 462372 657568
rect 485780 657620 485832 657626
rect 485780 657562 485832 657568
rect 466460 657552 466512 657558
rect 466460 657494 466512 657500
rect 466472 654922 466500 657494
rect 485792 654922 485820 657562
rect 514772 654922 514800 700334
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 541624 696992 541676 696998
rect 541624 696934 541676 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 52472 654894 52808 654922
rect 62132 654894 62376 654922
rect 81452 654894 81696 654922
rect 100772 654894 100924 654922
rect 120092 654894 120152 654922
rect 139412 654894 139472 654922
rect 167932 654894 168360 654922
rect 196912 654894 197248 654922
rect 216140 654894 216476 654922
rect 225800 654894 226136 654922
rect 235368 654894 235704 654922
rect 254596 654894 255024 654922
rect 273824 654894 274252 654922
rect 293052 654894 293480 654922
rect 312372 654894 312800 654922
rect 341260 654894 341688 654922
rect 370240 654894 370576 654922
rect 389468 654894 389804 654922
rect 399128 654894 399464 654922
rect 408696 654894 409032 654922
rect 428016 654894 428352 654922
rect 447244 654894 447580 654922
rect 466472 654894 466808 654922
rect 485792 654894 486128 654922
rect 514772 654894 515016 654922
rect 4896 632120 4948 632126
rect 4896 632062 4948 632068
rect 4804 187672 4856 187678
rect 4804 187614 4856 187620
rect 4908 164218 4936 632062
rect 17040 614100 17092 614106
rect 17040 614042 17092 614048
rect 17052 613465 17080 614042
rect 541636 613465 541664 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 558184 683188 558236 683194
rect 558184 683130 558236 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 556804 670744 556856 670750
rect 556804 670686 556856 670692
rect 17038 613456 17094 613465
rect 17038 613391 17094 613400
rect 541622 613456 541678 613465
rect 541622 613391 541678 613400
rect 542268 601656 542320 601662
rect 542266 601624 542268 601633
rect 542320 601624 542322 601633
rect 542266 601559 542322 601568
rect 541808 590708 541860 590714
rect 541808 590650 541860 590656
rect 17868 590640 17920 590646
rect 17868 590582 17920 590588
rect 17880 589801 17908 590582
rect 541820 589801 541848 590650
rect 17866 589792 17922 589801
rect 17866 589727 17922 589736
rect 541806 589792 541862 589801
rect 541806 589727 541862 589736
rect 8944 579828 8996 579834
rect 8944 579770 8996 579776
rect 4988 474972 5040 474978
rect 4988 474914 5040 474920
rect 4896 164212 4948 164218
rect 4896 164154 4948 164160
rect 3698 162888 3754 162897
rect 3698 162823 3754 162832
rect 3608 13660 3660 13666
rect 3608 13602 3660 13608
rect 3712 13598 3740 162823
rect 3790 110664 3846 110673
rect 3790 110599 3846 110608
rect 3700 13592 3752 13598
rect 3700 13534 3752 13540
rect 3804 13530 3832 110599
rect 5000 92478 5028 474914
rect 7564 470620 7616 470626
rect 7564 470562 7616 470568
rect 6184 371340 6236 371346
rect 6184 371282 6236 371288
rect 4988 92472 5040 92478
rect 4988 92414 5040 92420
rect 3882 71632 3938 71641
rect 3882 71567 3938 71576
rect 3896 22098 3924 71567
rect 6196 45558 6224 371282
rect 7576 346254 7604 470562
rect 7564 346248 7616 346254
rect 7564 346190 7616 346196
rect 8956 139398 8984 579770
rect 17866 565992 17922 566001
rect 15844 565956 15896 565962
rect 17866 565927 17868 565936
rect 15844 565898 15896 565904
rect 17920 565927 17922 565936
rect 541714 565992 541770 566001
rect 541714 565927 541770 565936
rect 17868 565898 17920 565904
rect 15856 554742 15884 565898
rect 15844 554736 15896 554742
rect 15844 554678 15896 554684
rect 541622 554160 541678 554169
rect 541622 554095 541678 554104
rect 17222 542328 17278 542337
rect 17222 542263 17278 542272
rect 17236 502314 17264 542263
rect 17406 518664 17462 518673
rect 17406 518599 17462 518608
rect 17224 502308 17276 502314
rect 17224 502250 17276 502256
rect 17222 494864 17278 494873
rect 17222 494799 17278 494808
rect 9036 422340 9088 422346
rect 9036 422282 9088 422288
rect 8944 139392 8996 139398
rect 8944 139334 8996 139340
rect 9048 69018 9076 422282
rect 17236 398818 17264 494799
rect 17314 459368 17370 459377
rect 17314 459303 17370 459312
rect 17224 398812 17276 398818
rect 17224 398754 17276 398760
rect 16764 376712 16816 376718
rect 16764 376654 16816 376660
rect 16776 376417 16804 376654
rect 16762 376408 16818 376417
rect 16762 376343 16818 376352
rect 17224 318844 17276 318850
rect 17224 318786 17276 318792
rect 16948 282872 17000 282878
rect 16948 282814 17000 282820
rect 16960 281625 16988 282814
rect 16946 281616 17002 281625
rect 16946 281551 17002 281560
rect 16764 247036 16816 247042
rect 16764 246978 16816 246984
rect 16776 245993 16804 246978
rect 16762 245984 16818 245993
rect 16762 245919 16818 245928
rect 16948 139392 17000 139398
rect 16946 139360 16948 139369
rect 17000 139360 17002 139369
rect 16946 139295 17002 139304
rect 9036 69012 9088 69018
rect 9036 68954 9088 68960
rect 6184 45552 6236 45558
rect 6184 45494 6236 45500
rect 16764 45552 16816 45558
rect 16764 45494 16816 45500
rect 16776 44577 16804 45494
rect 16762 44568 16818 44577
rect 16762 44503 16818 44512
rect 17236 32745 17264 318786
rect 17328 293962 17356 459303
rect 17420 449886 17448 518599
rect 541636 485790 541664 554095
rect 541728 538218 541756 565927
rect 541898 542328 541954 542337
rect 541898 542263 541954 542272
rect 541716 538212 541768 538218
rect 541716 538154 541768 538160
rect 541806 518664 541862 518673
rect 541806 518599 541862 518608
rect 541714 506832 541770 506841
rect 541714 506767 541770 506776
rect 541624 485784 541676 485790
rect 541624 485726 541676 485732
rect 541622 483032 541678 483041
rect 541622 482967 541678 482976
rect 17866 471200 17922 471209
rect 17866 471135 17922 471144
rect 17880 470626 17908 471135
rect 17868 470620 17920 470626
rect 17868 470562 17920 470568
rect 17408 449880 17460 449886
rect 17408 449822 17460 449828
rect 541438 447536 541494 447545
rect 541438 447471 541494 447480
rect 541452 447370 541480 447471
rect 541440 447364 541492 447370
rect 541440 447306 541492 447312
rect 17868 400172 17920 400178
rect 17868 400114 17920 400120
rect 17880 400081 17908 400114
rect 17866 400072 17922 400081
rect 17866 400007 17922 400016
rect 17868 353252 17920 353258
rect 17868 353194 17920 353200
rect 541256 353252 541308 353258
rect 541256 353194 541308 353200
rect 17880 352753 17908 353194
rect 541268 352753 541296 353194
rect 17866 352744 17922 352753
rect 17866 352679 17922 352688
rect 541254 352744 541310 352753
rect 541254 352679 541310 352688
rect 17868 329792 17920 329798
rect 17868 329734 17920 329740
rect 17880 328953 17908 329734
rect 17866 328944 17922 328953
rect 17866 328879 17922 328888
rect 17868 306332 17920 306338
rect 17868 306274 17920 306280
rect 17880 305289 17908 306274
rect 17866 305280 17922 305289
rect 17866 305215 17922 305224
rect 17316 293956 17368 293962
rect 17316 293898 17368 293904
rect 541348 293956 541400 293962
rect 541348 293898 541400 293904
rect 541360 293457 541388 293898
rect 541346 293448 541402 293457
rect 541346 293383 541402 293392
rect 17868 258052 17920 258058
rect 17868 257994 17920 258000
rect 17880 257825 17908 257994
rect 17866 257816 17922 257825
rect 17866 257751 17922 257760
rect 541636 233238 541664 482967
rect 541728 325650 541756 506767
rect 541820 379506 541848 518599
rect 541912 431934 541940 542263
rect 542266 494864 542322 494873
rect 542266 494799 542322 494808
rect 542280 494154 542308 494799
rect 542268 494148 542320 494154
rect 542268 494090 542320 494096
rect 548524 494148 548576 494154
rect 548524 494090 548576 494096
rect 542266 471200 542322 471209
rect 542266 471135 542268 471144
rect 542320 471135 542322 471144
rect 547144 471164 547196 471170
rect 542268 471106 542320 471112
rect 547144 471106 547196 471112
rect 542174 459368 542230 459377
rect 542174 459303 542230 459312
rect 542188 458250 542216 459303
rect 542176 458244 542228 458250
rect 542176 458186 542228 458192
rect 545764 458244 545816 458250
rect 545764 458186 545816 458192
rect 544384 447364 544436 447370
rect 544384 447306 544436 447312
rect 541900 431928 541952 431934
rect 541900 431870 541952 431876
rect 543004 404388 543056 404394
rect 543004 404330 543056 404336
rect 542268 400172 542320 400178
rect 542268 400114 542320 400120
rect 542280 400081 542308 400114
rect 542266 400072 542322 400081
rect 542266 400007 542322 400016
rect 542268 389156 542320 389162
rect 542268 389098 542320 389104
rect 542280 388249 542308 389098
rect 542266 388240 542322 388249
rect 542266 388175 542322 388184
rect 541808 379500 541860 379506
rect 541808 379442 541860 379448
rect 541900 376712 541952 376718
rect 541900 376654 541952 376660
rect 541912 376417 541940 376654
rect 541898 376408 541954 376417
rect 541898 376343 541954 376352
rect 541992 342236 542044 342242
rect 541992 342178 542044 342184
rect 542004 340921 542032 342178
rect 541990 340912 542046 340921
rect 541990 340847 542046 340856
rect 542268 329792 542320 329798
rect 542268 329734 542320 329740
rect 542280 328953 542308 329734
rect 542266 328944 542322 328953
rect 542266 328879 542322 328888
rect 541716 325644 541768 325650
rect 541716 325586 541768 325592
rect 541900 306332 541952 306338
rect 541900 306274 541952 306280
rect 541912 305289 541940 306274
rect 541898 305280 541954 305289
rect 541898 305215 541954 305224
rect 541714 281616 541770 281625
rect 541714 281551 541770 281560
rect 541728 259418 541756 281551
rect 541990 269784 542046 269793
rect 541990 269719 542046 269728
rect 541716 259412 541768 259418
rect 541716 259354 541768 259360
rect 541898 257816 541954 257825
rect 541898 257751 541954 257760
rect 541806 245984 541862 245993
rect 541806 245919 541862 245928
rect 541714 234152 541770 234161
rect 541714 234087 541770 234096
rect 541624 233232 541676 233238
rect 541624 233174 541676 233180
rect 17868 187672 17920 187678
rect 17868 187614 17920 187620
rect 17880 186833 17908 187614
rect 17866 186824 17922 186833
rect 17866 186759 17922 186768
rect 17868 164212 17920 164218
rect 17868 164154 17920 164160
rect 17880 163033 17908 164154
rect 17866 163024 17922 163033
rect 17866 162959 17922 162968
rect 17868 115932 17920 115938
rect 17868 115874 17920 115880
rect 17880 115705 17908 115874
rect 540980 115728 541032 115734
rect 17866 115696 17922 115705
rect 17866 115631 17922 115640
rect 540978 115696 540980 115705
rect 541032 115696 541034 115705
rect 540978 115631 541034 115640
rect 541728 100706 541756 234087
rect 541820 139398 541848 245919
rect 541912 179382 541940 257751
rect 542004 219434 542032 269719
rect 541992 219428 542044 219434
rect 541992 219370 542044 219376
rect 542268 187672 542320 187678
rect 542268 187614 542320 187620
rect 542280 186833 542308 187614
rect 542266 186824 542322 186833
rect 542266 186759 542322 186768
rect 541900 179376 541952 179382
rect 541900 179318 541952 179324
rect 542268 175228 542320 175234
rect 542268 175170 542320 175176
rect 542280 174865 542308 175170
rect 542266 174856 542322 174865
rect 542266 174791 542322 174800
rect 541992 164212 542044 164218
rect 541992 164154 542044 164160
rect 542004 163033 542032 164154
rect 541990 163024 542046 163033
rect 541990 162959 542046 162968
rect 541808 139392 541860 139398
rect 541808 139334 541860 139340
rect 542266 139360 542322 139369
rect 542266 139295 542268 139304
rect 542320 139295 542322 139304
rect 542268 139266 542320 139272
rect 542268 128308 542320 128314
rect 542268 128250 542320 128256
rect 542280 127537 542308 128250
rect 542266 127528 542322 127537
rect 542266 127463 542322 127472
rect 543016 115734 543044 404330
rect 543004 115728 543056 115734
rect 543004 115670 543056 115676
rect 544396 113150 544424 447306
rect 545776 153202 545804 458186
rect 547156 193186 547184 471106
rect 548536 273222 548564 494090
rect 548524 273216 548576 273222
rect 548524 273158 548576 273164
rect 547144 193180 547196 193186
rect 547144 193122 547196 193128
rect 556816 187678 556844 670686
rect 556896 456816 556948 456822
rect 556896 456758 556948 456764
rect 556804 187672 556856 187678
rect 556804 187614 556856 187620
rect 545764 153196 545816 153202
rect 545764 153138 545816 153144
rect 556908 128314 556936 456758
rect 558196 400178 558224 683130
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 573456 630692 573508 630698
rect 573456 630634 573508 630640
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 573364 616888 573416 616894
rect 573364 616830 573416 616836
rect 572076 576904 572128 576910
rect 572076 576846 572128 576852
rect 571984 563100 572036 563106
rect 571984 563042 572036 563048
rect 558276 524476 558328 524482
rect 558276 524418 558328 524424
rect 558184 400172 558236 400178
rect 558184 400114 558236 400120
rect 558288 353258 558316 524418
rect 558276 353252 558328 353258
rect 558276 353194 558328 353200
rect 558184 351960 558236 351966
rect 558184 351902 558236 351908
rect 556896 128308 556948 128314
rect 556896 128250 556948 128256
rect 544384 113144 544436 113150
rect 544384 113086 544436 113092
rect 541716 100700 541768 100706
rect 541716 100642 541768 100648
rect 558196 92478 558224 351902
rect 571996 164218 572024 563042
rect 572088 376718 572116 576846
rect 572076 376712 572128 376718
rect 572076 376654 572128 376660
rect 572076 298172 572128 298178
rect 572076 298114 572128 298120
rect 571984 164212 572036 164218
rect 571984 164154 572036 164160
rect 17868 92472 17920 92478
rect 17868 92414 17920 92420
rect 542268 92472 542320 92478
rect 542268 92414 542320 92420
rect 558184 92472 558236 92478
rect 558184 92414 558236 92420
rect 17880 91905 17908 92414
rect 542280 91905 542308 92414
rect 17866 91896 17922 91905
rect 17866 91831 17922 91840
rect 542266 91896 542322 91905
rect 542266 91831 542322 91840
rect 542266 80064 542322 80073
rect 572088 80034 572116 298114
rect 573376 175234 573404 616830
rect 573468 389162 573496 630634
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580276 601662 580304 643991
rect 580264 601656 580316 601662
rect 580264 601598 580316 601604
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580262 511320 580318 511329
rect 580262 511255 580318 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579620 431928 579672 431934
rect 579620 431870 579672 431876
rect 579632 431633 579660 431870
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 573456 389156 573508 389162
rect 573456 389098 573508 389104
rect 579804 379500 579856 379506
rect 579804 379442 579856 379448
rect 579816 378457 579844 379442
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 579986 298752 580042 298761
rect 579986 298687 580042 298696
rect 580000 298178 580028 298687
rect 579988 298172 580040 298178
rect 579988 298114 580040 298120
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 573456 244316 573508 244322
rect 573456 244258 573508 244264
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 573364 175228 573416 175234
rect 573364 175170 573416 175176
rect 542266 79999 542268 80008
rect 542320 79999 542322 80008
rect 572076 80028 572128 80034
rect 542268 79970 542320 79976
rect 572076 79970 572128 79976
rect 573468 69018 573496 244258
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580276 139330 580304 511255
rect 580354 471472 580410 471481
rect 580354 471407 580410 471416
rect 580368 342242 580396 471407
rect 580446 418296 580502 418305
rect 580446 418231 580502 418240
rect 580356 342236 580408 342242
rect 580356 342178 580408 342184
rect 580460 329798 580488 418231
rect 580538 365120 580594 365129
rect 580538 365055 580594 365064
rect 580448 329792 580500 329798
rect 580448 329734 580500 329740
rect 580354 312080 580410 312089
rect 580354 312015 580410 312024
rect 580368 293962 580396 312015
rect 580552 306338 580580 365055
rect 580540 306332 580592 306338
rect 580540 306274 580592 306280
rect 580356 293956 580408 293962
rect 580356 293898 580408 293904
rect 580354 205728 580410 205737
rect 580354 205663 580410 205672
rect 580170 139295 580226 139304
rect 580264 139324 580316 139330
rect 580264 139266 580316 139272
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 579712 100700 579764 100706
rect 579712 100642 579764 100648
rect 579724 99521 579752 100642
rect 579710 99512 579766 99521
rect 579710 99447 579766 99456
rect 17868 69012 17920 69018
rect 17868 68954 17920 68960
rect 542268 69012 542320 69018
rect 542268 68954 542320 68960
rect 573456 69012 573508 69018
rect 573456 68954 573508 68960
rect 17880 68241 17908 68954
rect 542280 68241 542308 68954
rect 17866 68232 17922 68241
rect 17866 68167 17922 68176
rect 542266 68232 542322 68241
rect 542266 68167 542322 68176
rect 542268 56568 542320 56574
rect 542268 56510 542320 56516
rect 542280 56409 542308 56510
rect 542266 56400 542322 56409
rect 542266 56335 542322 56344
rect 541900 45552 541952 45558
rect 541900 45494 541952 45500
rect 541912 44577 541940 45494
rect 541898 44568 541954 44577
rect 541898 44503 541954 44512
rect 580276 33114 580304 125967
rect 580368 56574 580396 205663
rect 580446 165880 580502 165889
rect 580446 165815 580502 165824
rect 580356 56568 580408 56574
rect 580356 56510 580408 56516
rect 580460 45558 580488 165815
rect 580538 86184 580594 86193
rect 580538 86119 580594 86128
rect 580448 45552 580500 45558
rect 580448 45494 580500 45500
rect 542268 33108 542320 33114
rect 542268 33050 542320 33056
rect 580264 33108 580316 33114
rect 580264 33050 580316 33056
rect 542280 32745 542308 33050
rect 17222 32736 17278 32745
rect 17222 32671 17278 32680
rect 542266 32736 542322 32745
rect 542266 32671 542322 32680
rect 580552 22098 580580 86119
rect 580630 59664 580686 59673
rect 580630 59599 580686 59608
rect 3884 22092 3936 22098
rect 3884 22034 3936 22040
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 541992 22092 542044 22098
rect 541992 22034 542044 22040
rect 580540 22092 580592 22098
rect 580540 22034 580592 22040
rect 17880 20913 17908 22034
rect 542004 20913 542032 22034
rect 17866 20904 17922 20913
rect 17866 20839 17922 20848
rect 541990 20904 542046 20913
rect 541990 20839 542046 20848
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 55876 15014 56212 15042
rect 130120 15014 130456 15042
rect 204364 15014 204700 15042
rect 279036 15014 279372 15042
rect 55876 13802 55904 15014
rect 55864 13796 55916 13802
rect 55864 13738 55916 13744
rect 130120 13530 130148 15014
rect 204364 13598 204392 15014
rect 279344 13802 279372 15014
rect 352944 15014 353280 15042
rect 427280 15014 427616 15042
rect 501860 15014 502196 15042
rect 279332 13796 279384 13802
rect 279332 13738 279384 13744
rect 352944 13666 352972 15014
rect 427280 13734 427308 15014
rect 502168 13734 502196 15014
rect 580276 13734 580304 19751
rect 580644 13802 580672 59599
rect 580632 13796 580684 13802
rect 580632 13738 580684 13744
rect 427268 13728 427320 13734
rect 427268 13670 427320 13676
rect 502156 13728 502208 13734
rect 502156 13670 502208 13676
rect 580264 13728 580316 13734
rect 580264 13670 580316 13676
rect 352932 13660 352984 13666
rect 352932 13602 352984 13608
rect 204352 13592 204404 13598
rect 204352 13534 204404 13540
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 130108 13524 130160 13530
rect 130108 13466 130160 13472
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3422 606056 3478 606112
rect 3146 579944 3202 580000
rect 2962 553832 3018 553888
rect 3422 527856 3478 527912
rect 3330 501744 3386 501800
rect 2778 475632 2834 475688
rect 3330 449520 3386 449576
rect 2962 423544 3018 423600
rect 3146 371340 3202 371376
rect 3146 371320 3148 371340
rect 3148 371320 3200 371340
rect 3200 371320 3202 371340
rect 3330 319232 3386 319288
rect 3606 619112 3662 619168
rect 3514 397432 3570 397488
rect 3698 566888 3754 566944
rect 3606 358400 3662 358456
rect 3514 345344 3570 345400
rect 3514 293120 3570 293176
rect 3514 267144 3570 267200
rect 3422 32408 3478 32464
rect 3790 514800 3846 514856
rect 3882 462576 3938 462632
rect 3974 410488 4030 410544
rect 3698 306176 3754 306232
rect 3606 214920 3662 214976
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 17038 613400 17094 613456
rect 541622 613400 541678 613456
rect 542266 601604 542268 601624
rect 542268 601604 542320 601624
rect 542320 601604 542322 601624
rect 542266 601568 542322 601604
rect 17866 589736 17922 589792
rect 541806 589736 541862 589792
rect 3698 162832 3754 162888
rect 3790 110608 3846 110664
rect 3882 71576 3938 71632
rect 17866 565956 17922 565992
rect 17866 565936 17868 565956
rect 17868 565936 17920 565956
rect 17920 565936 17922 565956
rect 541714 565936 541770 565992
rect 541622 554104 541678 554160
rect 17222 542272 17278 542328
rect 17406 518608 17462 518664
rect 17222 494808 17278 494864
rect 17314 459312 17370 459368
rect 16762 376352 16818 376408
rect 16946 281560 17002 281616
rect 16762 245928 16818 245984
rect 16946 139340 16948 139360
rect 16948 139340 17000 139360
rect 17000 139340 17002 139360
rect 16946 139304 17002 139340
rect 16762 44512 16818 44568
rect 541898 542272 541954 542328
rect 541806 518608 541862 518664
rect 541714 506776 541770 506832
rect 541622 482976 541678 483032
rect 17866 471144 17922 471200
rect 541438 447480 541494 447536
rect 17866 400016 17922 400072
rect 17866 352688 17922 352744
rect 541254 352688 541310 352744
rect 17866 328888 17922 328944
rect 17866 305224 17922 305280
rect 541346 293392 541402 293448
rect 17866 257760 17922 257816
rect 542266 494808 542322 494864
rect 542266 471164 542322 471200
rect 542266 471144 542268 471164
rect 542268 471144 542320 471164
rect 542320 471144 542322 471164
rect 542174 459312 542230 459368
rect 542266 400016 542322 400072
rect 542266 388184 542322 388240
rect 541898 376352 541954 376408
rect 541990 340856 542046 340912
rect 542266 328888 542322 328944
rect 541898 305224 541954 305280
rect 541714 281560 541770 281616
rect 541990 269728 542046 269784
rect 541898 257760 541954 257816
rect 541806 245928 541862 245984
rect 541714 234096 541770 234152
rect 17866 186768 17922 186824
rect 17866 162968 17922 163024
rect 17866 115640 17922 115696
rect 540978 115676 540980 115696
rect 540980 115676 541032 115696
rect 541032 115676 541034 115696
rect 540978 115640 541034 115676
rect 542266 186768 542322 186824
rect 542266 174800 542322 174856
rect 541990 162968 542046 163024
rect 542266 139324 542322 139360
rect 542266 139304 542268 139324
rect 542268 139304 542320 139324
rect 542320 139304 542322 139324
rect 542266 127472 542322 127528
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580262 644000 580318 644056
rect 579986 630808 580042 630864
rect 17866 91840 17922 91896
rect 542266 91840 542322 91896
rect 542266 80028 542322 80064
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580262 511264 580318 511320
rect 580170 484608 580226 484664
rect 580170 458088 580226 458144
rect 579618 431568 579674 431624
rect 580170 404912 580226 404968
rect 579802 378392 579858 378448
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 298696 580042 298752
rect 579894 272176 579950 272232
rect 579802 258848 579858 258904
rect 580170 245520 580226 245576
rect 542266 80008 542268 80028
rect 542268 80008 542320 80028
rect 542320 80008 542322 80028
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580354 471416 580410 471472
rect 580446 418240 580502 418296
rect 580538 365064 580594 365120
rect 580354 312024 580410 312080
rect 580354 205672 580410 205728
rect 580262 125976 580318 126032
rect 580170 112784 580226 112840
rect 579710 99456 579766 99512
rect 17866 68176 17922 68232
rect 542266 68176 542322 68232
rect 542266 56344 542322 56400
rect 541898 44512 541954 44568
rect 580446 165824 580502 165880
rect 580538 86128 580594 86184
rect 17222 32680 17278 32736
rect 542266 32680 542322 32736
rect 580630 59608 580686 59664
rect 17866 20848 17922 20904
rect 541990 20848 542046 20904
rect 580262 19760 580318 19816
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 17033 613458 17099 613461
rect 541617 613458 541683 613461
rect 17033 613456 19228 613458
rect 17033 613400 17038 613456
rect 17094 613400 19228 613456
rect 17033 613398 19228 613400
rect 539028 613456 541683 613458
rect 539028 613400 541622 613456
rect 541678 613400 541683 613456
rect 539028 613398 541683 613400
rect 17033 613395 17099 613398
rect 541617 613395 541683 613398
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect 542261 601626 542327 601629
rect 539028 601624 542327 601626
rect 539028 601568 542266 601624
rect 542322 601568 542327 601624
rect 539028 601566 542327 601568
rect 542261 601563 542327 601566
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 17861 589794 17927 589797
rect 541801 589794 541867 589797
rect 17861 589792 19228 589794
rect 17861 589736 17866 589792
rect 17922 589736 19228 589792
rect 17861 589734 19228 589736
rect 539028 589792 541867 589794
rect 539028 589736 541806 589792
rect 541862 589736 541867 589792
rect 539028 589734 541867 589736
rect 17861 589731 17927 589734
rect 541801 589731 541867 589734
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3693 566946 3759 566949
rect -960 566944 3759 566946
rect -960 566888 3698 566944
rect 3754 566888 3759 566944
rect -960 566886 3759 566888
rect -960 566796 480 566886
rect 3693 566883 3759 566886
rect 17861 565994 17927 565997
rect 541709 565994 541775 565997
rect 17861 565992 19228 565994
rect 17861 565936 17866 565992
rect 17922 565936 19228 565992
rect 17861 565934 19228 565936
rect 539028 565992 541775 565994
rect 539028 565936 541714 565992
rect 541770 565936 541775 565992
rect 539028 565934 541775 565936
rect 17861 565931 17927 565934
rect 541709 565931 541775 565934
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 541617 554162 541683 554165
rect 539028 554160 541683 554162
rect 539028 554104 541622 554160
rect 541678 554104 541683 554160
rect 539028 554102 541683 554104
rect 541617 554099 541683 554102
rect -960 553890 480 553980
rect 2957 553890 3023 553893
rect -960 553888 3023 553890
rect -960 553832 2962 553888
rect 3018 553832 3023 553888
rect -960 553830 3023 553832
rect -960 553740 480 553830
rect 2957 553827 3023 553830
rect 583520 551020 584960 551260
rect 17217 542330 17283 542333
rect 541893 542330 541959 542333
rect 17217 542328 19228 542330
rect 17217 542272 17222 542328
rect 17278 542272 19228 542328
rect 17217 542270 19228 542272
rect 539028 542328 541959 542330
rect 539028 542272 541898 542328
rect 541954 542272 541959 542328
rect 539028 542270 541959 542272
rect 17217 542267 17283 542270
rect 541893 542267 541959 542270
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 17401 518666 17467 518669
rect 541801 518666 541867 518669
rect 17401 518664 19228 518666
rect 17401 518608 17406 518664
rect 17462 518608 19228 518664
rect 17401 518606 19228 518608
rect 539028 518664 541867 518666
rect 539028 518608 541806 518664
rect 541862 518608 541867 518664
rect 539028 518606 541867 518608
rect 17401 518603 17467 518606
rect 541801 518603 541867 518606
rect -960 514858 480 514948
rect 3785 514858 3851 514861
rect -960 514856 3851 514858
rect -960 514800 3790 514856
rect 3846 514800 3851 514856
rect -960 514798 3851 514800
rect -960 514708 480 514798
rect 3785 514795 3851 514798
rect 580257 511322 580323 511325
rect 583520 511322 584960 511412
rect 580257 511320 584960 511322
rect 580257 511264 580262 511320
rect 580318 511264 584960 511320
rect 580257 511262 584960 511264
rect 580257 511259 580323 511262
rect 583520 511172 584960 511262
rect 541709 506834 541775 506837
rect 539028 506832 541775 506834
rect 539028 506776 541714 506832
rect 541770 506776 541775 506832
rect 539028 506774 541775 506776
rect 541709 506771 541775 506774
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect 17217 494866 17283 494869
rect 542261 494866 542327 494869
rect 17217 494864 19228 494866
rect 17217 494808 17222 494864
rect 17278 494808 19228 494864
rect 17217 494806 19228 494808
rect 539028 494864 542327 494866
rect 539028 494808 542266 494864
rect 542322 494808 542327 494864
rect 539028 494806 542327 494808
rect 17217 494803 17283 494806
rect 542261 494803 542327 494806
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 541617 483034 541683 483037
rect 539028 483032 541683 483034
rect 539028 482976 541622 483032
rect 541678 482976 541683 483032
rect 539028 482974 541683 482976
rect 541617 482971 541683 482974
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 580349 471474 580415 471477
rect 583520 471474 584960 471564
rect 580349 471472 584960 471474
rect 580349 471416 580354 471472
rect 580410 471416 584960 471472
rect 580349 471414 584960 471416
rect 580349 471411 580415 471414
rect 583520 471324 584960 471414
rect 17861 471202 17927 471205
rect 542261 471202 542327 471205
rect 17861 471200 19228 471202
rect 17861 471144 17866 471200
rect 17922 471144 19228 471200
rect 17861 471142 19228 471144
rect 539028 471200 542327 471202
rect 539028 471144 542266 471200
rect 542322 471144 542327 471200
rect 539028 471142 542327 471144
rect 17861 471139 17927 471142
rect 542261 471139 542327 471142
rect -960 462634 480 462724
rect 3877 462634 3943 462637
rect -960 462632 3943 462634
rect -960 462576 3882 462632
rect 3938 462576 3943 462632
rect -960 462574 3943 462576
rect -960 462484 480 462574
rect 3877 462571 3943 462574
rect 17309 459370 17375 459373
rect 542169 459370 542235 459373
rect 17309 459368 19228 459370
rect 17309 459312 17314 459368
rect 17370 459312 19228 459368
rect 17309 459310 19228 459312
rect 539028 459368 542235 459370
rect 539028 459312 542174 459368
rect 542230 459312 542235 459368
rect 539028 459310 542235 459312
rect 17309 459307 17375 459310
rect 542169 459307 542235 459310
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 541433 447538 541499 447541
rect 539028 447536 541499 447538
rect 539028 447480 541438 447536
rect 541494 447480 541499 447536
rect 539028 447478 541499 447480
rect 541433 447475 541499 447478
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2957 423602 3023 423605
rect -960 423600 3023 423602
rect -960 423544 2962 423600
rect 3018 423544 3023 423600
rect -960 423542 3023 423544
rect -960 423452 480 423542
rect 2957 423539 3023 423542
rect 580441 418298 580507 418301
rect 583520 418298 584960 418388
rect 580441 418296 584960 418298
rect 580441 418240 580446 418296
rect 580502 418240 584960 418296
rect 580441 418238 584960 418240
rect 580441 418235 580507 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 17861 400074 17927 400077
rect 542261 400074 542327 400077
rect 17861 400072 19228 400074
rect 17861 400016 17866 400072
rect 17922 400016 19228 400072
rect 17861 400014 19228 400016
rect 539028 400072 542327 400074
rect 539028 400016 542266 400072
rect 542322 400016 542327 400072
rect 539028 400014 542327 400016
rect 17861 400011 17927 400014
rect 542261 400011 542327 400014
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect 542261 388242 542327 388245
rect 539028 388240 542327 388242
rect 539028 388184 542266 388240
rect 542322 388184 542327 388240
rect 539028 388182 542327 388184
rect 542261 388179 542327 388182
rect -960 384284 480 384524
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect 16757 376410 16823 376413
rect 541893 376410 541959 376413
rect 16757 376408 19228 376410
rect 16757 376352 16762 376408
rect 16818 376352 19228 376408
rect 16757 376350 19228 376352
rect 539028 376408 541959 376410
rect 539028 376352 541898 376408
rect 541954 376352 541959 376408
rect 539028 376350 541959 376352
rect 16757 376347 16823 376350
rect 541893 376347 541959 376350
rect -960 371378 480 371468
rect 3141 371378 3207 371381
rect -960 371376 3207 371378
rect -960 371320 3146 371376
rect 3202 371320 3207 371376
rect -960 371318 3207 371320
rect -960 371228 480 371318
rect 3141 371315 3207 371318
rect 580533 365122 580599 365125
rect 583520 365122 584960 365212
rect 580533 365120 584960 365122
rect 580533 365064 580538 365120
rect 580594 365064 584960 365120
rect 580533 365062 584960 365064
rect 580533 365059 580599 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 17861 352746 17927 352749
rect 541249 352746 541315 352749
rect 17861 352744 19228 352746
rect 17861 352688 17866 352744
rect 17922 352688 19228 352744
rect 17861 352686 19228 352688
rect 539028 352744 541315 352746
rect 539028 352688 541254 352744
rect 541310 352688 541315 352744
rect 539028 352686 541315 352688
rect 17861 352683 17927 352686
rect 541249 352683 541315 352686
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 541985 340914 542051 340917
rect 539028 340912 542051 340914
rect 539028 340856 541990 340912
rect 542046 340856 542051 340912
rect 539028 340854 542051 340856
rect 541985 340851 542051 340854
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 17861 328946 17927 328949
rect 542261 328946 542327 328949
rect 17861 328944 19228 328946
rect 17861 328888 17866 328944
rect 17922 328888 19228 328944
rect 17861 328886 19228 328888
rect 539028 328944 542327 328946
rect 539028 328888 542266 328944
rect 542322 328888 542327 328944
rect 539028 328886 542327 328888
rect 17861 328883 17927 328886
rect 542261 328883 542327 328886
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580349 312082 580415 312085
rect 583520 312082 584960 312172
rect 580349 312080 584960 312082
rect 580349 312024 580354 312080
rect 580410 312024 584960 312080
rect 580349 312022 584960 312024
rect 580349 312019 580415 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3693 306234 3759 306237
rect -960 306232 3759 306234
rect -960 306176 3698 306232
rect 3754 306176 3759 306232
rect -960 306174 3759 306176
rect -960 306084 480 306174
rect 3693 306171 3759 306174
rect 17861 305282 17927 305285
rect 541893 305282 541959 305285
rect 17861 305280 19228 305282
rect 17861 305224 17866 305280
rect 17922 305224 19228 305280
rect 17861 305222 19228 305224
rect 539028 305280 541959 305282
rect 539028 305224 541898 305280
rect 541954 305224 541959 305280
rect 539028 305222 541959 305224
rect 17861 305219 17927 305222
rect 541893 305219 541959 305222
rect 579981 298754 580047 298757
rect 583520 298754 584960 298844
rect 579981 298752 584960 298754
rect 579981 298696 579986 298752
rect 580042 298696 584960 298752
rect 579981 298694 584960 298696
rect 579981 298691 580047 298694
rect 583520 298604 584960 298694
rect 541341 293450 541407 293453
rect 539028 293448 541407 293450
rect 539028 293392 541346 293448
rect 541402 293392 541407 293448
rect 539028 293390 541407 293392
rect 541341 293387 541407 293390
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect 16941 281618 17007 281621
rect 541709 281618 541775 281621
rect 16941 281616 19228 281618
rect 16941 281560 16946 281616
rect 17002 281560 19228 281616
rect 16941 281558 19228 281560
rect 539028 281616 541775 281618
rect 539028 281560 541714 281616
rect 541770 281560 541775 281616
rect 539028 281558 541775 281560
rect 16941 281555 17007 281558
rect 541709 281555 541775 281558
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect 541985 269786 542051 269789
rect 539028 269784 542051 269786
rect 539028 269728 541990 269784
rect 542046 269728 542051 269784
rect 539028 269726 542051 269728
rect 541985 269723 542051 269726
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect 17861 257818 17927 257821
rect 541893 257818 541959 257821
rect 17861 257816 19228 257818
rect 17861 257760 17866 257816
rect 17922 257760 19228 257816
rect 17861 257758 19228 257760
rect 539028 257816 541959 257818
rect 539028 257760 541898 257816
rect 541954 257760 541959 257816
rect 539028 257758 541959 257760
rect 17861 257755 17927 257758
rect 541893 257755 541959 257758
rect -960 253996 480 254236
rect 16757 245986 16823 245989
rect 541801 245986 541867 245989
rect 16757 245984 19228 245986
rect 16757 245928 16762 245984
rect 16818 245928 19228 245984
rect 16757 245926 19228 245928
rect 539028 245984 541867 245986
rect 539028 245928 541806 245984
rect 541862 245928 541867 245984
rect 539028 245926 541867 245928
rect 16757 245923 16823 245926
rect 541801 245923 541867 245926
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 240940 480 241180
rect 541709 234154 541775 234157
rect 539028 234152 541775 234154
rect 539028 234096 541714 234152
rect 541770 234096 541775 234152
rect 539028 234094 541775 234096
rect 541709 234091 541775 234094
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3601 214978 3667 214981
rect -960 214976 3667 214978
rect -960 214920 3606 214976
rect 3662 214920 3667 214976
rect -960 214918 3667 214920
rect -960 214828 480 214918
rect 3601 214915 3667 214918
rect 580349 205730 580415 205733
rect 583520 205730 584960 205820
rect 580349 205728 584960 205730
rect 580349 205672 580354 205728
rect 580410 205672 584960 205728
rect 580349 205670 584960 205672
rect 580349 205667 580415 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 17861 186826 17927 186829
rect 542261 186826 542327 186829
rect 17861 186824 19228 186826
rect 17861 186768 17866 186824
rect 17922 186768 19228 186824
rect 17861 186766 19228 186768
rect 539028 186824 542327 186826
rect 539028 186768 542266 186824
rect 542322 186768 542327 186824
rect 539028 186766 542327 186768
rect 17861 186763 17927 186766
rect 542261 186763 542327 186766
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 542261 174858 542327 174861
rect 539028 174856 542327 174858
rect 539028 174800 542266 174856
rect 542322 174800 542327 174856
rect 539028 174798 542327 174800
rect 542261 174795 542327 174798
rect 580441 165882 580507 165885
rect 583520 165882 584960 165972
rect 580441 165880 584960 165882
rect 580441 165824 580446 165880
rect 580502 165824 584960 165880
rect 580441 165822 584960 165824
rect 580441 165819 580507 165822
rect 583520 165732 584960 165822
rect 17861 163026 17927 163029
rect 541985 163026 542051 163029
rect 17861 163024 19228 163026
rect -960 162890 480 162980
rect 17861 162968 17866 163024
rect 17922 162968 19228 163024
rect 17861 162966 19228 162968
rect 539028 163024 542051 163026
rect 539028 162968 541990 163024
rect 542046 162968 542051 163024
rect 539028 162966 542051 162968
rect 17861 162963 17927 162966
rect 541985 162963 542051 162966
rect 3693 162890 3759 162893
rect -960 162888 3759 162890
rect -960 162832 3698 162888
rect 3754 162832 3759 162888
rect -960 162830 3759 162832
rect -960 162740 480 162830
rect 3693 162827 3759 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149684 480 149924
rect 16941 139362 17007 139365
rect 542261 139362 542327 139365
rect 16941 139360 19228 139362
rect 16941 139304 16946 139360
rect 17002 139304 19228 139360
rect 16941 139302 19228 139304
rect 539028 139360 542327 139362
rect 539028 139304 542266 139360
rect 542322 139304 542327 139360
rect 539028 139302 542327 139304
rect 16941 139299 17007 139302
rect 542261 139299 542327 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136628 480 136868
rect 542261 127530 542327 127533
rect 539028 127528 542327 127530
rect 539028 127472 542266 127528
rect 542322 127472 542327 127528
rect 539028 127470 542327 127472
rect 542261 127467 542327 127470
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 580257 125971 580323 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 17861 115698 17927 115701
rect 540973 115698 541039 115701
rect 17861 115696 19228 115698
rect 17861 115640 17866 115696
rect 17922 115640 19228 115696
rect 17861 115638 19228 115640
rect 539028 115696 541039 115698
rect 539028 115640 540978 115696
rect 541034 115640 541039 115696
rect 539028 115638 541039 115640
rect 17861 115635 17927 115638
rect 540973 115635 541039 115638
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3785 110666 3851 110669
rect -960 110664 3851 110666
rect -960 110608 3790 110664
rect 3846 110608 3851 110664
rect -960 110606 3851 110608
rect -960 110516 480 110606
rect 3785 110603 3851 110606
rect 579705 99514 579771 99517
rect 583520 99514 584960 99604
rect 579705 99512 584960 99514
rect 579705 99456 579710 99512
rect 579766 99456 584960 99512
rect 579705 99454 584960 99456
rect 579705 99451 579771 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 17861 91898 17927 91901
rect 542261 91898 542327 91901
rect 17861 91896 19228 91898
rect 17861 91840 17866 91896
rect 17922 91840 19228 91896
rect 17861 91838 19228 91840
rect 539028 91896 542327 91898
rect 539028 91840 542266 91896
rect 542322 91840 542327 91896
rect 539028 91838 542327 91840
rect 17861 91835 17927 91838
rect 542261 91835 542327 91838
rect 580533 86186 580599 86189
rect 583520 86186 584960 86276
rect 580533 86184 584960 86186
rect 580533 86128 580538 86184
rect 580594 86128 584960 86184
rect 580533 86126 584960 86128
rect 580533 86123 580599 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 542261 80066 542327 80069
rect 539028 80064 542327 80066
rect 539028 80008 542266 80064
rect 542322 80008 542327 80064
rect 539028 80006 542327 80008
rect 542261 80003 542327 80006
rect 583520 72844 584960 73084
rect -960 71634 480 71724
rect 3877 71634 3943 71637
rect -960 71632 3943 71634
rect -960 71576 3882 71632
rect 3938 71576 3943 71632
rect -960 71574 3943 71576
rect -960 71484 480 71574
rect 3877 71571 3943 71574
rect 17861 68234 17927 68237
rect 542261 68234 542327 68237
rect 17861 68232 19228 68234
rect 17861 68176 17866 68232
rect 17922 68176 19228 68232
rect 17861 68174 19228 68176
rect 539028 68232 542327 68234
rect 539028 68176 542266 68232
rect 542322 68176 542327 68232
rect 539028 68174 542327 68176
rect 17861 68171 17927 68174
rect 542261 68171 542327 68174
rect 580625 59666 580691 59669
rect 583520 59666 584960 59756
rect 580625 59664 584960 59666
rect 580625 59608 580630 59664
rect 580686 59608 584960 59664
rect 580625 59606 584960 59608
rect 580625 59603 580691 59606
rect 583520 59516 584960 59606
rect -960 58428 480 58668
rect 542261 56402 542327 56405
rect 539028 56400 542327 56402
rect 539028 56344 542266 56400
rect 542322 56344 542327 56400
rect 539028 56342 542327 56344
rect 542261 56339 542327 56342
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 16757 44570 16823 44573
rect 541893 44570 541959 44573
rect 16757 44568 19228 44570
rect 16757 44512 16762 44568
rect 16818 44512 19228 44568
rect 16757 44510 19228 44512
rect 539028 44568 541959 44570
rect 539028 44512 541898 44568
rect 541954 44512 541959 44568
rect 539028 44510 541959 44512
rect 16757 44507 16823 44510
rect 541893 44507 541959 44510
rect 583520 32996 584960 33236
rect 17217 32738 17283 32741
rect 542261 32738 542327 32741
rect 17217 32736 19228 32738
rect 17217 32680 17222 32736
rect 17278 32680 19228 32736
rect 17217 32678 19228 32680
rect 539028 32736 542327 32738
rect 539028 32680 542266 32736
rect 542322 32680 542327 32736
rect 539028 32678 542327 32680
rect 17217 32675 17283 32678
rect 542261 32675 542327 32678
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 17861 20906 17927 20909
rect 541985 20906 542051 20909
rect 17861 20904 19228 20906
rect 17861 20848 17866 20904
rect 17922 20848 19228 20904
rect 17861 20846 19228 20848
rect 539028 20904 542051 20906
rect 539028 20848 541990 20904
rect 542046 20848 542051 20904
rect 539028 20846 542051 20848
rect 17861 20843 17927 20846
rect 541985 20843 542051 20846
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 6914 705798 7534 705830
rect 6914 705562 6946 705798
rect 7182 705562 7266 705798
rect 7502 705562 7534 705798
rect 6914 705478 7534 705562
rect 6914 705242 6946 705478
rect 7182 705242 7266 705478
rect 7502 705242 7534 705478
rect 6914 669454 7534 705242
rect 6914 669218 6946 669454
rect 7182 669218 7266 669454
rect 7502 669218 7534 669454
rect 6914 669134 7534 669218
rect 6914 668898 6946 669134
rect 7182 668898 7266 669134
rect 7502 668898 7534 669134
rect 6914 633454 7534 668898
rect 6914 633218 6946 633454
rect 7182 633218 7266 633454
rect 7502 633218 7534 633454
rect 6914 633134 7534 633218
rect 6914 632898 6946 633134
rect 7182 632898 7266 633134
rect 7502 632898 7534 633134
rect 6914 597454 7534 632898
rect 6914 597218 6946 597454
rect 7182 597218 7266 597454
rect 7502 597218 7534 597454
rect 6914 597134 7534 597218
rect 6914 596898 6946 597134
rect 7182 596898 7266 597134
rect 7502 596898 7534 597134
rect 6914 561454 7534 596898
rect 6914 561218 6946 561454
rect 7182 561218 7266 561454
rect 7502 561218 7534 561454
rect 6914 561134 7534 561218
rect 6914 560898 6946 561134
rect 7182 560898 7266 561134
rect 7502 560898 7534 561134
rect 6914 525454 7534 560898
rect 6914 525218 6946 525454
rect 7182 525218 7266 525454
rect 7502 525218 7534 525454
rect 6914 525134 7534 525218
rect 6914 524898 6946 525134
rect 7182 524898 7266 525134
rect 7502 524898 7534 525134
rect 6914 489454 7534 524898
rect 6914 489218 6946 489454
rect 7182 489218 7266 489454
rect 7502 489218 7534 489454
rect 6914 489134 7534 489218
rect 6914 488898 6946 489134
rect 7182 488898 7266 489134
rect 7502 488898 7534 489134
rect 6914 453454 7534 488898
rect 6914 453218 6946 453454
rect 7182 453218 7266 453454
rect 7502 453218 7534 453454
rect 6914 453134 7534 453218
rect 6914 452898 6946 453134
rect 7182 452898 7266 453134
rect 7502 452898 7534 453134
rect 6914 417454 7534 452898
rect 6914 417218 6946 417454
rect 7182 417218 7266 417454
rect 7502 417218 7534 417454
rect 6914 417134 7534 417218
rect 6914 416898 6946 417134
rect 7182 416898 7266 417134
rect 7502 416898 7534 417134
rect 6914 381454 7534 416898
rect 6914 381218 6946 381454
rect 7182 381218 7266 381454
rect 7502 381218 7534 381454
rect 6914 381134 7534 381218
rect 6914 380898 6946 381134
rect 7182 380898 7266 381134
rect 7502 380898 7534 381134
rect 6914 345454 7534 380898
rect 6914 345218 6946 345454
rect 7182 345218 7266 345454
rect 7502 345218 7534 345454
rect 6914 345134 7534 345218
rect 6914 344898 6946 345134
rect 7182 344898 7266 345134
rect 7502 344898 7534 345134
rect 6914 309454 7534 344898
rect 6914 309218 6946 309454
rect 7182 309218 7266 309454
rect 7502 309218 7534 309454
rect 6914 309134 7534 309218
rect 6914 308898 6946 309134
rect 7182 308898 7266 309134
rect 7502 308898 7534 309134
rect 6914 273454 7534 308898
rect 6914 273218 6946 273454
rect 7182 273218 7266 273454
rect 7502 273218 7534 273454
rect 6914 273134 7534 273218
rect 6914 272898 6946 273134
rect 7182 272898 7266 273134
rect 7502 272898 7534 273134
rect 6914 237454 7534 272898
rect 6914 237218 6946 237454
rect 7182 237218 7266 237454
rect 7502 237218 7534 237454
rect 6914 237134 7534 237218
rect 6914 236898 6946 237134
rect 7182 236898 7266 237134
rect 7502 236898 7534 237134
rect 6914 201454 7534 236898
rect 6914 201218 6946 201454
rect 7182 201218 7266 201454
rect 7502 201218 7534 201454
rect 6914 201134 7534 201218
rect 6914 200898 6946 201134
rect 7182 200898 7266 201134
rect 7502 200898 7534 201134
rect 6914 165454 7534 200898
rect 6914 165218 6946 165454
rect 7182 165218 7266 165454
rect 7502 165218 7534 165454
rect 6914 165134 7534 165218
rect 6914 164898 6946 165134
rect 7182 164898 7266 165134
rect 7502 164898 7534 165134
rect 6914 129454 7534 164898
rect 6914 129218 6946 129454
rect 7182 129218 7266 129454
rect 7502 129218 7534 129454
rect 6914 129134 7534 129218
rect 6914 128898 6946 129134
rect 7182 128898 7266 129134
rect 7502 128898 7534 129134
rect 6914 93454 7534 128898
rect 6914 93218 6946 93454
rect 7182 93218 7266 93454
rect 7502 93218 7534 93454
rect 6914 93134 7534 93218
rect 6914 92898 6946 93134
rect 7182 92898 7266 93134
rect 7502 92898 7534 93134
rect 6914 57454 7534 92898
rect 6914 57218 6946 57454
rect 7182 57218 7266 57454
rect 7502 57218 7534 57454
rect 6914 57134 7534 57218
rect 6914 56898 6946 57134
rect 7182 56898 7266 57134
rect 7502 56898 7534 57134
rect 6914 21454 7534 56898
rect 6914 21218 6946 21454
rect 7182 21218 7266 21454
rect 7502 21218 7534 21454
rect 6914 21134 7534 21218
rect 6914 20898 6946 21134
rect 7182 20898 7266 21134
rect 7502 20898 7534 21134
rect 6914 -1306 7534 20898
rect 6914 -1542 6946 -1306
rect 7182 -1542 7266 -1306
rect 7502 -1542 7534 -1306
rect 6914 -1626 7534 -1542
rect 6914 -1862 6946 -1626
rect 7182 -1862 7266 -1626
rect 7502 -1862 7534 -1626
rect 6914 -1894 7534 -1862
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 10634 707718 11254 707750
rect 10634 707482 10666 707718
rect 10902 707482 10986 707718
rect 11222 707482 11254 707718
rect 10634 707398 11254 707482
rect 10634 707162 10666 707398
rect 10902 707162 10986 707398
rect 11222 707162 11254 707398
rect 10634 673174 11254 707162
rect 10634 672938 10666 673174
rect 10902 672938 10986 673174
rect 11222 672938 11254 673174
rect 10634 672854 11254 672938
rect 10634 672618 10666 672854
rect 10902 672618 10986 672854
rect 11222 672618 11254 672854
rect 10634 637174 11254 672618
rect 10634 636938 10666 637174
rect 10902 636938 10986 637174
rect 11222 636938 11254 637174
rect 10634 636854 11254 636938
rect 10634 636618 10666 636854
rect 10902 636618 10986 636854
rect 11222 636618 11254 636854
rect 10634 601174 11254 636618
rect 10634 600938 10666 601174
rect 10902 600938 10986 601174
rect 11222 600938 11254 601174
rect 10634 600854 11254 600938
rect 10634 600618 10666 600854
rect 10902 600618 10986 600854
rect 11222 600618 11254 600854
rect 10634 565174 11254 600618
rect 10634 564938 10666 565174
rect 10902 564938 10986 565174
rect 11222 564938 11254 565174
rect 10634 564854 11254 564938
rect 10634 564618 10666 564854
rect 10902 564618 10986 564854
rect 11222 564618 11254 564854
rect 10634 529174 11254 564618
rect 10634 528938 10666 529174
rect 10902 528938 10986 529174
rect 11222 528938 11254 529174
rect 10634 528854 11254 528938
rect 10634 528618 10666 528854
rect 10902 528618 10986 528854
rect 11222 528618 11254 528854
rect 10634 493174 11254 528618
rect 10634 492938 10666 493174
rect 10902 492938 10986 493174
rect 11222 492938 11254 493174
rect 10634 492854 11254 492938
rect 10634 492618 10666 492854
rect 10902 492618 10986 492854
rect 11222 492618 11254 492854
rect 10634 457174 11254 492618
rect 10634 456938 10666 457174
rect 10902 456938 10986 457174
rect 11222 456938 11254 457174
rect 10634 456854 11254 456938
rect 10634 456618 10666 456854
rect 10902 456618 10986 456854
rect 11222 456618 11254 456854
rect 10634 421174 11254 456618
rect 10634 420938 10666 421174
rect 10902 420938 10986 421174
rect 11222 420938 11254 421174
rect 10634 420854 11254 420938
rect 10634 420618 10666 420854
rect 10902 420618 10986 420854
rect 11222 420618 11254 420854
rect 10634 385174 11254 420618
rect 10634 384938 10666 385174
rect 10902 384938 10986 385174
rect 11222 384938 11254 385174
rect 10634 384854 11254 384938
rect 10634 384618 10666 384854
rect 10902 384618 10986 384854
rect 11222 384618 11254 384854
rect 10634 349174 11254 384618
rect 10634 348938 10666 349174
rect 10902 348938 10986 349174
rect 11222 348938 11254 349174
rect 10634 348854 11254 348938
rect 10634 348618 10666 348854
rect 10902 348618 10986 348854
rect 11222 348618 11254 348854
rect 10634 313174 11254 348618
rect 10634 312938 10666 313174
rect 10902 312938 10986 313174
rect 11222 312938 11254 313174
rect 10634 312854 11254 312938
rect 10634 312618 10666 312854
rect 10902 312618 10986 312854
rect 11222 312618 11254 312854
rect 10634 277174 11254 312618
rect 10634 276938 10666 277174
rect 10902 276938 10986 277174
rect 11222 276938 11254 277174
rect 10634 276854 11254 276938
rect 10634 276618 10666 276854
rect 10902 276618 10986 276854
rect 11222 276618 11254 276854
rect 10634 241174 11254 276618
rect 10634 240938 10666 241174
rect 10902 240938 10986 241174
rect 11222 240938 11254 241174
rect 10634 240854 11254 240938
rect 10634 240618 10666 240854
rect 10902 240618 10986 240854
rect 11222 240618 11254 240854
rect 10634 205174 11254 240618
rect 10634 204938 10666 205174
rect 10902 204938 10986 205174
rect 11222 204938 11254 205174
rect 10634 204854 11254 204938
rect 10634 204618 10666 204854
rect 10902 204618 10986 204854
rect 11222 204618 11254 204854
rect 10634 169174 11254 204618
rect 10634 168938 10666 169174
rect 10902 168938 10986 169174
rect 11222 168938 11254 169174
rect 10634 168854 11254 168938
rect 10634 168618 10666 168854
rect 10902 168618 10986 168854
rect 11222 168618 11254 168854
rect 10634 133174 11254 168618
rect 10634 132938 10666 133174
rect 10902 132938 10986 133174
rect 11222 132938 11254 133174
rect 10634 132854 11254 132938
rect 10634 132618 10666 132854
rect 10902 132618 10986 132854
rect 11222 132618 11254 132854
rect 10634 97174 11254 132618
rect 10634 96938 10666 97174
rect 10902 96938 10986 97174
rect 11222 96938 11254 97174
rect 10634 96854 11254 96938
rect 10634 96618 10666 96854
rect 10902 96618 10986 96854
rect 11222 96618 11254 96854
rect 10634 61174 11254 96618
rect 10634 60938 10666 61174
rect 10902 60938 10986 61174
rect 11222 60938 11254 61174
rect 10634 60854 11254 60938
rect 10634 60618 10666 60854
rect 10902 60618 10986 60854
rect 11222 60618 11254 60854
rect 10634 25174 11254 60618
rect 10634 24938 10666 25174
rect 10902 24938 10986 25174
rect 11222 24938 11254 25174
rect 10634 24854 11254 24938
rect 10634 24618 10666 24854
rect 10902 24618 10986 24854
rect 11222 24618 11254 24854
rect 10634 -3226 11254 24618
rect 12034 704838 12654 705830
rect 12034 704602 12066 704838
rect 12302 704602 12386 704838
rect 12622 704602 12654 704838
rect 12034 704518 12654 704602
rect 12034 704282 12066 704518
rect 12302 704282 12386 704518
rect 12622 704282 12654 704518
rect 12034 687454 12654 704282
rect 12034 687218 12066 687454
rect 12302 687218 12386 687454
rect 12622 687218 12654 687454
rect 12034 687134 12654 687218
rect 12034 686898 12066 687134
rect 12302 686898 12386 687134
rect 12622 686898 12654 687134
rect 12034 651454 12654 686898
rect 12034 651218 12066 651454
rect 12302 651218 12386 651454
rect 12622 651218 12654 651454
rect 12034 651134 12654 651218
rect 12034 650898 12066 651134
rect 12302 650898 12386 651134
rect 12622 650898 12654 651134
rect 12034 615454 12654 650898
rect 12034 615218 12066 615454
rect 12302 615218 12386 615454
rect 12622 615218 12654 615454
rect 12034 615134 12654 615218
rect 12034 614898 12066 615134
rect 12302 614898 12386 615134
rect 12622 614898 12654 615134
rect 12034 579454 12654 614898
rect 12034 579218 12066 579454
rect 12302 579218 12386 579454
rect 12622 579218 12654 579454
rect 12034 579134 12654 579218
rect 12034 578898 12066 579134
rect 12302 578898 12386 579134
rect 12622 578898 12654 579134
rect 12034 543454 12654 578898
rect 12034 543218 12066 543454
rect 12302 543218 12386 543454
rect 12622 543218 12654 543454
rect 12034 543134 12654 543218
rect 12034 542898 12066 543134
rect 12302 542898 12386 543134
rect 12622 542898 12654 543134
rect 12034 507454 12654 542898
rect 12034 507218 12066 507454
rect 12302 507218 12386 507454
rect 12622 507218 12654 507454
rect 12034 507134 12654 507218
rect 12034 506898 12066 507134
rect 12302 506898 12386 507134
rect 12622 506898 12654 507134
rect 12034 471454 12654 506898
rect 12034 471218 12066 471454
rect 12302 471218 12386 471454
rect 12622 471218 12654 471454
rect 12034 471134 12654 471218
rect 12034 470898 12066 471134
rect 12302 470898 12386 471134
rect 12622 470898 12654 471134
rect 12034 435454 12654 470898
rect 12034 435218 12066 435454
rect 12302 435218 12386 435454
rect 12622 435218 12654 435454
rect 12034 435134 12654 435218
rect 12034 434898 12066 435134
rect 12302 434898 12386 435134
rect 12622 434898 12654 435134
rect 12034 399454 12654 434898
rect 12034 399218 12066 399454
rect 12302 399218 12386 399454
rect 12622 399218 12654 399454
rect 12034 399134 12654 399218
rect 12034 398898 12066 399134
rect 12302 398898 12386 399134
rect 12622 398898 12654 399134
rect 12034 363454 12654 398898
rect 12034 363218 12066 363454
rect 12302 363218 12386 363454
rect 12622 363218 12654 363454
rect 12034 363134 12654 363218
rect 12034 362898 12066 363134
rect 12302 362898 12386 363134
rect 12622 362898 12654 363134
rect 12034 327454 12654 362898
rect 12034 327218 12066 327454
rect 12302 327218 12386 327454
rect 12622 327218 12654 327454
rect 12034 327134 12654 327218
rect 12034 326898 12066 327134
rect 12302 326898 12386 327134
rect 12622 326898 12654 327134
rect 12034 291454 12654 326898
rect 12034 291218 12066 291454
rect 12302 291218 12386 291454
rect 12622 291218 12654 291454
rect 12034 291134 12654 291218
rect 12034 290898 12066 291134
rect 12302 290898 12386 291134
rect 12622 290898 12654 291134
rect 12034 255454 12654 290898
rect 12034 255218 12066 255454
rect 12302 255218 12386 255454
rect 12622 255218 12654 255454
rect 12034 255134 12654 255218
rect 12034 254898 12066 255134
rect 12302 254898 12386 255134
rect 12622 254898 12654 255134
rect 12034 219454 12654 254898
rect 12034 219218 12066 219454
rect 12302 219218 12386 219454
rect 12622 219218 12654 219454
rect 12034 219134 12654 219218
rect 12034 218898 12066 219134
rect 12302 218898 12386 219134
rect 12622 218898 12654 219134
rect 12034 183454 12654 218898
rect 12034 183218 12066 183454
rect 12302 183218 12386 183454
rect 12622 183218 12654 183454
rect 12034 183134 12654 183218
rect 12034 182898 12066 183134
rect 12302 182898 12386 183134
rect 12622 182898 12654 183134
rect 12034 147454 12654 182898
rect 12034 147218 12066 147454
rect 12302 147218 12386 147454
rect 12622 147218 12654 147454
rect 12034 147134 12654 147218
rect 12034 146898 12066 147134
rect 12302 146898 12386 147134
rect 12622 146898 12654 147134
rect 12034 111454 12654 146898
rect 12034 111218 12066 111454
rect 12302 111218 12386 111454
rect 12622 111218 12654 111454
rect 12034 111134 12654 111218
rect 12034 110898 12066 111134
rect 12302 110898 12386 111134
rect 12622 110898 12654 111134
rect 12034 75454 12654 110898
rect 12034 75218 12066 75454
rect 12302 75218 12386 75454
rect 12622 75218 12654 75454
rect 12034 75134 12654 75218
rect 12034 74898 12066 75134
rect 12302 74898 12386 75134
rect 12622 74898 12654 75134
rect 12034 39454 12654 74898
rect 12034 39218 12066 39454
rect 12302 39218 12386 39454
rect 12622 39218 12654 39454
rect 12034 39134 12654 39218
rect 12034 38898 12066 39134
rect 12302 38898 12386 39134
rect 12622 38898 12654 39134
rect 12034 3454 12654 38898
rect 12034 3218 12066 3454
rect 12302 3218 12386 3454
rect 12622 3218 12654 3454
rect 12034 3134 12654 3218
rect 12034 2898 12066 3134
rect 12302 2898 12386 3134
rect 12622 2898 12654 3134
rect 12034 -346 12654 2898
rect 12034 -582 12066 -346
rect 12302 -582 12386 -346
rect 12622 -582 12654 -346
rect 12034 -666 12654 -582
rect 12034 -902 12066 -666
rect 12302 -902 12386 -666
rect 12622 -902 12654 -666
rect 12034 -1894 12654 -902
rect 12954 698614 13574 710042
rect 18074 711558 18694 711590
rect 18074 711322 18106 711558
rect 18342 711322 18426 711558
rect 18662 711322 18694 711558
rect 18074 711238 18694 711322
rect 18074 711002 18106 711238
rect 18342 711002 18426 711238
rect 18662 711002 18694 711238
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 10634 -3462 10666 -3226
rect 10902 -3462 10986 -3226
rect 11222 -3462 11254 -3226
rect 10634 -3546 11254 -3462
rect 10634 -3782 10666 -3546
rect 10902 -3782 10986 -3546
rect 11222 -3782 11254 -3546
rect 10634 -3814 11254 -3782
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 14354 709638 14974 709670
rect 14354 709402 14386 709638
rect 14622 709402 14706 709638
rect 14942 709402 14974 709638
rect 14354 709318 14974 709402
rect 14354 709082 14386 709318
rect 14622 709082 14706 709318
rect 14942 709082 14974 709318
rect 14354 676894 14974 709082
rect 14354 676658 14386 676894
rect 14622 676658 14706 676894
rect 14942 676658 14974 676894
rect 14354 676574 14974 676658
rect 14354 676338 14386 676574
rect 14622 676338 14706 676574
rect 14942 676338 14974 676574
rect 14354 640894 14974 676338
rect 14354 640658 14386 640894
rect 14622 640658 14706 640894
rect 14942 640658 14974 640894
rect 14354 640574 14974 640658
rect 14354 640338 14386 640574
rect 14622 640338 14706 640574
rect 14942 640338 14974 640574
rect 14354 604894 14974 640338
rect 14354 604658 14386 604894
rect 14622 604658 14706 604894
rect 14942 604658 14974 604894
rect 14354 604574 14974 604658
rect 14354 604338 14386 604574
rect 14622 604338 14706 604574
rect 14942 604338 14974 604574
rect 14354 568894 14974 604338
rect 14354 568658 14386 568894
rect 14622 568658 14706 568894
rect 14942 568658 14974 568894
rect 14354 568574 14974 568658
rect 14354 568338 14386 568574
rect 14622 568338 14706 568574
rect 14942 568338 14974 568574
rect 14354 532894 14974 568338
rect 14354 532658 14386 532894
rect 14622 532658 14706 532894
rect 14942 532658 14974 532894
rect 14354 532574 14974 532658
rect 14354 532338 14386 532574
rect 14622 532338 14706 532574
rect 14942 532338 14974 532574
rect 14354 496894 14974 532338
rect 14354 496658 14386 496894
rect 14622 496658 14706 496894
rect 14942 496658 14974 496894
rect 14354 496574 14974 496658
rect 14354 496338 14386 496574
rect 14622 496338 14706 496574
rect 14942 496338 14974 496574
rect 14354 460894 14974 496338
rect 14354 460658 14386 460894
rect 14622 460658 14706 460894
rect 14942 460658 14974 460894
rect 14354 460574 14974 460658
rect 14354 460338 14386 460574
rect 14622 460338 14706 460574
rect 14942 460338 14974 460574
rect 14354 424894 14974 460338
rect 14354 424658 14386 424894
rect 14622 424658 14706 424894
rect 14942 424658 14974 424894
rect 14354 424574 14974 424658
rect 14354 424338 14386 424574
rect 14622 424338 14706 424574
rect 14942 424338 14974 424574
rect 14354 388894 14974 424338
rect 14354 388658 14386 388894
rect 14622 388658 14706 388894
rect 14942 388658 14974 388894
rect 14354 388574 14974 388658
rect 14354 388338 14386 388574
rect 14622 388338 14706 388574
rect 14942 388338 14974 388574
rect 14354 352894 14974 388338
rect 14354 352658 14386 352894
rect 14622 352658 14706 352894
rect 14942 352658 14974 352894
rect 14354 352574 14974 352658
rect 14354 352338 14386 352574
rect 14622 352338 14706 352574
rect 14942 352338 14974 352574
rect 14354 316894 14974 352338
rect 14354 316658 14386 316894
rect 14622 316658 14706 316894
rect 14942 316658 14974 316894
rect 14354 316574 14974 316658
rect 14354 316338 14386 316574
rect 14622 316338 14706 316574
rect 14942 316338 14974 316574
rect 14354 280894 14974 316338
rect 14354 280658 14386 280894
rect 14622 280658 14706 280894
rect 14942 280658 14974 280894
rect 14354 280574 14974 280658
rect 14354 280338 14386 280574
rect 14622 280338 14706 280574
rect 14942 280338 14974 280574
rect 14354 244894 14974 280338
rect 14354 244658 14386 244894
rect 14622 244658 14706 244894
rect 14942 244658 14974 244894
rect 14354 244574 14974 244658
rect 14354 244338 14386 244574
rect 14622 244338 14706 244574
rect 14942 244338 14974 244574
rect 14354 208894 14974 244338
rect 14354 208658 14386 208894
rect 14622 208658 14706 208894
rect 14942 208658 14974 208894
rect 14354 208574 14974 208658
rect 14354 208338 14386 208574
rect 14622 208338 14706 208574
rect 14942 208338 14974 208574
rect 14354 172894 14974 208338
rect 14354 172658 14386 172894
rect 14622 172658 14706 172894
rect 14942 172658 14974 172894
rect 14354 172574 14974 172658
rect 14354 172338 14386 172574
rect 14622 172338 14706 172574
rect 14942 172338 14974 172574
rect 14354 136894 14974 172338
rect 14354 136658 14386 136894
rect 14622 136658 14706 136894
rect 14942 136658 14974 136894
rect 14354 136574 14974 136658
rect 14354 136338 14386 136574
rect 14622 136338 14706 136574
rect 14942 136338 14974 136574
rect 14354 100894 14974 136338
rect 14354 100658 14386 100894
rect 14622 100658 14706 100894
rect 14942 100658 14974 100894
rect 14354 100574 14974 100658
rect 14354 100338 14386 100574
rect 14622 100338 14706 100574
rect 14942 100338 14974 100574
rect 14354 64894 14974 100338
rect 14354 64658 14386 64894
rect 14622 64658 14706 64894
rect 14942 64658 14974 64894
rect 14354 64574 14974 64658
rect 14354 64338 14386 64574
rect 14622 64338 14706 64574
rect 14942 64338 14974 64574
rect 14354 28894 14974 64338
rect 14354 28658 14386 28894
rect 14622 28658 14706 28894
rect 14942 28658 14974 28894
rect 14354 28574 14974 28658
rect 14354 28338 14386 28574
rect 14622 28338 14706 28574
rect 14942 28338 14974 28574
rect 14354 -5146 14974 28338
rect 15754 706758 16374 707750
rect 15754 706522 15786 706758
rect 16022 706522 16106 706758
rect 16342 706522 16374 706758
rect 15754 706438 16374 706522
rect 15754 706202 15786 706438
rect 16022 706202 16106 706438
rect 16342 706202 16374 706438
rect 15754 691174 16374 706202
rect 15754 690938 15786 691174
rect 16022 690938 16106 691174
rect 16342 690938 16374 691174
rect 15754 690854 16374 690938
rect 15754 690618 15786 690854
rect 16022 690618 16106 690854
rect 16342 690618 16374 690854
rect 15754 655174 16374 690618
rect 17154 705798 17774 705830
rect 17154 705562 17186 705798
rect 17422 705562 17506 705798
rect 17742 705562 17774 705798
rect 17154 705478 17774 705562
rect 17154 705242 17186 705478
rect 17422 705242 17506 705478
rect 17742 705242 17774 705478
rect 17154 669454 17774 705242
rect 17154 669218 17186 669454
rect 17422 669218 17506 669454
rect 17742 669218 17774 669454
rect 17154 669134 17774 669218
rect 17154 668898 17186 669134
rect 17422 668898 17506 669134
rect 17742 668898 17774 669134
rect 17154 657000 17774 668898
rect 18074 680614 18694 711002
rect 23194 710598 23814 711590
rect 23194 710362 23226 710598
rect 23462 710362 23546 710598
rect 23782 710362 23814 710598
rect 23194 710278 23814 710362
rect 23194 710042 23226 710278
rect 23462 710042 23546 710278
rect 23782 710042 23814 710278
rect 18074 680378 18106 680614
rect 18342 680378 18426 680614
rect 18662 680378 18694 680614
rect 18074 680294 18694 680378
rect 18074 680058 18106 680294
rect 18342 680058 18426 680294
rect 18662 680058 18694 680294
rect 18074 657000 18694 680058
rect 19474 708678 20094 709670
rect 19474 708442 19506 708678
rect 19742 708442 19826 708678
rect 20062 708442 20094 708678
rect 19474 708358 20094 708442
rect 19474 708122 19506 708358
rect 19742 708122 19826 708358
rect 20062 708122 20094 708358
rect 19474 694894 20094 708122
rect 19474 694658 19506 694894
rect 19742 694658 19826 694894
rect 20062 694658 20094 694894
rect 19474 694574 20094 694658
rect 19474 694338 19506 694574
rect 19742 694338 19826 694574
rect 20062 694338 20094 694574
rect 19474 658894 20094 694338
rect 19474 658658 19506 658894
rect 19742 658658 19826 658894
rect 20062 658658 20094 658894
rect 19474 658574 20094 658658
rect 19474 658338 19506 658574
rect 19742 658338 19826 658574
rect 20062 658338 20094 658574
rect 19474 657000 20094 658338
rect 20874 707718 21494 707750
rect 20874 707482 20906 707718
rect 21142 707482 21226 707718
rect 21462 707482 21494 707718
rect 20874 707398 21494 707482
rect 20874 707162 20906 707398
rect 21142 707162 21226 707398
rect 21462 707162 21494 707398
rect 20874 673174 21494 707162
rect 20874 672938 20906 673174
rect 21142 672938 21226 673174
rect 21462 672938 21494 673174
rect 20874 672854 21494 672938
rect 20874 672618 20906 672854
rect 21142 672618 21226 672854
rect 21462 672618 21494 672854
rect 20874 657000 21494 672618
rect 22274 704838 22894 705830
rect 22274 704602 22306 704838
rect 22542 704602 22626 704838
rect 22862 704602 22894 704838
rect 22274 704518 22894 704602
rect 22274 704282 22306 704518
rect 22542 704282 22626 704518
rect 22862 704282 22894 704518
rect 22274 687454 22894 704282
rect 22274 687218 22306 687454
rect 22542 687218 22626 687454
rect 22862 687218 22894 687454
rect 22274 687134 22894 687218
rect 22274 686898 22306 687134
rect 22542 686898 22626 687134
rect 22862 686898 22894 687134
rect 22274 657000 22894 686898
rect 23194 698614 23814 710042
rect 28314 711558 28934 711590
rect 28314 711322 28346 711558
rect 28582 711322 28666 711558
rect 28902 711322 28934 711558
rect 28314 711238 28934 711322
rect 28314 711002 28346 711238
rect 28582 711002 28666 711238
rect 28902 711002 28934 711238
rect 23194 698378 23226 698614
rect 23462 698378 23546 698614
rect 23782 698378 23814 698614
rect 23194 698294 23814 698378
rect 23194 698058 23226 698294
rect 23462 698058 23546 698294
rect 23782 698058 23814 698294
rect 23194 662614 23814 698058
rect 23194 662378 23226 662614
rect 23462 662378 23546 662614
rect 23782 662378 23814 662614
rect 23194 662294 23814 662378
rect 23194 662058 23226 662294
rect 23462 662058 23546 662294
rect 23782 662058 23814 662294
rect 23194 657000 23814 662058
rect 24594 709638 25214 709670
rect 24594 709402 24626 709638
rect 24862 709402 24946 709638
rect 25182 709402 25214 709638
rect 24594 709318 25214 709402
rect 24594 709082 24626 709318
rect 24862 709082 24946 709318
rect 25182 709082 25214 709318
rect 24594 676894 25214 709082
rect 24594 676658 24626 676894
rect 24862 676658 24946 676894
rect 25182 676658 25214 676894
rect 24594 676574 25214 676658
rect 24594 676338 24626 676574
rect 24862 676338 24946 676574
rect 25182 676338 25214 676574
rect 24594 657000 25214 676338
rect 25994 706758 26614 707750
rect 25994 706522 26026 706758
rect 26262 706522 26346 706758
rect 26582 706522 26614 706758
rect 25994 706438 26614 706522
rect 25994 706202 26026 706438
rect 26262 706202 26346 706438
rect 26582 706202 26614 706438
rect 25994 691174 26614 706202
rect 25994 690938 26026 691174
rect 26262 690938 26346 691174
rect 26582 690938 26614 691174
rect 25994 690854 26614 690938
rect 25994 690618 26026 690854
rect 26262 690618 26346 690854
rect 26582 690618 26614 690854
rect 25994 657000 26614 690618
rect 27394 705798 28014 705830
rect 27394 705562 27426 705798
rect 27662 705562 27746 705798
rect 27982 705562 28014 705798
rect 27394 705478 28014 705562
rect 27394 705242 27426 705478
rect 27662 705242 27746 705478
rect 27982 705242 28014 705478
rect 27394 669454 28014 705242
rect 27394 669218 27426 669454
rect 27662 669218 27746 669454
rect 27982 669218 28014 669454
rect 27394 669134 28014 669218
rect 27394 668898 27426 669134
rect 27662 668898 27746 669134
rect 27982 668898 28014 669134
rect 27394 657000 28014 668898
rect 28314 680614 28934 711002
rect 33434 710598 34054 711590
rect 33434 710362 33466 710598
rect 33702 710362 33786 710598
rect 34022 710362 34054 710598
rect 33434 710278 34054 710362
rect 33434 710042 33466 710278
rect 33702 710042 33786 710278
rect 34022 710042 34054 710278
rect 28314 680378 28346 680614
rect 28582 680378 28666 680614
rect 28902 680378 28934 680614
rect 28314 680294 28934 680378
rect 28314 680058 28346 680294
rect 28582 680058 28666 680294
rect 28902 680058 28934 680294
rect 28314 657000 28934 680058
rect 29714 708678 30334 709670
rect 29714 708442 29746 708678
rect 29982 708442 30066 708678
rect 30302 708442 30334 708678
rect 29714 708358 30334 708442
rect 29714 708122 29746 708358
rect 29982 708122 30066 708358
rect 30302 708122 30334 708358
rect 29714 694894 30334 708122
rect 29714 694658 29746 694894
rect 29982 694658 30066 694894
rect 30302 694658 30334 694894
rect 29714 694574 30334 694658
rect 29714 694338 29746 694574
rect 29982 694338 30066 694574
rect 30302 694338 30334 694574
rect 29714 658894 30334 694338
rect 29714 658658 29746 658894
rect 29982 658658 30066 658894
rect 30302 658658 30334 658894
rect 29714 658574 30334 658658
rect 29714 658338 29746 658574
rect 29982 658338 30066 658574
rect 30302 658338 30334 658574
rect 29714 657000 30334 658338
rect 31114 707718 31734 707750
rect 31114 707482 31146 707718
rect 31382 707482 31466 707718
rect 31702 707482 31734 707718
rect 31114 707398 31734 707482
rect 31114 707162 31146 707398
rect 31382 707162 31466 707398
rect 31702 707162 31734 707398
rect 31114 673174 31734 707162
rect 31114 672938 31146 673174
rect 31382 672938 31466 673174
rect 31702 672938 31734 673174
rect 31114 672854 31734 672938
rect 31114 672618 31146 672854
rect 31382 672618 31466 672854
rect 31702 672618 31734 672854
rect 31114 657000 31734 672618
rect 32514 704838 33134 705830
rect 32514 704602 32546 704838
rect 32782 704602 32866 704838
rect 33102 704602 33134 704838
rect 32514 704518 33134 704602
rect 32514 704282 32546 704518
rect 32782 704282 32866 704518
rect 33102 704282 33134 704518
rect 32514 687454 33134 704282
rect 32514 687218 32546 687454
rect 32782 687218 32866 687454
rect 33102 687218 33134 687454
rect 32514 687134 33134 687218
rect 32514 686898 32546 687134
rect 32782 686898 32866 687134
rect 33102 686898 33134 687134
rect 32514 657000 33134 686898
rect 33434 698614 34054 710042
rect 38554 711558 39174 711590
rect 38554 711322 38586 711558
rect 38822 711322 38906 711558
rect 39142 711322 39174 711558
rect 38554 711238 39174 711322
rect 38554 711002 38586 711238
rect 38822 711002 38906 711238
rect 39142 711002 39174 711238
rect 33434 698378 33466 698614
rect 33702 698378 33786 698614
rect 34022 698378 34054 698614
rect 33434 698294 34054 698378
rect 33434 698058 33466 698294
rect 33702 698058 33786 698294
rect 34022 698058 34054 698294
rect 33434 662614 34054 698058
rect 33434 662378 33466 662614
rect 33702 662378 33786 662614
rect 34022 662378 34054 662614
rect 33434 662294 34054 662378
rect 33434 662058 33466 662294
rect 33702 662058 33786 662294
rect 34022 662058 34054 662294
rect 33434 657000 34054 662058
rect 34834 709638 35454 709670
rect 34834 709402 34866 709638
rect 35102 709402 35186 709638
rect 35422 709402 35454 709638
rect 34834 709318 35454 709402
rect 34834 709082 34866 709318
rect 35102 709082 35186 709318
rect 35422 709082 35454 709318
rect 34834 676894 35454 709082
rect 34834 676658 34866 676894
rect 35102 676658 35186 676894
rect 35422 676658 35454 676894
rect 34834 676574 35454 676658
rect 34834 676338 34866 676574
rect 35102 676338 35186 676574
rect 35422 676338 35454 676574
rect 34834 657000 35454 676338
rect 36234 706758 36854 707750
rect 36234 706522 36266 706758
rect 36502 706522 36586 706758
rect 36822 706522 36854 706758
rect 36234 706438 36854 706522
rect 36234 706202 36266 706438
rect 36502 706202 36586 706438
rect 36822 706202 36854 706438
rect 36234 691174 36854 706202
rect 36234 690938 36266 691174
rect 36502 690938 36586 691174
rect 36822 690938 36854 691174
rect 36234 690854 36854 690938
rect 36234 690618 36266 690854
rect 36502 690618 36586 690854
rect 36822 690618 36854 690854
rect 36234 657000 36854 690618
rect 37634 705798 38254 705830
rect 37634 705562 37666 705798
rect 37902 705562 37986 705798
rect 38222 705562 38254 705798
rect 37634 705478 38254 705562
rect 37634 705242 37666 705478
rect 37902 705242 37986 705478
rect 38222 705242 38254 705478
rect 37634 669454 38254 705242
rect 37634 669218 37666 669454
rect 37902 669218 37986 669454
rect 38222 669218 38254 669454
rect 37634 669134 38254 669218
rect 37634 668898 37666 669134
rect 37902 668898 37986 669134
rect 38222 668898 38254 669134
rect 37634 657000 38254 668898
rect 38554 680614 39174 711002
rect 43674 710598 44294 711590
rect 43674 710362 43706 710598
rect 43942 710362 44026 710598
rect 44262 710362 44294 710598
rect 43674 710278 44294 710362
rect 43674 710042 43706 710278
rect 43942 710042 44026 710278
rect 44262 710042 44294 710278
rect 38554 680378 38586 680614
rect 38822 680378 38906 680614
rect 39142 680378 39174 680614
rect 38554 680294 39174 680378
rect 38554 680058 38586 680294
rect 38822 680058 38906 680294
rect 39142 680058 39174 680294
rect 38554 657000 39174 680058
rect 39954 708678 40574 709670
rect 39954 708442 39986 708678
rect 40222 708442 40306 708678
rect 40542 708442 40574 708678
rect 39954 708358 40574 708442
rect 39954 708122 39986 708358
rect 40222 708122 40306 708358
rect 40542 708122 40574 708358
rect 39954 694894 40574 708122
rect 39954 694658 39986 694894
rect 40222 694658 40306 694894
rect 40542 694658 40574 694894
rect 39954 694574 40574 694658
rect 39954 694338 39986 694574
rect 40222 694338 40306 694574
rect 40542 694338 40574 694574
rect 39954 658894 40574 694338
rect 39954 658658 39986 658894
rect 40222 658658 40306 658894
rect 40542 658658 40574 658894
rect 39954 658574 40574 658658
rect 39954 658338 39986 658574
rect 40222 658338 40306 658574
rect 40542 658338 40574 658574
rect 39954 657000 40574 658338
rect 41354 707718 41974 707750
rect 41354 707482 41386 707718
rect 41622 707482 41706 707718
rect 41942 707482 41974 707718
rect 41354 707398 41974 707482
rect 41354 707162 41386 707398
rect 41622 707162 41706 707398
rect 41942 707162 41974 707398
rect 41354 673174 41974 707162
rect 41354 672938 41386 673174
rect 41622 672938 41706 673174
rect 41942 672938 41974 673174
rect 41354 672854 41974 672938
rect 41354 672618 41386 672854
rect 41622 672618 41706 672854
rect 41942 672618 41974 672854
rect 41354 657000 41974 672618
rect 42754 704838 43374 705830
rect 42754 704602 42786 704838
rect 43022 704602 43106 704838
rect 43342 704602 43374 704838
rect 42754 704518 43374 704602
rect 42754 704282 42786 704518
rect 43022 704282 43106 704518
rect 43342 704282 43374 704518
rect 42754 687454 43374 704282
rect 42754 687218 42786 687454
rect 43022 687218 43106 687454
rect 43342 687218 43374 687454
rect 42754 687134 43374 687218
rect 42754 686898 42786 687134
rect 43022 686898 43106 687134
rect 43342 686898 43374 687134
rect 42754 657000 43374 686898
rect 43674 698614 44294 710042
rect 48794 711558 49414 711590
rect 48794 711322 48826 711558
rect 49062 711322 49146 711558
rect 49382 711322 49414 711558
rect 48794 711238 49414 711322
rect 48794 711002 48826 711238
rect 49062 711002 49146 711238
rect 49382 711002 49414 711238
rect 43674 698378 43706 698614
rect 43942 698378 44026 698614
rect 44262 698378 44294 698614
rect 43674 698294 44294 698378
rect 43674 698058 43706 698294
rect 43942 698058 44026 698294
rect 44262 698058 44294 698294
rect 43674 662614 44294 698058
rect 43674 662378 43706 662614
rect 43942 662378 44026 662614
rect 44262 662378 44294 662614
rect 43674 662294 44294 662378
rect 43674 662058 43706 662294
rect 43942 662058 44026 662294
rect 44262 662058 44294 662294
rect 43674 657000 44294 662058
rect 45074 709638 45694 709670
rect 45074 709402 45106 709638
rect 45342 709402 45426 709638
rect 45662 709402 45694 709638
rect 45074 709318 45694 709402
rect 45074 709082 45106 709318
rect 45342 709082 45426 709318
rect 45662 709082 45694 709318
rect 45074 676894 45694 709082
rect 45074 676658 45106 676894
rect 45342 676658 45426 676894
rect 45662 676658 45694 676894
rect 45074 676574 45694 676658
rect 45074 676338 45106 676574
rect 45342 676338 45426 676574
rect 45662 676338 45694 676574
rect 45074 657000 45694 676338
rect 46474 706758 47094 707750
rect 46474 706522 46506 706758
rect 46742 706522 46826 706758
rect 47062 706522 47094 706758
rect 46474 706438 47094 706522
rect 46474 706202 46506 706438
rect 46742 706202 46826 706438
rect 47062 706202 47094 706438
rect 46474 691174 47094 706202
rect 46474 690938 46506 691174
rect 46742 690938 46826 691174
rect 47062 690938 47094 691174
rect 46474 690854 47094 690938
rect 46474 690618 46506 690854
rect 46742 690618 46826 690854
rect 47062 690618 47094 690854
rect 46474 657000 47094 690618
rect 47874 705798 48494 705830
rect 47874 705562 47906 705798
rect 48142 705562 48226 705798
rect 48462 705562 48494 705798
rect 47874 705478 48494 705562
rect 47874 705242 47906 705478
rect 48142 705242 48226 705478
rect 48462 705242 48494 705478
rect 47874 669454 48494 705242
rect 47874 669218 47906 669454
rect 48142 669218 48226 669454
rect 48462 669218 48494 669454
rect 47874 669134 48494 669218
rect 47874 668898 47906 669134
rect 48142 668898 48226 669134
rect 48462 668898 48494 669134
rect 47874 657000 48494 668898
rect 48794 680614 49414 711002
rect 53914 710598 54534 711590
rect 53914 710362 53946 710598
rect 54182 710362 54266 710598
rect 54502 710362 54534 710598
rect 53914 710278 54534 710362
rect 53914 710042 53946 710278
rect 54182 710042 54266 710278
rect 54502 710042 54534 710278
rect 48794 680378 48826 680614
rect 49062 680378 49146 680614
rect 49382 680378 49414 680614
rect 48794 680294 49414 680378
rect 48794 680058 48826 680294
rect 49062 680058 49146 680294
rect 49382 680058 49414 680294
rect 48794 657000 49414 680058
rect 50194 708678 50814 709670
rect 50194 708442 50226 708678
rect 50462 708442 50546 708678
rect 50782 708442 50814 708678
rect 50194 708358 50814 708442
rect 50194 708122 50226 708358
rect 50462 708122 50546 708358
rect 50782 708122 50814 708358
rect 50194 694894 50814 708122
rect 50194 694658 50226 694894
rect 50462 694658 50546 694894
rect 50782 694658 50814 694894
rect 50194 694574 50814 694658
rect 50194 694338 50226 694574
rect 50462 694338 50546 694574
rect 50782 694338 50814 694574
rect 50194 658894 50814 694338
rect 50194 658658 50226 658894
rect 50462 658658 50546 658894
rect 50782 658658 50814 658894
rect 50194 658574 50814 658658
rect 50194 658338 50226 658574
rect 50462 658338 50546 658574
rect 50782 658338 50814 658574
rect 50194 657000 50814 658338
rect 51594 707718 52214 707750
rect 51594 707482 51626 707718
rect 51862 707482 51946 707718
rect 52182 707482 52214 707718
rect 51594 707398 52214 707482
rect 51594 707162 51626 707398
rect 51862 707162 51946 707398
rect 52182 707162 52214 707398
rect 51594 673174 52214 707162
rect 51594 672938 51626 673174
rect 51862 672938 51946 673174
rect 52182 672938 52214 673174
rect 51594 672854 52214 672938
rect 51594 672618 51626 672854
rect 51862 672618 51946 672854
rect 52182 672618 52214 672854
rect 51594 657000 52214 672618
rect 52994 704838 53614 705830
rect 52994 704602 53026 704838
rect 53262 704602 53346 704838
rect 53582 704602 53614 704838
rect 52994 704518 53614 704602
rect 52994 704282 53026 704518
rect 53262 704282 53346 704518
rect 53582 704282 53614 704518
rect 52994 687454 53614 704282
rect 52994 687218 53026 687454
rect 53262 687218 53346 687454
rect 53582 687218 53614 687454
rect 52994 687134 53614 687218
rect 52994 686898 53026 687134
rect 53262 686898 53346 687134
rect 53582 686898 53614 687134
rect 52994 657000 53614 686898
rect 53914 698614 54534 710042
rect 59034 711558 59654 711590
rect 59034 711322 59066 711558
rect 59302 711322 59386 711558
rect 59622 711322 59654 711558
rect 59034 711238 59654 711322
rect 59034 711002 59066 711238
rect 59302 711002 59386 711238
rect 59622 711002 59654 711238
rect 53914 698378 53946 698614
rect 54182 698378 54266 698614
rect 54502 698378 54534 698614
rect 53914 698294 54534 698378
rect 53914 698058 53946 698294
rect 54182 698058 54266 698294
rect 54502 698058 54534 698294
rect 53914 662614 54534 698058
rect 53914 662378 53946 662614
rect 54182 662378 54266 662614
rect 54502 662378 54534 662614
rect 53914 662294 54534 662378
rect 53914 662058 53946 662294
rect 54182 662058 54266 662294
rect 54502 662058 54534 662294
rect 53914 657000 54534 662058
rect 55314 709638 55934 709670
rect 55314 709402 55346 709638
rect 55582 709402 55666 709638
rect 55902 709402 55934 709638
rect 55314 709318 55934 709402
rect 55314 709082 55346 709318
rect 55582 709082 55666 709318
rect 55902 709082 55934 709318
rect 55314 676894 55934 709082
rect 55314 676658 55346 676894
rect 55582 676658 55666 676894
rect 55902 676658 55934 676894
rect 55314 676574 55934 676658
rect 55314 676338 55346 676574
rect 55582 676338 55666 676574
rect 55902 676338 55934 676574
rect 55314 657000 55934 676338
rect 56714 706758 57334 707750
rect 56714 706522 56746 706758
rect 56982 706522 57066 706758
rect 57302 706522 57334 706758
rect 56714 706438 57334 706522
rect 56714 706202 56746 706438
rect 56982 706202 57066 706438
rect 57302 706202 57334 706438
rect 56714 691174 57334 706202
rect 56714 690938 56746 691174
rect 56982 690938 57066 691174
rect 57302 690938 57334 691174
rect 56714 690854 57334 690938
rect 56714 690618 56746 690854
rect 56982 690618 57066 690854
rect 57302 690618 57334 690854
rect 56714 657000 57334 690618
rect 58114 705798 58734 705830
rect 58114 705562 58146 705798
rect 58382 705562 58466 705798
rect 58702 705562 58734 705798
rect 58114 705478 58734 705562
rect 58114 705242 58146 705478
rect 58382 705242 58466 705478
rect 58702 705242 58734 705478
rect 58114 669454 58734 705242
rect 58114 669218 58146 669454
rect 58382 669218 58466 669454
rect 58702 669218 58734 669454
rect 58114 669134 58734 669218
rect 58114 668898 58146 669134
rect 58382 668898 58466 669134
rect 58702 668898 58734 669134
rect 58114 657000 58734 668898
rect 59034 680614 59654 711002
rect 64154 710598 64774 711590
rect 64154 710362 64186 710598
rect 64422 710362 64506 710598
rect 64742 710362 64774 710598
rect 64154 710278 64774 710362
rect 64154 710042 64186 710278
rect 64422 710042 64506 710278
rect 64742 710042 64774 710278
rect 59034 680378 59066 680614
rect 59302 680378 59386 680614
rect 59622 680378 59654 680614
rect 59034 680294 59654 680378
rect 59034 680058 59066 680294
rect 59302 680058 59386 680294
rect 59622 680058 59654 680294
rect 59034 657000 59654 680058
rect 60434 708678 61054 709670
rect 60434 708442 60466 708678
rect 60702 708442 60786 708678
rect 61022 708442 61054 708678
rect 60434 708358 61054 708442
rect 60434 708122 60466 708358
rect 60702 708122 60786 708358
rect 61022 708122 61054 708358
rect 60434 694894 61054 708122
rect 60434 694658 60466 694894
rect 60702 694658 60786 694894
rect 61022 694658 61054 694894
rect 60434 694574 61054 694658
rect 60434 694338 60466 694574
rect 60702 694338 60786 694574
rect 61022 694338 61054 694574
rect 60434 658894 61054 694338
rect 60434 658658 60466 658894
rect 60702 658658 60786 658894
rect 61022 658658 61054 658894
rect 60434 658574 61054 658658
rect 60434 658338 60466 658574
rect 60702 658338 60786 658574
rect 61022 658338 61054 658574
rect 60434 657000 61054 658338
rect 61834 707718 62454 707750
rect 61834 707482 61866 707718
rect 62102 707482 62186 707718
rect 62422 707482 62454 707718
rect 61834 707398 62454 707482
rect 61834 707162 61866 707398
rect 62102 707162 62186 707398
rect 62422 707162 62454 707398
rect 61834 673174 62454 707162
rect 61834 672938 61866 673174
rect 62102 672938 62186 673174
rect 62422 672938 62454 673174
rect 61834 672854 62454 672938
rect 61834 672618 61866 672854
rect 62102 672618 62186 672854
rect 62422 672618 62454 672854
rect 61834 657000 62454 672618
rect 63234 704838 63854 705830
rect 63234 704602 63266 704838
rect 63502 704602 63586 704838
rect 63822 704602 63854 704838
rect 63234 704518 63854 704602
rect 63234 704282 63266 704518
rect 63502 704282 63586 704518
rect 63822 704282 63854 704518
rect 63234 687454 63854 704282
rect 63234 687218 63266 687454
rect 63502 687218 63586 687454
rect 63822 687218 63854 687454
rect 63234 687134 63854 687218
rect 63234 686898 63266 687134
rect 63502 686898 63586 687134
rect 63822 686898 63854 687134
rect 63234 657000 63854 686898
rect 64154 698614 64774 710042
rect 69274 711558 69894 711590
rect 69274 711322 69306 711558
rect 69542 711322 69626 711558
rect 69862 711322 69894 711558
rect 69274 711238 69894 711322
rect 69274 711002 69306 711238
rect 69542 711002 69626 711238
rect 69862 711002 69894 711238
rect 64154 698378 64186 698614
rect 64422 698378 64506 698614
rect 64742 698378 64774 698614
rect 64154 698294 64774 698378
rect 64154 698058 64186 698294
rect 64422 698058 64506 698294
rect 64742 698058 64774 698294
rect 64154 662614 64774 698058
rect 64154 662378 64186 662614
rect 64422 662378 64506 662614
rect 64742 662378 64774 662614
rect 64154 662294 64774 662378
rect 64154 662058 64186 662294
rect 64422 662058 64506 662294
rect 64742 662058 64774 662294
rect 64154 657000 64774 662058
rect 65554 709638 66174 709670
rect 65554 709402 65586 709638
rect 65822 709402 65906 709638
rect 66142 709402 66174 709638
rect 65554 709318 66174 709402
rect 65554 709082 65586 709318
rect 65822 709082 65906 709318
rect 66142 709082 66174 709318
rect 65554 676894 66174 709082
rect 65554 676658 65586 676894
rect 65822 676658 65906 676894
rect 66142 676658 66174 676894
rect 65554 676574 66174 676658
rect 65554 676338 65586 676574
rect 65822 676338 65906 676574
rect 66142 676338 66174 676574
rect 65554 657000 66174 676338
rect 66954 706758 67574 707750
rect 66954 706522 66986 706758
rect 67222 706522 67306 706758
rect 67542 706522 67574 706758
rect 66954 706438 67574 706522
rect 66954 706202 66986 706438
rect 67222 706202 67306 706438
rect 67542 706202 67574 706438
rect 66954 691174 67574 706202
rect 66954 690938 66986 691174
rect 67222 690938 67306 691174
rect 67542 690938 67574 691174
rect 66954 690854 67574 690938
rect 66954 690618 66986 690854
rect 67222 690618 67306 690854
rect 67542 690618 67574 690854
rect 66954 657000 67574 690618
rect 68354 705798 68974 705830
rect 68354 705562 68386 705798
rect 68622 705562 68706 705798
rect 68942 705562 68974 705798
rect 68354 705478 68974 705562
rect 68354 705242 68386 705478
rect 68622 705242 68706 705478
rect 68942 705242 68974 705478
rect 68354 669454 68974 705242
rect 68354 669218 68386 669454
rect 68622 669218 68706 669454
rect 68942 669218 68974 669454
rect 68354 669134 68974 669218
rect 68354 668898 68386 669134
rect 68622 668898 68706 669134
rect 68942 668898 68974 669134
rect 68354 657000 68974 668898
rect 69274 680614 69894 711002
rect 74394 710598 75014 711590
rect 74394 710362 74426 710598
rect 74662 710362 74746 710598
rect 74982 710362 75014 710598
rect 74394 710278 75014 710362
rect 74394 710042 74426 710278
rect 74662 710042 74746 710278
rect 74982 710042 75014 710278
rect 69274 680378 69306 680614
rect 69542 680378 69626 680614
rect 69862 680378 69894 680614
rect 69274 680294 69894 680378
rect 69274 680058 69306 680294
rect 69542 680058 69626 680294
rect 69862 680058 69894 680294
rect 69274 657000 69894 680058
rect 70674 708678 71294 709670
rect 70674 708442 70706 708678
rect 70942 708442 71026 708678
rect 71262 708442 71294 708678
rect 70674 708358 71294 708442
rect 70674 708122 70706 708358
rect 70942 708122 71026 708358
rect 71262 708122 71294 708358
rect 70674 694894 71294 708122
rect 70674 694658 70706 694894
rect 70942 694658 71026 694894
rect 71262 694658 71294 694894
rect 70674 694574 71294 694658
rect 70674 694338 70706 694574
rect 70942 694338 71026 694574
rect 71262 694338 71294 694574
rect 70674 658894 71294 694338
rect 70674 658658 70706 658894
rect 70942 658658 71026 658894
rect 71262 658658 71294 658894
rect 70674 658574 71294 658658
rect 70674 658338 70706 658574
rect 70942 658338 71026 658574
rect 71262 658338 71294 658574
rect 70674 657000 71294 658338
rect 72074 707718 72694 707750
rect 72074 707482 72106 707718
rect 72342 707482 72426 707718
rect 72662 707482 72694 707718
rect 72074 707398 72694 707482
rect 72074 707162 72106 707398
rect 72342 707162 72426 707398
rect 72662 707162 72694 707398
rect 72074 673174 72694 707162
rect 72074 672938 72106 673174
rect 72342 672938 72426 673174
rect 72662 672938 72694 673174
rect 72074 672854 72694 672938
rect 72074 672618 72106 672854
rect 72342 672618 72426 672854
rect 72662 672618 72694 672854
rect 72074 657000 72694 672618
rect 73474 704838 74094 705830
rect 73474 704602 73506 704838
rect 73742 704602 73826 704838
rect 74062 704602 74094 704838
rect 73474 704518 74094 704602
rect 73474 704282 73506 704518
rect 73742 704282 73826 704518
rect 74062 704282 74094 704518
rect 73474 687454 74094 704282
rect 73474 687218 73506 687454
rect 73742 687218 73826 687454
rect 74062 687218 74094 687454
rect 73474 687134 74094 687218
rect 73474 686898 73506 687134
rect 73742 686898 73826 687134
rect 74062 686898 74094 687134
rect 73474 657000 74094 686898
rect 74394 698614 75014 710042
rect 79514 711558 80134 711590
rect 79514 711322 79546 711558
rect 79782 711322 79866 711558
rect 80102 711322 80134 711558
rect 79514 711238 80134 711322
rect 79514 711002 79546 711238
rect 79782 711002 79866 711238
rect 80102 711002 80134 711238
rect 74394 698378 74426 698614
rect 74662 698378 74746 698614
rect 74982 698378 75014 698614
rect 74394 698294 75014 698378
rect 74394 698058 74426 698294
rect 74662 698058 74746 698294
rect 74982 698058 75014 698294
rect 74394 662614 75014 698058
rect 74394 662378 74426 662614
rect 74662 662378 74746 662614
rect 74982 662378 75014 662614
rect 74394 662294 75014 662378
rect 74394 662058 74426 662294
rect 74662 662058 74746 662294
rect 74982 662058 75014 662294
rect 74394 657000 75014 662058
rect 75794 709638 76414 709670
rect 75794 709402 75826 709638
rect 76062 709402 76146 709638
rect 76382 709402 76414 709638
rect 75794 709318 76414 709402
rect 75794 709082 75826 709318
rect 76062 709082 76146 709318
rect 76382 709082 76414 709318
rect 75794 676894 76414 709082
rect 75794 676658 75826 676894
rect 76062 676658 76146 676894
rect 76382 676658 76414 676894
rect 75794 676574 76414 676658
rect 75794 676338 75826 676574
rect 76062 676338 76146 676574
rect 76382 676338 76414 676574
rect 75794 657000 76414 676338
rect 77194 706758 77814 707750
rect 77194 706522 77226 706758
rect 77462 706522 77546 706758
rect 77782 706522 77814 706758
rect 77194 706438 77814 706522
rect 77194 706202 77226 706438
rect 77462 706202 77546 706438
rect 77782 706202 77814 706438
rect 77194 691174 77814 706202
rect 77194 690938 77226 691174
rect 77462 690938 77546 691174
rect 77782 690938 77814 691174
rect 77194 690854 77814 690938
rect 77194 690618 77226 690854
rect 77462 690618 77546 690854
rect 77782 690618 77814 690854
rect 77194 657000 77814 690618
rect 78594 705798 79214 705830
rect 78594 705562 78626 705798
rect 78862 705562 78946 705798
rect 79182 705562 79214 705798
rect 78594 705478 79214 705562
rect 78594 705242 78626 705478
rect 78862 705242 78946 705478
rect 79182 705242 79214 705478
rect 78594 669454 79214 705242
rect 78594 669218 78626 669454
rect 78862 669218 78946 669454
rect 79182 669218 79214 669454
rect 78594 669134 79214 669218
rect 78594 668898 78626 669134
rect 78862 668898 78946 669134
rect 79182 668898 79214 669134
rect 78594 657000 79214 668898
rect 79514 680614 80134 711002
rect 84634 710598 85254 711590
rect 84634 710362 84666 710598
rect 84902 710362 84986 710598
rect 85222 710362 85254 710598
rect 84634 710278 85254 710362
rect 84634 710042 84666 710278
rect 84902 710042 84986 710278
rect 85222 710042 85254 710278
rect 79514 680378 79546 680614
rect 79782 680378 79866 680614
rect 80102 680378 80134 680614
rect 79514 680294 80134 680378
rect 79514 680058 79546 680294
rect 79782 680058 79866 680294
rect 80102 680058 80134 680294
rect 79514 657000 80134 680058
rect 80914 708678 81534 709670
rect 80914 708442 80946 708678
rect 81182 708442 81266 708678
rect 81502 708442 81534 708678
rect 80914 708358 81534 708442
rect 80914 708122 80946 708358
rect 81182 708122 81266 708358
rect 81502 708122 81534 708358
rect 80914 694894 81534 708122
rect 80914 694658 80946 694894
rect 81182 694658 81266 694894
rect 81502 694658 81534 694894
rect 80914 694574 81534 694658
rect 80914 694338 80946 694574
rect 81182 694338 81266 694574
rect 81502 694338 81534 694574
rect 80914 658894 81534 694338
rect 80914 658658 80946 658894
rect 81182 658658 81266 658894
rect 81502 658658 81534 658894
rect 80914 658574 81534 658658
rect 80914 658338 80946 658574
rect 81182 658338 81266 658574
rect 81502 658338 81534 658574
rect 80914 657000 81534 658338
rect 82314 707718 82934 707750
rect 82314 707482 82346 707718
rect 82582 707482 82666 707718
rect 82902 707482 82934 707718
rect 82314 707398 82934 707482
rect 82314 707162 82346 707398
rect 82582 707162 82666 707398
rect 82902 707162 82934 707398
rect 82314 673174 82934 707162
rect 82314 672938 82346 673174
rect 82582 672938 82666 673174
rect 82902 672938 82934 673174
rect 82314 672854 82934 672938
rect 82314 672618 82346 672854
rect 82582 672618 82666 672854
rect 82902 672618 82934 672854
rect 82314 657000 82934 672618
rect 83714 704838 84334 705830
rect 83714 704602 83746 704838
rect 83982 704602 84066 704838
rect 84302 704602 84334 704838
rect 83714 704518 84334 704602
rect 83714 704282 83746 704518
rect 83982 704282 84066 704518
rect 84302 704282 84334 704518
rect 83714 687454 84334 704282
rect 83714 687218 83746 687454
rect 83982 687218 84066 687454
rect 84302 687218 84334 687454
rect 83714 687134 84334 687218
rect 83714 686898 83746 687134
rect 83982 686898 84066 687134
rect 84302 686898 84334 687134
rect 83714 657000 84334 686898
rect 84634 698614 85254 710042
rect 89754 711558 90374 711590
rect 89754 711322 89786 711558
rect 90022 711322 90106 711558
rect 90342 711322 90374 711558
rect 89754 711238 90374 711322
rect 89754 711002 89786 711238
rect 90022 711002 90106 711238
rect 90342 711002 90374 711238
rect 84634 698378 84666 698614
rect 84902 698378 84986 698614
rect 85222 698378 85254 698614
rect 84634 698294 85254 698378
rect 84634 698058 84666 698294
rect 84902 698058 84986 698294
rect 85222 698058 85254 698294
rect 84634 662614 85254 698058
rect 84634 662378 84666 662614
rect 84902 662378 84986 662614
rect 85222 662378 85254 662614
rect 84634 662294 85254 662378
rect 84634 662058 84666 662294
rect 84902 662058 84986 662294
rect 85222 662058 85254 662294
rect 84634 657000 85254 662058
rect 86034 709638 86654 709670
rect 86034 709402 86066 709638
rect 86302 709402 86386 709638
rect 86622 709402 86654 709638
rect 86034 709318 86654 709402
rect 86034 709082 86066 709318
rect 86302 709082 86386 709318
rect 86622 709082 86654 709318
rect 86034 676894 86654 709082
rect 86034 676658 86066 676894
rect 86302 676658 86386 676894
rect 86622 676658 86654 676894
rect 86034 676574 86654 676658
rect 86034 676338 86066 676574
rect 86302 676338 86386 676574
rect 86622 676338 86654 676574
rect 86034 657000 86654 676338
rect 87434 706758 88054 707750
rect 87434 706522 87466 706758
rect 87702 706522 87786 706758
rect 88022 706522 88054 706758
rect 87434 706438 88054 706522
rect 87434 706202 87466 706438
rect 87702 706202 87786 706438
rect 88022 706202 88054 706438
rect 87434 691174 88054 706202
rect 87434 690938 87466 691174
rect 87702 690938 87786 691174
rect 88022 690938 88054 691174
rect 87434 690854 88054 690938
rect 87434 690618 87466 690854
rect 87702 690618 87786 690854
rect 88022 690618 88054 690854
rect 87434 657000 88054 690618
rect 88834 705798 89454 705830
rect 88834 705562 88866 705798
rect 89102 705562 89186 705798
rect 89422 705562 89454 705798
rect 88834 705478 89454 705562
rect 88834 705242 88866 705478
rect 89102 705242 89186 705478
rect 89422 705242 89454 705478
rect 88834 669454 89454 705242
rect 88834 669218 88866 669454
rect 89102 669218 89186 669454
rect 89422 669218 89454 669454
rect 88834 669134 89454 669218
rect 88834 668898 88866 669134
rect 89102 668898 89186 669134
rect 89422 668898 89454 669134
rect 88834 657000 89454 668898
rect 89754 680614 90374 711002
rect 94874 710598 95494 711590
rect 94874 710362 94906 710598
rect 95142 710362 95226 710598
rect 95462 710362 95494 710598
rect 94874 710278 95494 710362
rect 94874 710042 94906 710278
rect 95142 710042 95226 710278
rect 95462 710042 95494 710278
rect 89754 680378 89786 680614
rect 90022 680378 90106 680614
rect 90342 680378 90374 680614
rect 89754 680294 90374 680378
rect 89754 680058 89786 680294
rect 90022 680058 90106 680294
rect 90342 680058 90374 680294
rect 89754 657000 90374 680058
rect 91154 708678 91774 709670
rect 91154 708442 91186 708678
rect 91422 708442 91506 708678
rect 91742 708442 91774 708678
rect 91154 708358 91774 708442
rect 91154 708122 91186 708358
rect 91422 708122 91506 708358
rect 91742 708122 91774 708358
rect 91154 694894 91774 708122
rect 91154 694658 91186 694894
rect 91422 694658 91506 694894
rect 91742 694658 91774 694894
rect 91154 694574 91774 694658
rect 91154 694338 91186 694574
rect 91422 694338 91506 694574
rect 91742 694338 91774 694574
rect 91154 658894 91774 694338
rect 91154 658658 91186 658894
rect 91422 658658 91506 658894
rect 91742 658658 91774 658894
rect 91154 658574 91774 658658
rect 91154 658338 91186 658574
rect 91422 658338 91506 658574
rect 91742 658338 91774 658574
rect 91154 657000 91774 658338
rect 92554 707718 93174 707750
rect 92554 707482 92586 707718
rect 92822 707482 92906 707718
rect 93142 707482 93174 707718
rect 92554 707398 93174 707482
rect 92554 707162 92586 707398
rect 92822 707162 92906 707398
rect 93142 707162 93174 707398
rect 92554 673174 93174 707162
rect 92554 672938 92586 673174
rect 92822 672938 92906 673174
rect 93142 672938 93174 673174
rect 92554 672854 93174 672938
rect 92554 672618 92586 672854
rect 92822 672618 92906 672854
rect 93142 672618 93174 672854
rect 92554 657000 93174 672618
rect 93954 704838 94574 705830
rect 93954 704602 93986 704838
rect 94222 704602 94306 704838
rect 94542 704602 94574 704838
rect 93954 704518 94574 704602
rect 93954 704282 93986 704518
rect 94222 704282 94306 704518
rect 94542 704282 94574 704518
rect 93954 687454 94574 704282
rect 93954 687218 93986 687454
rect 94222 687218 94306 687454
rect 94542 687218 94574 687454
rect 93954 687134 94574 687218
rect 93954 686898 93986 687134
rect 94222 686898 94306 687134
rect 94542 686898 94574 687134
rect 93954 657000 94574 686898
rect 94874 698614 95494 710042
rect 99994 711558 100614 711590
rect 99994 711322 100026 711558
rect 100262 711322 100346 711558
rect 100582 711322 100614 711558
rect 99994 711238 100614 711322
rect 99994 711002 100026 711238
rect 100262 711002 100346 711238
rect 100582 711002 100614 711238
rect 94874 698378 94906 698614
rect 95142 698378 95226 698614
rect 95462 698378 95494 698614
rect 94874 698294 95494 698378
rect 94874 698058 94906 698294
rect 95142 698058 95226 698294
rect 95462 698058 95494 698294
rect 94874 662614 95494 698058
rect 94874 662378 94906 662614
rect 95142 662378 95226 662614
rect 95462 662378 95494 662614
rect 94874 662294 95494 662378
rect 94874 662058 94906 662294
rect 95142 662058 95226 662294
rect 95462 662058 95494 662294
rect 94874 657000 95494 662058
rect 96274 709638 96894 709670
rect 96274 709402 96306 709638
rect 96542 709402 96626 709638
rect 96862 709402 96894 709638
rect 96274 709318 96894 709402
rect 96274 709082 96306 709318
rect 96542 709082 96626 709318
rect 96862 709082 96894 709318
rect 96274 676894 96894 709082
rect 96274 676658 96306 676894
rect 96542 676658 96626 676894
rect 96862 676658 96894 676894
rect 96274 676574 96894 676658
rect 96274 676338 96306 676574
rect 96542 676338 96626 676574
rect 96862 676338 96894 676574
rect 96274 657000 96894 676338
rect 97674 706758 98294 707750
rect 97674 706522 97706 706758
rect 97942 706522 98026 706758
rect 98262 706522 98294 706758
rect 97674 706438 98294 706522
rect 97674 706202 97706 706438
rect 97942 706202 98026 706438
rect 98262 706202 98294 706438
rect 97674 691174 98294 706202
rect 97674 690938 97706 691174
rect 97942 690938 98026 691174
rect 98262 690938 98294 691174
rect 97674 690854 98294 690938
rect 97674 690618 97706 690854
rect 97942 690618 98026 690854
rect 98262 690618 98294 690854
rect 97674 657000 98294 690618
rect 99074 705798 99694 705830
rect 99074 705562 99106 705798
rect 99342 705562 99426 705798
rect 99662 705562 99694 705798
rect 99074 705478 99694 705562
rect 99074 705242 99106 705478
rect 99342 705242 99426 705478
rect 99662 705242 99694 705478
rect 99074 669454 99694 705242
rect 99074 669218 99106 669454
rect 99342 669218 99426 669454
rect 99662 669218 99694 669454
rect 99074 669134 99694 669218
rect 99074 668898 99106 669134
rect 99342 668898 99426 669134
rect 99662 668898 99694 669134
rect 99074 657000 99694 668898
rect 99994 680614 100614 711002
rect 105114 710598 105734 711590
rect 105114 710362 105146 710598
rect 105382 710362 105466 710598
rect 105702 710362 105734 710598
rect 105114 710278 105734 710362
rect 105114 710042 105146 710278
rect 105382 710042 105466 710278
rect 105702 710042 105734 710278
rect 99994 680378 100026 680614
rect 100262 680378 100346 680614
rect 100582 680378 100614 680614
rect 99994 680294 100614 680378
rect 99994 680058 100026 680294
rect 100262 680058 100346 680294
rect 100582 680058 100614 680294
rect 99994 657000 100614 680058
rect 101394 708678 102014 709670
rect 101394 708442 101426 708678
rect 101662 708442 101746 708678
rect 101982 708442 102014 708678
rect 101394 708358 102014 708442
rect 101394 708122 101426 708358
rect 101662 708122 101746 708358
rect 101982 708122 102014 708358
rect 101394 694894 102014 708122
rect 101394 694658 101426 694894
rect 101662 694658 101746 694894
rect 101982 694658 102014 694894
rect 101394 694574 102014 694658
rect 101394 694338 101426 694574
rect 101662 694338 101746 694574
rect 101982 694338 102014 694574
rect 101394 658894 102014 694338
rect 101394 658658 101426 658894
rect 101662 658658 101746 658894
rect 101982 658658 102014 658894
rect 101394 658574 102014 658658
rect 101394 658338 101426 658574
rect 101662 658338 101746 658574
rect 101982 658338 102014 658574
rect 101394 657000 102014 658338
rect 102794 707718 103414 707750
rect 102794 707482 102826 707718
rect 103062 707482 103146 707718
rect 103382 707482 103414 707718
rect 102794 707398 103414 707482
rect 102794 707162 102826 707398
rect 103062 707162 103146 707398
rect 103382 707162 103414 707398
rect 102794 673174 103414 707162
rect 102794 672938 102826 673174
rect 103062 672938 103146 673174
rect 103382 672938 103414 673174
rect 102794 672854 103414 672938
rect 102794 672618 102826 672854
rect 103062 672618 103146 672854
rect 103382 672618 103414 672854
rect 102794 657000 103414 672618
rect 104194 704838 104814 705830
rect 104194 704602 104226 704838
rect 104462 704602 104546 704838
rect 104782 704602 104814 704838
rect 104194 704518 104814 704602
rect 104194 704282 104226 704518
rect 104462 704282 104546 704518
rect 104782 704282 104814 704518
rect 104194 687454 104814 704282
rect 104194 687218 104226 687454
rect 104462 687218 104546 687454
rect 104782 687218 104814 687454
rect 104194 687134 104814 687218
rect 104194 686898 104226 687134
rect 104462 686898 104546 687134
rect 104782 686898 104814 687134
rect 104194 657000 104814 686898
rect 105114 698614 105734 710042
rect 110234 711558 110854 711590
rect 110234 711322 110266 711558
rect 110502 711322 110586 711558
rect 110822 711322 110854 711558
rect 110234 711238 110854 711322
rect 110234 711002 110266 711238
rect 110502 711002 110586 711238
rect 110822 711002 110854 711238
rect 105114 698378 105146 698614
rect 105382 698378 105466 698614
rect 105702 698378 105734 698614
rect 105114 698294 105734 698378
rect 105114 698058 105146 698294
rect 105382 698058 105466 698294
rect 105702 698058 105734 698294
rect 105114 662614 105734 698058
rect 105114 662378 105146 662614
rect 105382 662378 105466 662614
rect 105702 662378 105734 662614
rect 105114 662294 105734 662378
rect 105114 662058 105146 662294
rect 105382 662058 105466 662294
rect 105702 662058 105734 662294
rect 105114 657000 105734 662058
rect 106514 709638 107134 709670
rect 106514 709402 106546 709638
rect 106782 709402 106866 709638
rect 107102 709402 107134 709638
rect 106514 709318 107134 709402
rect 106514 709082 106546 709318
rect 106782 709082 106866 709318
rect 107102 709082 107134 709318
rect 106514 676894 107134 709082
rect 106514 676658 106546 676894
rect 106782 676658 106866 676894
rect 107102 676658 107134 676894
rect 106514 676574 107134 676658
rect 106514 676338 106546 676574
rect 106782 676338 106866 676574
rect 107102 676338 107134 676574
rect 106514 657000 107134 676338
rect 107914 706758 108534 707750
rect 107914 706522 107946 706758
rect 108182 706522 108266 706758
rect 108502 706522 108534 706758
rect 107914 706438 108534 706522
rect 107914 706202 107946 706438
rect 108182 706202 108266 706438
rect 108502 706202 108534 706438
rect 107914 691174 108534 706202
rect 107914 690938 107946 691174
rect 108182 690938 108266 691174
rect 108502 690938 108534 691174
rect 107914 690854 108534 690938
rect 107914 690618 107946 690854
rect 108182 690618 108266 690854
rect 108502 690618 108534 690854
rect 107914 657000 108534 690618
rect 109314 705798 109934 705830
rect 109314 705562 109346 705798
rect 109582 705562 109666 705798
rect 109902 705562 109934 705798
rect 109314 705478 109934 705562
rect 109314 705242 109346 705478
rect 109582 705242 109666 705478
rect 109902 705242 109934 705478
rect 109314 669454 109934 705242
rect 109314 669218 109346 669454
rect 109582 669218 109666 669454
rect 109902 669218 109934 669454
rect 109314 669134 109934 669218
rect 109314 668898 109346 669134
rect 109582 668898 109666 669134
rect 109902 668898 109934 669134
rect 109314 657000 109934 668898
rect 110234 680614 110854 711002
rect 115354 710598 115974 711590
rect 115354 710362 115386 710598
rect 115622 710362 115706 710598
rect 115942 710362 115974 710598
rect 115354 710278 115974 710362
rect 115354 710042 115386 710278
rect 115622 710042 115706 710278
rect 115942 710042 115974 710278
rect 110234 680378 110266 680614
rect 110502 680378 110586 680614
rect 110822 680378 110854 680614
rect 110234 680294 110854 680378
rect 110234 680058 110266 680294
rect 110502 680058 110586 680294
rect 110822 680058 110854 680294
rect 110234 657000 110854 680058
rect 111634 708678 112254 709670
rect 111634 708442 111666 708678
rect 111902 708442 111986 708678
rect 112222 708442 112254 708678
rect 111634 708358 112254 708442
rect 111634 708122 111666 708358
rect 111902 708122 111986 708358
rect 112222 708122 112254 708358
rect 111634 694894 112254 708122
rect 111634 694658 111666 694894
rect 111902 694658 111986 694894
rect 112222 694658 112254 694894
rect 111634 694574 112254 694658
rect 111634 694338 111666 694574
rect 111902 694338 111986 694574
rect 112222 694338 112254 694574
rect 111634 658894 112254 694338
rect 111634 658658 111666 658894
rect 111902 658658 111986 658894
rect 112222 658658 112254 658894
rect 111634 658574 112254 658658
rect 111634 658338 111666 658574
rect 111902 658338 111986 658574
rect 112222 658338 112254 658574
rect 111634 657000 112254 658338
rect 113034 707718 113654 707750
rect 113034 707482 113066 707718
rect 113302 707482 113386 707718
rect 113622 707482 113654 707718
rect 113034 707398 113654 707482
rect 113034 707162 113066 707398
rect 113302 707162 113386 707398
rect 113622 707162 113654 707398
rect 113034 673174 113654 707162
rect 113034 672938 113066 673174
rect 113302 672938 113386 673174
rect 113622 672938 113654 673174
rect 113034 672854 113654 672938
rect 113034 672618 113066 672854
rect 113302 672618 113386 672854
rect 113622 672618 113654 672854
rect 113034 657000 113654 672618
rect 114434 704838 115054 705830
rect 114434 704602 114466 704838
rect 114702 704602 114786 704838
rect 115022 704602 115054 704838
rect 114434 704518 115054 704602
rect 114434 704282 114466 704518
rect 114702 704282 114786 704518
rect 115022 704282 115054 704518
rect 114434 687454 115054 704282
rect 114434 687218 114466 687454
rect 114702 687218 114786 687454
rect 115022 687218 115054 687454
rect 114434 687134 115054 687218
rect 114434 686898 114466 687134
rect 114702 686898 114786 687134
rect 115022 686898 115054 687134
rect 114434 657000 115054 686898
rect 115354 698614 115974 710042
rect 120474 711558 121094 711590
rect 120474 711322 120506 711558
rect 120742 711322 120826 711558
rect 121062 711322 121094 711558
rect 120474 711238 121094 711322
rect 120474 711002 120506 711238
rect 120742 711002 120826 711238
rect 121062 711002 121094 711238
rect 115354 698378 115386 698614
rect 115622 698378 115706 698614
rect 115942 698378 115974 698614
rect 115354 698294 115974 698378
rect 115354 698058 115386 698294
rect 115622 698058 115706 698294
rect 115942 698058 115974 698294
rect 115354 662614 115974 698058
rect 115354 662378 115386 662614
rect 115622 662378 115706 662614
rect 115942 662378 115974 662614
rect 115354 662294 115974 662378
rect 115354 662058 115386 662294
rect 115622 662058 115706 662294
rect 115942 662058 115974 662294
rect 115354 657000 115974 662058
rect 116754 709638 117374 709670
rect 116754 709402 116786 709638
rect 117022 709402 117106 709638
rect 117342 709402 117374 709638
rect 116754 709318 117374 709402
rect 116754 709082 116786 709318
rect 117022 709082 117106 709318
rect 117342 709082 117374 709318
rect 116754 676894 117374 709082
rect 116754 676658 116786 676894
rect 117022 676658 117106 676894
rect 117342 676658 117374 676894
rect 116754 676574 117374 676658
rect 116754 676338 116786 676574
rect 117022 676338 117106 676574
rect 117342 676338 117374 676574
rect 116754 657000 117374 676338
rect 118154 706758 118774 707750
rect 118154 706522 118186 706758
rect 118422 706522 118506 706758
rect 118742 706522 118774 706758
rect 118154 706438 118774 706522
rect 118154 706202 118186 706438
rect 118422 706202 118506 706438
rect 118742 706202 118774 706438
rect 118154 691174 118774 706202
rect 118154 690938 118186 691174
rect 118422 690938 118506 691174
rect 118742 690938 118774 691174
rect 118154 690854 118774 690938
rect 118154 690618 118186 690854
rect 118422 690618 118506 690854
rect 118742 690618 118774 690854
rect 118154 657000 118774 690618
rect 119554 705798 120174 705830
rect 119554 705562 119586 705798
rect 119822 705562 119906 705798
rect 120142 705562 120174 705798
rect 119554 705478 120174 705562
rect 119554 705242 119586 705478
rect 119822 705242 119906 705478
rect 120142 705242 120174 705478
rect 119554 669454 120174 705242
rect 119554 669218 119586 669454
rect 119822 669218 119906 669454
rect 120142 669218 120174 669454
rect 119554 669134 120174 669218
rect 119554 668898 119586 669134
rect 119822 668898 119906 669134
rect 120142 668898 120174 669134
rect 119554 657000 120174 668898
rect 120474 680614 121094 711002
rect 125594 710598 126214 711590
rect 125594 710362 125626 710598
rect 125862 710362 125946 710598
rect 126182 710362 126214 710598
rect 125594 710278 126214 710362
rect 125594 710042 125626 710278
rect 125862 710042 125946 710278
rect 126182 710042 126214 710278
rect 120474 680378 120506 680614
rect 120742 680378 120826 680614
rect 121062 680378 121094 680614
rect 120474 680294 121094 680378
rect 120474 680058 120506 680294
rect 120742 680058 120826 680294
rect 121062 680058 121094 680294
rect 120474 657000 121094 680058
rect 121874 708678 122494 709670
rect 121874 708442 121906 708678
rect 122142 708442 122226 708678
rect 122462 708442 122494 708678
rect 121874 708358 122494 708442
rect 121874 708122 121906 708358
rect 122142 708122 122226 708358
rect 122462 708122 122494 708358
rect 121874 694894 122494 708122
rect 121874 694658 121906 694894
rect 122142 694658 122226 694894
rect 122462 694658 122494 694894
rect 121874 694574 122494 694658
rect 121874 694338 121906 694574
rect 122142 694338 122226 694574
rect 122462 694338 122494 694574
rect 121874 658894 122494 694338
rect 121874 658658 121906 658894
rect 122142 658658 122226 658894
rect 122462 658658 122494 658894
rect 121874 658574 122494 658658
rect 121874 658338 121906 658574
rect 122142 658338 122226 658574
rect 122462 658338 122494 658574
rect 121874 657000 122494 658338
rect 123274 707718 123894 707750
rect 123274 707482 123306 707718
rect 123542 707482 123626 707718
rect 123862 707482 123894 707718
rect 123274 707398 123894 707482
rect 123274 707162 123306 707398
rect 123542 707162 123626 707398
rect 123862 707162 123894 707398
rect 123274 673174 123894 707162
rect 123274 672938 123306 673174
rect 123542 672938 123626 673174
rect 123862 672938 123894 673174
rect 123274 672854 123894 672938
rect 123274 672618 123306 672854
rect 123542 672618 123626 672854
rect 123862 672618 123894 672854
rect 123274 657000 123894 672618
rect 124674 704838 125294 705830
rect 124674 704602 124706 704838
rect 124942 704602 125026 704838
rect 125262 704602 125294 704838
rect 124674 704518 125294 704602
rect 124674 704282 124706 704518
rect 124942 704282 125026 704518
rect 125262 704282 125294 704518
rect 124674 687454 125294 704282
rect 124674 687218 124706 687454
rect 124942 687218 125026 687454
rect 125262 687218 125294 687454
rect 124674 687134 125294 687218
rect 124674 686898 124706 687134
rect 124942 686898 125026 687134
rect 125262 686898 125294 687134
rect 124674 657000 125294 686898
rect 125594 698614 126214 710042
rect 130714 711558 131334 711590
rect 130714 711322 130746 711558
rect 130982 711322 131066 711558
rect 131302 711322 131334 711558
rect 130714 711238 131334 711322
rect 130714 711002 130746 711238
rect 130982 711002 131066 711238
rect 131302 711002 131334 711238
rect 125594 698378 125626 698614
rect 125862 698378 125946 698614
rect 126182 698378 126214 698614
rect 125594 698294 126214 698378
rect 125594 698058 125626 698294
rect 125862 698058 125946 698294
rect 126182 698058 126214 698294
rect 125594 662614 126214 698058
rect 125594 662378 125626 662614
rect 125862 662378 125946 662614
rect 126182 662378 126214 662614
rect 125594 662294 126214 662378
rect 125594 662058 125626 662294
rect 125862 662058 125946 662294
rect 126182 662058 126214 662294
rect 125594 657000 126214 662058
rect 126994 709638 127614 709670
rect 126994 709402 127026 709638
rect 127262 709402 127346 709638
rect 127582 709402 127614 709638
rect 126994 709318 127614 709402
rect 126994 709082 127026 709318
rect 127262 709082 127346 709318
rect 127582 709082 127614 709318
rect 126994 676894 127614 709082
rect 126994 676658 127026 676894
rect 127262 676658 127346 676894
rect 127582 676658 127614 676894
rect 126994 676574 127614 676658
rect 126994 676338 127026 676574
rect 127262 676338 127346 676574
rect 127582 676338 127614 676574
rect 126994 657000 127614 676338
rect 128394 706758 129014 707750
rect 128394 706522 128426 706758
rect 128662 706522 128746 706758
rect 128982 706522 129014 706758
rect 128394 706438 129014 706522
rect 128394 706202 128426 706438
rect 128662 706202 128746 706438
rect 128982 706202 129014 706438
rect 128394 691174 129014 706202
rect 128394 690938 128426 691174
rect 128662 690938 128746 691174
rect 128982 690938 129014 691174
rect 128394 690854 129014 690938
rect 128394 690618 128426 690854
rect 128662 690618 128746 690854
rect 128982 690618 129014 690854
rect 128394 657000 129014 690618
rect 129794 705798 130414 705830
rect 129794 705562 129826 705798
rect 130062 705562 130146 705798
rect 130382 705562 130414 705798
rect 129794 705478 130414 705562
rect 129794 705242 129826 705478
rect 130062 705242 130146 705478
rect 130382 705242 130414 705478
rect 129794 669454 130414 705242
rect 129794 669218 129826 669454
rect 130062 669218 130146 669454
rect 130382 669218 130414 669454
rect 129794 669134 130414 669218
rect 129794 668898 129826 669134
rect 130062 668898 130146 669134
rect 130382 668898 130414 669134
rect 129794 657000 130414 668898
rect 130714 680614 131334 711002
rect 135834 710598 136454 711590
rect 135834 710362 135866 710598
rect 136102 710362 136186 710598
rect 136422 710362 136454 710598
rect 135834 710278 136454 710362
rect 135834 710042 135866 710278
rect 136102 710042 136186 710278
rect 136422 710042 136454 710278
rect 130714 680378 130746 680614
rect 130982 680378 131066 680614
rect 131302 680378 131334 680614
rect 130714 680294 131334 680378
rect 130714 680058 130746 680294
rect 130982 680058 131066 680294
rect 131302 680058 131334 680294
rect 130714 657000 131334 680058
rect 132114 708678 132734 709670
rect 132114 708442 132146 708678
rect 132382 708442 132466 708678
rect 132702 708442 132734 708678
rect 132114 708358 132734 708442
rect 132114 708122 132146 708358
rect 132382 708122 132466 708358
rect 132702 708122 132734 708358
rect 132114 694894 132734 708122
rect 132114 694658 132146 694894
rect 132382 694658 132466 694894
rect 132702 694658 132734 694894
rect 132114 694574 132734 694658
rect 132114 694338 132146 694574
rect 132382 694338 132466 694574
rect 132702 694338 132734 694574
rect 132114 658894 132734 694338
rect 132114 658658 132146 658894
rect 132382 658658 132466 658894
rect 132702 658658 132734 658894
rect 132114 658574 132734 658658
rect 132114 658338 132146 658574
rect 132382 658338 132466 658574
rect 132702 658338 132734 658574
rect 132114 657000 132734 658338
rect 133514 707718 134134 707750
rect 133514 707482 133546 707718
rect 133782 707482 133866 707718
rect 134102 707482 134134 707718
rect 133514 707398 134134 707482
rect 133514 707162 133546 707398
rect 133782 707162 133866 707398
rect 134102 707162 134134 707398
rect 133514 673174 134134 707162
rect 133514 672938 133546 673174
rect 133782 672938 133866 673174
rect 134102 672938 134134 673174
rect 133514 672854 134134 672938
rect 133514 672618 133546 672854
rect 133782 672618 133866 672854
rect 134102 672618 134134 672854
rect 133514 657000 134134 672618
rect 134914 704838 135534 705830
rect 134914 704602 134946 704838
rect 135182 704602 135266 704838
rect 135502 704602 135534 704838
rect 134914 704518 135534 704602
rect 134914 704282 134946 704518
rect 135182 704282 135266 704518
rect 135502 704282 135534 704518
rect 134914 687454 135534 704282
rect 134914 687218 134946 687454
rect 135182 687218 135266 687454
rect 135502 687218 135534 687454
rect 134914 687134 135534 687218
rect 134914 686898 134946 687134
rect 135182 686898 135266 687134
rect 135502 686898 135534 687134
rect 134914 657000 135534 686898
rect 135834 698614 136454 710042
rect 140954 711558 141574 711590
rect 140954 711322 140986 711558
rect 141222 711322 141306 711558
rect 141542 711322 141574 711558
rect 140954 711238 141574 711322
rect 140954 711002 140986 711238
rect 141222 711002 141306 711238
rect 141542 711002 141574 711238
rect 135834 698378 135866 698614
rect 136102 698378 136186 698614
rect 136422 698378 136454 698614
rect 135834 698294 136454 698378
rect 135834 698058 135866 698294
rect 136102 698058 136186 698294
rect 136422 698058 136454 698294
rect 135834 662614 136454 698058
rect 135834 662378 135866 662614
rect 136102 662378 136186 662614
rect 136422 662378 136454 662614
rect 135834 662294 136454 662378
rect 135834 662058 135866 662294
rect 136102 662058 136186 662294
rect 136422 662058 136454 662294
rect 135834 657000 136454 662058
rect 137234 709638 137854 709670
rect 137234 709402 137266 709638
rect 137502 709402 137586 709638
rect 137822 709402 137854 709638
rect 137234 709318 137854 709402
rect 137234 709082 137266 709318
rect 137502 709082 137586 709318
rect 137822 709082 137854 709318
rect 137234 676894 137854 709082
rect 137234 676658 137266 676894
rect 137502 676658 137586 676894
rect 137822 676658 137854 676894
rect 137234 676574 137854 676658
rect 137234 676338 137266 676574
rect 137502 676338 137586 676574
rect 137822 676338 137854 676574
rect 137234 657000 137854 676338
rect 138634 706758 139254 707750
rect 138634 706522 138666 706758
rect 138902 706522 138986 706758
rect 139222 706522 139254 706758
rect 138634 706438 139254 706522
rect 138634 706202 138666 706438
rect 138902 706202 138986 706438
rect 139222 706202 139254 706438
rect 138634 691174 139254 706202
rect 138634 690938 138666 691174
rect 138902 690938 138986 691174
rect 139222 690938 139254 691174
rect 138634 690854 139254 690938
rect 138634 690618 138666 690854
rect 138902 690618 138986 690854
rect 139222 690618 139254 690854
rect 138634 657000 139254 690618
rect 140034 705798 140654 705830
rect 140034 705562 140066 705798
rect 140302 705562 140386 705798
rect 140622 705562 140654 705798
rect 140034 705478 140654 705562
rect 140034 705242 140066 705478
rect 140302 705242 140386 705478
rect 140622 705242 140654 705478
rect 140034 669454 140654 705242
rect 140034 669218 140066 669454
rect 140302 669218 140386 669454
rect 140622 669218 140654 669454
rect 140034 669134 140654 669218
rect 140034 668898 140066 669134
rect 140302 668898 140386 669134
rect 140622 668898 140654 669134
rect 140034 657000 140654 668898
rect 140954 680614 141574 711002
rect 146074 710598 146694 711590
rect 146074 710362 146106 710598
rect 146342 710362 146426 710598
rect 146662 710362 146694 710598
rect 146074 710278 146694 710362
rect 146074 710042 146106 710278
rect 146342 710042 146426 710278
rect 146662 710042 146694 710278
rect 140954 680378 140986 680614
rect 141222 680378 141306 680614
rect 141542 680378 141574 680614
rect 140954 680294 141574 680378
rect 140954 680058 140986 680294
rect 141222 680058 141306 680294
rect 141542 680058 141574 680294
rect 140954 657000 141574 680058
rect 142354 708678 142974 709670
rect 142354 708442 142386 708678
rect 142622 708442 142706 708678
rect 142942 708442 142974 708678
rect 142354 708358 142974 708442
rect 142354 708122 142386 708358
rect 142622 708122 142706 708358
rect 142942 708122 142974 708358
rect 142354 694894 142974 708122
rect 142354 694658 142386 694894
rect 142622 694658 142706 694894
rect 142942 694658 142974 694894
rect 142354 694574 142974 694658
rect 142354 694338 142386 694574
rect 142622 694338 142706 694574
rect 142942 694338 142974 694574
rect 142354 658894 142974 694338
rect 142354 658658 142386 658894
rect 142622 658658 142706 658894
rect 142942 658658 142974 658894
rect 142354 658574 142974 658658
rect 142354 658338 142386 658574
rect 142622 658338 142706 658574
rect 142942 658338 142974 658574
rect 142354 657000 142974 658338
rect 143754 707718 144374 707750
rect 143754 707482 143786 707718
rect 144022 707482 144106 707718
rect 144342 707482 144374 707718
rect 143754 707398 144374 707482
rect 143754 707162 143786 707398
rect 144022 707162 144106 707398
rect 144342 707162 144374 707398
rect 143754 673174 144374 707162
rect 143754 672938 143786 673174
rect 144022 672938 144106 673174
rect 144342 672938 144374 673174
rect 143754 672854 144374 672938
rect 143754 672618 143786 672854
rect 144022 672618 144106 672854
rect 144342 672618 144374 672854
rect 143754 657000 144374 672618
rect 145154 704838 145774 705830
rect 145154 704602 145186 704838
rect 145422 704602 145506 704838
rect 145742 704602 145774 704838
rect 145154 704518 145774 704602
rect 145154 704282 145186 704518
rect 145422 704282 145506 704518
rect 145742 704282 145774 704518
rect 145154 687454 145774 704282
rect 145154 687218 145186 687454
rect 145422 687218 145506 687454
rect 145742 687218 145774 687454
rect 145154 687134 145774 687218
rect 145154 686898 145186 687134
rect 145422 686898 145506 687134
rect 145742 686898 145774 687134
rect 145154 657000 145774 686898
rect 146074 698614 146694 710042
rect 151194 711558 151814 711590
rect 151194 711322 151226 711558
rect 151462 711322 151546 711558
rect 151782 711322 151814 711558
rect 151194 711238 151814 711322
rect 151194 711002 151226 711238
rect 151462 711002 151546 711238
rect 151782 711002 151814 711238
rect 146074 698378 146106 698614
rect 146342 698378 146426 698614
rect 146662 698378 146694 698614
rect 146074 698294 146694 698378
rect 146074 698058 146106 698294
rect 146342 698058 146426 698294
rect 146662 698058 146694 698294
rect 146074 662614 146694 698058
rect 146074 662378 146106 662614
rect 146342 662378 146426 662614
rect 146662 662378 146694 662614
rect 146074 662294 146694 662378
rect 146074 662058 146106 662294
rect 146342 662058 146426 662294
rect 146662 662058 146694 662294
rect 146074 657000 146694 662058
rect 147474 709638 148094 709670
rect 147474 709402 147506 709638
rect 147742 709402 147826 709638
rect 148062 709402 148094 709638
rect 147474 709318 148094 709402
rect 147474 709082 147506 709318
rect 147742 709082 147826 709318
rect 148062 709082 148094 709318
rect 147474 676894 148094 709082
rect 147474 676658 147506 676894
rect 147742 676658 147826 676894
rect 148062 676658 148094 676894
rect 147474 676574 148094 676658
rect 147474 676338 147506 676574
rect 147742 676338 147826 676574
rect 148062 676338 148094 676574
rect 147474 657000 148094 676338
rect 148874 706758 149494 707750
rect 148874 706522 148906 706758
rect 149142 706522 149226 706758
rect 149462 706522 149494 706758
rect 148874 706438 149494 706522
rect 148874 706202 148906 706438
rect 149142 706202 149226 706438
rect 149462 706202 149494 706438
rect 148874 691174 149494 706202
rect 148874 690938 148906 691174
rect 149142 690938 149226 691174
rect 149462 690938 149494 691174
rect 148874 690854 149494 690938
rect 148874 690618 148906 690854
rect 149142 690618 149226 690854
rect 149462 690618 149494 690854
rect 148874 657000 149494 690618
rect 150274 705798 150894 705830
rect 150274 705562 150306 705798
rect 150542 705562 150626 705798
rect 150862 705562 150894 705798
rect 150274 705478 150894 705562
rect 150274 705242 150306 705478
rect 150542 705242 150626 705478
rect 150862 705242 150894 705478
rect 150274 669454 150894 705242
rect 150274 669218 150306 669454
rect 150542 669218 150626 669454
rect 150862 669218 150894 669454
rect 150274 669134 150894 669218
rect 150274 668898 150306 669134
rect 150542 668898 150626 669134
rect 150862 668898 150894 669134
rect 150274 657000 150894 668898
rect 151194 680614 151814 711002
rect 156314 710598 156934 711590
rect 156314 710362 156346 710598
rect 156582 710362 156666 710598
rect 156902 710362 156934 710598
rect 156314 710278 156934 710362
rect 156314 710042 156346 710278
rect 156582 710042 156666 710278
rect 156902 710042 156934 710278
rect 151194 680378 151226 680614
rect 151462 680378 151546 680614
rect 151782 680378 151814 680614
rect 151194 680294 151814 680378
rect 151194 680058 151226 680294
rect 151462 680058 151546 680294
rect 151782 680058 151814 680294
rect 151194 657000 151814 680058
rect 152594 708678 153214 709670
rect 152594 708442 152626 708678
rect 152862 708442 152946 708678
rect 153182 708442 153214 708678
rect 152594 708358 153214 708442
rect 152594 708122 152626 708358
rect 152862 708122 152946 708358
rect 153182 708122 153214 708358
rect 152594 694894 153214 708122
rect 152594 694658 152626 694894
rect 152862 694658 152946 694894
rect 153182 694658 153214 694894
rect 152594 694574 153214 694658
rect 152594 694338 152626 694574
rect 152862 694338 152946 694574
rect 153182 694338 153214 694574
rect 152594 658894 153214 694338
rect 152594 658658 152626 658894
rect 152862 658658 152946 658894
rect 153182 658658 153214 658894
rect 152594 658574 153214 658658
rect 152594 658338 152626 658574
rect 152862 658338 152946 658574
rect 153182 658338 153214 658574
rect 152594 657000 153214 658338
rect 153994 707718 154614 707750
rect 153994 707482 154026 707718
rect 154262 707482 154346 707718
rect 154582 707482 154614 707718
rect 153994 707398 154614 707482
rect 153994 707162 154026 707398
rect 154262 707162 154346 707398
rect 154582 707162 154614 707398
rect 153994 673174 154614 707162
rect 153994 672938 154026 673174
rect 154262 672938 154346 673174
rect 154582 672938 154614 673174
rect 153994 672854 154614 672938
rect 153994 672618 154026 672854
rect 154262 672618 154346 672854
rect 154582 672618 154614 672854
rect 153994 657000 154614 672618
rect 155394 704838 156014 705830
rect 155394 704602 155426 704838
rect 155662 704602 155746 704838
rect 155982 704602 156014 704838
rect 155394 704518 156014 704602
rect 155394 704282 155426 704518
rect 155662 704282 155746 704518
rect 155982 704282 156014 704518
rect 155394 687454 156014 704282
rect 155394 687218 155426 687454
rect 155662 687218 155746 687454
rect 155982 687218 156014 687454
rect 155394 687134 156014 687218
rect 155394 686898 155426 687134
rect 155662 686898 155746 687134
rect 155982 686898 156014 687134
rect 155394 657000 156014 686898
rect 156314 698614 156934 710042
rect 161434 711558 162054 711590
rect 161434 711322 161466 711558
rect 161702 711322 161786 711558
rect 162022 711322 162054 711558
rect 161434 711238 162054 711322
rect 161434 711002 161466 711238
rect 161702 711002 161786 711238
rect 162022 711002 162054 711238
rect 156314 698378 156346 698614
rect 156582 698378 156666 698614
rect 156902 698378 156934 698614
rect 156314 698294 156934 698378
rect 156314 698058 156346 698294
rect 156582 698058 156666 698294
rect 156902 698058 156934 698294
rect 156314 662614 156934 698058
rect 156314 662378 156346 662614
rect 156582 662378 156666 662614
rect 156902 662378 156934 662614
rect 156314 662294 156934 662378
rect 156314 662058 156346 662294
rect 156582 662058 156666 662294
rect 156902 662058 156934 662294
rect 156314 657000 156934 662058
rect 157714 709638 158334 709670
rect 157714 709402 157746 709638
rect 157982 709402 158066 709638
rect 158302 709402 158334 709638
rect 157714 709318 158334 709402
rect 157714 709082 157746 709318
rect 157982 709082 158066 709318
rect 158302 709082 158334 709318
rect 157714 676894 158334 709082
rect 157714 676658 157746 676894
rect 157982 676658 158066 676894
rect 158302 676658 158334 676894
rect 157714 676574 158334 676658
rect 157714 676338 157746 676574
rect 157982 676338 158066 676574
rect 158302 676338 158334 676574
rect 157714 657000 158334 676338
rect 159114 706758 159734 707750
rect 159114 706522 159146 706758
rect 159382 706522 159466 706758
rect 159702 706522 159734 706758
rect 159114 706438 159734 706522
rect 159114 706202 159146 706438
rect 159382 706202 159466 706438
rect 159702 706202 159734 706438
rect 159114 691174 159734 706202
rect 159114 690938 159146 691174
rect 159382 690938 159466 691174
rect 159702 690938 159734 691174
rect 159114 690854 159734 690938
rect 159114 690618 159146 690854
rect 159382 690618 159466 690854
rect 159702 690618 159734 690854
rect 159114 657000 159734 690618
rect 160514 705798 161134 705830
rect 160514 705562 160546 705798
rect 160782 705562 160866 705798
rect 161102 705562 161134 705798
rect 160514 705478 161134 705562
rect 160514 705242 160546 705478
rect 160782 705242 160866 705478
rect 161102 705242 161134 705478
rect 160514 669454 161134 705242
rect 160514 669218 160546 669454
rect 160782 669218 160866 669454
rect 161102 669218 161134 669454
rect 160514 669134 161134 669218
rect 160514 668898 160546 669134
rect 160782 668898 160866 669134
rect 161102 668898 161134 669134
rect 160514 657000 161134 668898
rect 161434 680614 162054 711002
rect 166554 710598 167174 711590
rect 166554 710362 166586 710598
rect 166822 710362 166906 710598
rect 167142 710362 167174 710598
rect 166554 710278 167174 710362
rect 166554 710042 166586 710278
rect 166822 710042 166906 710278
rect 167142 710042 167174 710278
rect 161434 680378 161466 680614
rect 161702 680378 161786 680614
rect 162022 680378 162054 680614
rect 161434 680294 162054 680378
rect 161434 680058 161466 680294
rect 161702 680058 161786 680294
rect 162022 680058 162054 680294
rect 161434 657000 162054 680058
rect 162834 708678 163454 709670
rect 162834 708442 162866 708678
rect 163102 708442 163186 708678
rect 163422 708442 163454 708678
rect 162834 708358 163454 708442
rect 162834 708122 162866 708358
rect 163102 708122 163186 708358
rect 163422 708122 163454 708358
rect 162834 694894 163454 708122
rect 162834 694658 162866 694894
rect 163102 694658 163186 694894
rect 163422 694658 163454 694894
rect 162834 694574 163454 694658
rect 162834 694338 162866 694574
rect 163102 694338 163186 694574
rect 163422 694338 163454 694574
rect 162834 658894 163454 694338
rect 162834 658658 162866 658894
rect 163102 658658 163186 658894
rect 163422 658658 163454 658894
rect 162834 658574 163454 658658
rect 162834 658338 162866 658574
rect 163102 658338 163186 658574
rect 163422 658338 163454 658574
rect 162834 657000 163454 658338
rect 164234 707718 164854 707750
rect 164234 707482 164266 707718
rect 164502 707482 164586 707718
rect 164822 707482 164854 707718
rect 164234 707398 164854 707482
rect 164234 707162 164266 707398
rect 164502 707162 164586 707398
rect 164822 707162 164854 707398
rect 164234 673174 164854 707162
rect 164234 672938 164266 673174
rect 164502 672938 164586 673174
rect 164822 672938 164854 673174
rect 164234 672854 164854 672938
rect 164234 672618 164266 672854
rect 164502 672618 164586 672854
rect 164822 672618 164854 672854
rect 164234 657000 164854 672618
rect 165634 704838 166254 705830
rect 165634 704602 165666 704838
rect 165902 704602 165986 704838
rect 166222 704602 166254 704838
rect 165634 704518 166254 704602
rect 165634 704282 165666 704518
rect 165902 704282 165986 704518
rect 166222 704282 166254 704518
rect 165634 687454 166254 704282
rect 165634 687218 165666 687454
rect 165902 687218 165986 687454
rect 166222 687218 166254 687454
rect 165634 687134 166254 687218
rect 165634 686898 165666 687134
rect 165902 686898 165986 687134
rect 166222 686898 166254 687134
rect 165634 657000 166254 686898
rect 166554 698614 167174 710042
rect 171674 711558 172294 711590
rect 171674 711322 171706 711558
rect 171942 711322 172026 711558
rect 172262 711322 172294 711558
rect 171674 711238 172294 711322
rect 171674 711002 171706 711238
rect 171942 711002 172026 711238
rect 172262 711002 172294 711238
rect 166554 698378 166586 698614
rect 166822 698378 166906 698614
rect 167142 698378 167174 698614
rect 166554 698294 167174 698378
rect 166554 698058 166586 698294
rect 166822 698058 166906 698294
rect 167142 698058 167174 698294
rect 166554 662614 167174 698058
rect 166554 662378 166586 662614
rect 166822 662378 166906 662614
rect 167142 662378 167174 662614
rect 166554 662294 167174 662378
rect 166554 662058 166586 662294
rect 166822 662058 166906 662294
rect 167142 662058 167174 662294
rect 166554 657000 167174 662058
rect 167954 709638 168574 709670
rect 167954 709402 167986 709638
rect 168222 709402 168306 709638
rect 168542 709402 168574 709638
rect 167954 709318 168574 709402
rect 167954 709082 167986 709318
rect 168222 709082 168306 709318
rect 168542 709082 168574 709318
rect 167954 676894 168574 709082
rect 167954 676658 167986 676894
rect 168222 676658 168306 676894
rect 168542 676658 168574 676894
rect 167954 676574 168574 676658
rect 167954 676338 167986 676574
rect 168222 676338 168306 676574
rect 168542 676338 168574 676574
rect 167954 657000 168574 676338
rect 169354 706758 169974 707750
rect 169354 706522 169386 706758
rect 169622 706522 169706 706758
rect 169942 706522 169974 706758
rect 169354 706438 169974 706522
rect 169354 706202 169386 706438
rect 169622 706202 169706 706438
rect 169942 706202 169974 706438
rect 169354 691174 169974 706202
rect 169354 690938 169386 691174
rect 169622 690938 169706 691174
rect 169942 690938 169974 691174
rect 169354 690854 169974 690938
rect 169354 690618 169386 690854
rect 169622 690618 169706 690854
rect 169942 690618 169974 690854
rect 169354 657000 169974 690618
rect 170754 705798 171374 705830
rect 170754 705562 170786 705798
rect 171022 705562 171106 705798
rect 171342 705562 171374 705798
rect 170754 705478 171374 705562
rect 170754 705242 170786 705478
rect 171022 705242 171106 705478
rect 171342 705242 171374 705478
rect 170754 669454 171374 705242
rect 170754 669218 170786 669454
rect 171022 669218 171106 669454
rect 171342 669218 171374 669454
rect 170754 669134 171374 669218
rect 170754 668898 170786 669134
rect 171022 668898 171106 669134
rect 171342 668898 171374 669134
rect 170754 657000 171374 668898
rect 171674 680614 172294 711002
rect 176794 710598 177414 711590
rect 176794 710362 176826 710598
rect 177062 710362 177146 710598
rect 177382 710362 177414 710598
rect 176794 710278 177414 710362
rect 176794 710042 176826 710278
rect 177062 710042 177146 710278
rect 177382 710042 177414 710278
rect 171674 680378 171706 680614
rect 171942 680378 172026 680614
rect 172262 680378 172294 680614
rect 171674 680294 172294 680378
rect 171674 680058 171706 680294
rect 171942 680058 172026 680294
rect 172262 680058 172294 680294
rect 171674 657000 172294 680058
rect 173074 708678 173694 709670
rect 173074 708442 173106 708678
rect 173342 708442 173426 708678
rect 173662 708442 173694 708678
rect 173074 708358 173694 708442
rect 173074 708122 173106 708358
rect 173342 708122 173426 708358
rect 173662 708122 173694 708358
rect 173074 694894 173694 708122
rect 173074 694658 173106 694894
rect 173342 694658 173426 694894
rect 173662 694658 173694 694894
rect 173074 694574 173694 694658
rect 173074 694338 173106 694574
rect 173342 694338 173426 694574
rect 173662 694338 173694 694574
rect 173074 658894 173694 694338
rect 173074 658658 173106 658894
rect 173342 658658 173426 658894
rect 173662 658658 173694 658894
rect 173074 658574 173694 658658
rect 173074 658338 173106 658574
rect 173342 658338 173426 658574
rect 173662 658338 173694 658574
rect 173074 657000 173694 658338
rect 174474 707718 175094 707750
rect 174474 707482 174506 707718
rect 174742 707482 174826 707718
rect 175062 707482 175094 707718
rect 174474 707398 175094 707482
rect 174474 707162 174506 707398
rect 174742 707162 174826 707398
rect 175062 707162 175094 707398
rect 174474 673174 175094 707162
rect 174474 672938 174506 673174
rect 174742 672938 174826 673174
rect 175062 672938 175094 673174
rect 174474 672854 175094 672938
rect 174474 672618 174506 672854
rect 174742 672618 174826 672854
rect 175062 672618 175094 672854
rect 174474 657000 175094 672618
rect 175874 704838 176494 705830
rect 175874 704602 175906 704838
rect 176142 704602 176226 704838
rect 176462 704602 176494 704838
rect 175874 704518 176494 704602
rect 175874 704282 175906 704518
rect 176142 704282 176226 704518
rect 176462 704282 176494 704518
rect 175874 687454 176494 704282
rect 175874 687218 175906 687454
rect 176142 687218 176226 687454
rect 176462 687218 176494 687454
rect 175874 687134 176494 687218
rect 175874 686898 175906 687134
rect 176142 686898 176226 687134
rect 176462 686898 176494 687134
rect 175874 657000 176494 686898
rect 176794 698614 177414 710042
rect 181914 711558 182534 711590
rect 181914 711322 181946 711558
rect 182182 711322 182266 711558
rect 182502 711322 182534 711558
rect 181914 711238 182534 711322
rect 181914 711002 181946 711238
rect 182182 711002 182266 711238
rect 182502 711002 182534 711238
rect 176794 698378 176826 698614
rect 177062 698378 177146 698614
rect 177382 698378 177414 698614
rect 176794 698294 177414 698378
rect 176794 698058 176826 698294
rect 177062 698058 177146 698294
rect 177382 698058 177414 698294
rect 176794 662614 177414 698058
rect 176794 662378 176826 662614
rect 177062 662378 177146 662614
rect 177382 662378 177414 662614
rect 176794 662294 177414 662378
rect 176794 662058 176826 662294
rect 177062 662058 177146 662294
rect 177382 662058 177414 662294
rect 176794 657000 177414 662058
rect 178194 709638 178814 709670
rect 178194 709402 178226 709638
rect 178462 709402 178546 709638
rect 178782 709402 178814 709638
rect 178194 709318 178814 709402
rect 178194 709082 178226 709318
rect 178462 709082 178546 709318
rect 178782 709082 178814 709318
rect 178194 676894 178814 709082
rect 178194 676658 178226 676894
rect 178462 676658 178546 676894
rect 178782 676658 178814 676894
rect 178194 676574 178814 676658
rect 178194 676338 178226 676574
rect 178462 676338 178546 676574
rect 178782 676338 178814 676574
rect 178194 657000 178814 676338
rect 179594 706758 180214 707750
rect 179594 706522 179626 706758
rect 179862 706522 179946 706758
rect 180182 706522 180214 706758
rect 179594 706438 180214 706522
rect 179594 706202 179626 706438
rect 179862 706202 179946 706438
rect 180182 706202 180214 706438
rect 179594 691174 180214 706202
rect 179594 690938 179626 691174
rect 179862 690938 179946 691174
rect 180182 690938 180214 691174
rect 179594 690854 180214 690938
rect 179594 690618 179626 690854
rect 179862 690618 179946 690854
rect 180182 690618 180214 690854
rect 179594 657000 180214 690618
rect 180994 705798 181614 705830
rect 180994 705562 181026 705798
rect 181262 705562 181346 705798
rect 181582 705562 181614 705798
rect 180994 705478 181614 705562
rect 180994 705242 181026 705478
rect 181262 705242 181346 705478
rect 181582 705242 181614 705478
rect 180994 669454 181614 705242
rect 180994 669218 181026 669454
rect 181262 669218 181346 669454
rect 181582 669218 181614 669454
rect 180994 669134 181614 669218
rect 180994 668898 181026 669134
rect 181262 668898 181346 669134
rect 181582 668898 181614 669134
rect 180994 657000 181614 668898
rect 181914 680614 182534 711002
rect 187034 710598 187654 711590
rect 187034 710362 187066 710598
rect 187302 710362 187386 710598
rect 187622 710362 187654 710598
rect 187034 710278 187654 710362
rect 187034 710042 187066 710278
rect 187302 710042 187386 710278
rect 187622 710042 187654 710278
rect 181914 680378 181946 680614
rect 182182 680378 182266 680614
rect 182502 680378 182534 680614
rect 181914 680294 182534 680378
rect 181914 680058 181946 680294
rect 182182 680058 182266 680294
rect 182502 680058 182534 680294
rect 181914 657000 182534 680058
rect 183314 708678 183934 709670
rect 183314 708442 183346 708678
rect 183582 708442 183666 708678
rect 183902 708442 183934 708678
rect 183314 708358 183934 708442
rect 183314 708122 183346 708358
rect 183582 708122 183666 708358
rect 183902 708122 183934 708358
rect 183314 694894 183934 708122
rect 183314 694658 183346 694894
rect 183582 694658 183666 694894
rect 183902 694658 183934 694894
rect 183314 694574 183934 694658
rect 183314 694338 183346 694574
rect 183582 694338 183666 694574
rect 183902 694338 183934 694574
rect 183314 658894 183934 694338
rect 183314 658658 183346 658894
rect 183582 658658 183666 658894
rect 183902 658658 183934 658894
rect 183314 658574 183934 658658
rect 183314 658338 183346 658574
rect 183582 658338 183666 658574
rect 183902 658338 183934 658574
rect 183314 657000 183934 658338
rect 184714 707718 185334 707750
rect 184714 707482 184746 707718
rect 184982 707482 185066 707718
rect 185302 707482 185334 707718
rect 184714 707398 185334 707482
rect 184714 707162 184746 707398
rect 184982 707162 185066 707398
rect 185302 707162 185334 707398
rect 184714 673174 185334 707162
rect 184714 672938 184746 673174
rect 184982 672938 185066 673174
rect 185302 672938 185334 673174
rect 184714 672854 185334 672938
rect 184714 672618 184746 672854
rect 184982 672618 185066 672854
rect 185302 672618 185334 672854
rect 184714 657000 185334 672618
rect 186114 704838 186734 705830
rect 186114 704602 186146 704838
rect 186382 704602 186466 704838
rect 186702 704602 186734 704838
rect 186114 704518 186734 704602
rect 186114 704282 186146 704518
rect 186382 704282 186466 704518
rect 186702 704282 186734 704518
rect 186114 687454 186734 704282
rect 186114 687218 186146 687454
rect 186382 687218 186466 687454
rect 186702 687218 186734 687454
rect 186114 687134 186734 687218
rect 186114 686898 186146 687134
rect 186382 686898 186466 687134
rect 186702 686898 186734 687134
rect 186114 657000 186734 686898
rect 187034 698614 187654 710042
rect 192154 711558 192774 711590
rect 192154 711322 192186 711558
rect 192422 711322 192506 711558
rect 192742 711322 192774 711558
rect 192154 711238 192774 711322
rect 192154 711002 192186 711238
rect 192422 711002 192506 711238
rect 192742 711002 192774 711238
rect 187034 698378 187066 698614
rect 187302 698378 187386 698614
rect 187622 698378 187654 698614
rect 187034 698294 187654 698378
rect 187034 698058 187066 698294
rect 187302 698058 187386 698294
rect 187622 698058 187654 698294
rect 187034 662614 187654 698058
rect 187034 662378 187066 662614
rect 187302 662378 187386 662614
rect 187622 662378 187654 662614
rect 187034 662294 187654 662378
rect 187034 662058 187066 662294
rect 187302 662058 187386 662294
rect 187622 662058 187654 662294
rect 187034 657000 187654 662058
rect 188434 709638 189054 709670
rect 188434 709402 188466 709638
rect 188702 709402 188786 709638
rect 189022 709402 189054 709638
rect 188434 709318 189054 709402
rect 188434 709082 188466 709318
rect 188702 709082 188786 709318
rect 189022 709082 189054 709318
rect 188434 676894 189054 709082
rect 188434 676658 188466 676894
rect 188702 676658 188786 676894
rect 189022 676658 189054 676894
rect 188434 676574 189054 676658
rect 188434 676338 188466 676574
rect 188702 676338 188786 676574
rect 189022 676338 189054 676574
rect 188434 657000 189054 676338
rect 189834 706758 190454 707750
rect 189834 706522 189866 706758
rect 190102 706522 190186 706758
rect 190422 706522 190454 706758
rect 189834 706438 190454 706522
rect 189834 706202 189866 706438
rect 190102 706202 190186 706438
rect 190422 706202 190454 706438
rect 189834 691174 190454 706202
rect 189834 690938 189866 691174
rect 190102 690938 190186 691174
rect 190422 690938 190454 691174
rect 189834 690854 190454 690938
rect 189834 690618 189866 690854
rect 190102 690618 190186 690854
rect 190422 690618 190454 690854
rect 189834 657000 190454 690618
rect 191234 705798 191854 705830
rect 191234 705562 191266 705798
rect 191502 705562 191586 705798
rect 191822 705562 191854 705798
rect 191234 705478 191854 705562
rect 191234 705242 191266 705478
rect 191502 705242 191586 705478
rect 191822 705242 191854 705478
rect 191234 669454 191854 705242
rect 191234 669218 191266 669454
rect 191502 669218 191586 669454
rect 191822 669218 191854 669454
rect 191234 669134 191854 669218
rect 191234 668898 191266 669134
rect 191502 668898 191586 669134
rect 191822 668898 191854 669134
rect 191234 657000 191854 668898
rect 192154 680614 192774 711002
rect 197274 710598 197894 711590
rect 197274 710362 197306 710598
rect 197542 710362 197626 710598
rect 197862 710362 197894 710598
rect 197274 710278 197894 710362
rect 197274 710042 197306 710278
rect 197542 710042 197626 710278
rect 197862 710042 197894 710278
rect 192154 680378 192186 680614
rect 192422 680378 192506 680614
rect 192742 680378 192774 680614
rect 192154 680294 192774 680378
rect 192154 680058 192186 680294
rect 192422 680058 192506 680294
rect 192742 680058 192774 680294
rect 192154 657000 192774 680058
rect 193554 708678 194174 709670
rect 193554 708442 193586 708678
rect 193822 708442 193906 708678
rect 194142 708442 194174 708678
rect 193554 708358 194174 708442
rect 193554 708122 193586 708358
rect 193822 708122 193906 708358
rect 194142 708122 194174 708358
rect 193554 694894 194174 708122
rect 193554 694658 193586 694894
rect 193822 694658 193906 694894
rect 194142 694658 194174 694894
rect 193554 694574 194174 694658
rect 193554 694338 193586 694574
rect 193822 694338 193906 694574
rect 194142 694338 194174 694574
rect 193554 658894 194174 694338
rect 193554 658658 193586 658894
rect 193822 658658 193906 658894
rect 194142 658658 194174 658894
rect 193554 658574 194174 658658
rect 193554 658338 193586 658574
rect 193822 658338 193906 658574
rect 194142 658338 194174 658574
rect 193554 657000 194174 658338
rect 194954 707718 195574 707750
rect 194954 707482 194986 707718
rect 195222 707482 195306 707718
rect 195542 707482 195574 707718
rect 194954 707398 195574 707482
rect 194954 707162 194986 707398
rect 195222 707162 195306 707398
rect 195542 707162 195574 707398
rect 194954 673174 195574 707162
rect 194954 672938 194986 673174
rect 195222 672938 195306 673174
rect 195542 672938 195574 673174
rect 194954 672854 195574 672938
rect 194954 672618 194986 672854
rect 195222 672618 195306 672854
rect 195542 672618 195574 672854
rect 194954 657000 195574 672618
rect 196354 704838 196974 705830
rect 196354 704602 196386 704838
rect 196622 704602 196706 704838
rect 196942 704602 196974 704838
rect 196354 704518 196974 704602
rect 196354 704282 196386 704518
rect 196622 704282 196706 704518
rect 196942 704282 196974 704518
rect 196354 687454 196974 704282
rect 196354 687218 196386 687454
rect 196622 687218 196706 687454
rect 196942 687218 196974 687454
rect 196354 687134 196974 687218
rect 196354 686898 196386 687134
rect 196622 686898 196706 687134
rect 196942 686898 196974 687134
rect 196354 657000 196974 686898
rect 197274 698614 197894 710042
rect 202394 711558 203014 711590
rect 202394 711322 202426 711558
rect 202662 711322 202746 711558
rect 202982 711322 203014 711558
rect 202394 711238 203014 711322
rect 202394 711002 202426 711238
rect 202662 711002 202746 711238
rect 202982 711002 203014 711238
rect 197274 698378 197306 698614
rect 197542 698378 197626 698614
rect 197862 698378 197894 698614
rect 197274 698294 197894 698378
rect 197274 698058 197306 698294
rect 197542 698058 197626 698294
rect 197862 698058 197894 698294
rect 197274 662614 197894 698058
rect 197274 662378 197306 662614
rect 197542 662378 197626 662614
rect 197862 662378 197894 662614
rect 197274 662294 197894 662378
rect 197274 662058 197306 662294
rect 197542 662058 197626 662294
rect 197862 662058 197894 662294
rect 197274 657000 197894 662058
rect 198674 709638 199294 709670
rect 198674 709402 198706 709638
rect 198942 709402 199026 709638
rect 199262 709402 199294 709638
rect 198674 709318 199294 709402
rect 198674 709082 198706 709318
rect 198942 709082 199026 709318
rect 199262 709082 199294 709318
rect 198674 676894 199294 709082
rect 198674 676658 198706 676894
rect 198942 676658 199026 676894
rect 199262 676658 199294 676894
rect 198674 676574 199294 676658
rect 198674 676338 198706 676574
rect 198942 676338 199026 676574
rect 199262 676338 199294 676574
rect 198674 657000 199294 676338
rect 200074 706758 200694 707750
rect 200074 706522 200106 706758
rect 200342 706522 200426 706758
rect 200662 706522 200694 706758
rect 200074 706438 200694 706522
rect 200074 706202 200106 706438
rect 200342 706202 200426 706438
rect 200662 706202 200694 706438
rect 200074 691174 200694 706202
rect 200074 690938 200106 691174
rect 200342 690938 200426 691174
rect 200662 690938 200694 691174
rect 200074 690854 200694 690938
rect 200074 690618 200106 690854
rect 200342 690618 200426 690854
rect 200662 690618 200694 690854
rect 200074 657000 200694 690618
rect 201474 705798 202094 705830
rect 201474 705562 201506 705798
rect 201742 705562 201826 705798
rect 202062 705562 202094 705798
rect 201474 705478 202094 705562
rect 201474 705242 201506 705478
rect 201742 705242 201826 705478
rect 202062 705242 202094 705478
rect 201474 669454 202094 705242
rect 201474 669218 201506 669454
rect 201742 669218 201826 669454
rect 202062 669218 202094 669454
rect 201474 669134 202094 669218
rect 201474 668898 201506 669134
rect 201742 668898 201826 669134
rect 202062 668898 202094 669134
rect 201474 657000 202094 668898
rect 202394 680614 203014 711002
rect 207514 710598 208134 711590
rect 207514 710362 207546 710598
rect 207782 710362 207866 710598
rect 208102 710362 208134 710598
rect 207514 710278 208134 710362
rect 207514 710042 207546 710278
rect 207782 710042 207866 710278
rect 208102 710042 208134 710278
rect 202394 680378 202426 680614
rect 202662 680378 202746 680614
rect 202982 680378 203014 680614
rect 202394 680294 203014 680378
rect 202394 680058 202426 680294
rect 202662 680058 202746 680294
rect 202982 680058 203014 680294
rect 202394 657000 203014 680058
rect 203794 708678 204414 709670
rect 203794 708442 203826 708678
rect 204062 708442 204146 708678
rect 204382 708442 204414 708678
rect 203794 708358 204414 708442
rect 203794 708122 203826 708358
rect 204062 708122 204146 708358
rect 204382 708122 204414 708358
rect 203794 694894 204414 708122
rect 203794 694658 203826 694894
rect 204062 694658 204146 694894
rect 204382 694658 204414 694894
rect 203794 694574 204414 694658
rect 203794 694338 203826 694574
rect 204062 694338 204146 694574
rect 204382 694338 204414 694574
rect 203794 658894 204414 694338
rect 203794 658658 203826 658894
rect 204062 658658 204146 658894
rect 204382 658658 204414 658894
rect 203794 658574 204414 658658
rect 203794 658338 203826 658574
rect 204062 658338 204146 658574
rect 204382 658338 204414 658574
rect 203794 657000 204414 658338
rect 205194 707718 205814 707750
rect 205194 707482 205226 707718
rect 205462 707482 205546 707718
rect 205782 707482 205814 707718
rect 205194 707398 205814 707482
rect 205194 707162 205226 707398
rect 205462 707162 205546 707398
rect 205782 707162 205814 707398
rect 205194 673174 205814 707162
rect 205194 672938 205226 673174
rect 205462 672938 205546 673174
rect 205782 672938 205814 673174
rect 205194 672854 205814 672938
rect 205194 672618 205226 672854
rect 205462 672618 205546 672854
rect 205782 672618 205814 672854
rect 205194 657000 205814 672618
rect 206594 704838 207214 705830
rect 206594 704602 206626 704838
rect 206862 704602 206946 704838
rect 207182 704602 207214 704838
rect 206594 704518 207214 704602
rect 206594 704282 206626 704518
rect 206862 704282 206946 704518
rect 207182 704282 207214 704518
rect 206594 687454 207214 704282
rect 206594 687218 206626 687454
rect 206862 687218 206946 687454
rect 207182 687218 207214 687454
rect 206594 687134 207214 687218
rect 206594 686898 206626 687134
rect 206862 686898 206946 687134
rect 207182 686898 207214 687134
rect 206594 657000 207214 686898
rect 207514 698614 208134 710042
rect 212634 711558 213254 711590
rect 212634 711322 212666 711558
rect 212902 711322 212986 711558
rect 213222 711322 213254 711558
rect 212634 711238 213254 711322
rect 212634 711002 212666 711238
rect 212902 711002 212986 711238
rect 213222 711002 213254 711238
rect 207514 698378 207546 698614
rect 207782 698378 207866 698614
rect 208102 698378 208134 698614
rect 207514 698294 208134 698378
rect 207514 698058 207546 698294
rect 207782 698058 207866 698294
rect 208102 698058 208134 698294
rect 207514 662614 208134 698058
rect 207514 662378 207546 662614
rect 207782 662378 207866 662614
rect 208102 662378 208134 662614
rect 207514 662294 208134 662378
rect 207514 662058 207546 662294
rect 207782 662058 207866 662294
rect 208102 662058 208134 662294
rect 207514 657000 208134 662058
rect 208914 709638 209534 709670
rect 208914 709402 208946 709638
rect 209182 709402 209266 709638
rect 209502 709402 209534 709638
rect 208914 709318 209534 709402
rect 208914 709082 208946 709318
rect 209182 709082 209266 709318
rect 209502 709082 209534 709318
rect 208914 676894 209534 709082
rect 208914 676658 208946 676894
rect 209182 676658 209266 676894
rect 209502 676658 209534 676894
rect 208914 676574 209534 676658
rect 208914 676338 208946 676574
rect 209182 676338 209266 676574
rect 209502 676338 209534 676574
rect 208914 657000 209534 676338
rect 210314 706758 210934 707750
rect 210314 706522 210346 706758
rect 210582 706522 210666 706758
rect 210902 706522 210934 706758
rect 210314 706438 210934 706522
rect 210314 706202 210346 706438
rect 210582 706202 210666 706438
rect 210902 706202 210934 706438
rect 210314 691174 210934 706202
rect 210314 690938 210346 691174
rect 210582 690938 210666 691174
rect 210902 690938 210934 691174
rect 210314 690854 210934 690938
rect 210314 690618 210346 690854
rect 210582 690618 210666 690854
rect 210902 690618 210934 690854
rect 210314 657000 210934 690618
rect 211714 705798 212334 705830
rect 211714 705562 211746 705798
rect 211982 705562 212066 705798
rect 212302 705562 212334 705798
rect 211714 705478 212334 705562
rect 211714 705242 211746 705478
rect 211982 705242 212066 705478
rect 212302 705242 212334 705478
rect 211714 669454 212334 705242
rect 211714 669218 211746 669454
rect 211982 669218 212066 669454
rect 212302 669218 212334 669454
rect 211714 669134 212334 669218
rect 211714 668898 211746 669134
rect 211982 668898 212066 669134
rect 212302 668898 212334 669134
rect 211714 657000 212334 668898
rect 212634 680614 213254 711002
rect 217754 710598 218374 711590
rect 217754 710362 217786 710598
rect 218022 710362 218106 710598
rect 218342 710362 218374 710598
rect 217754 710278 218374 710362
rect 217754 710042 217786 710278
rect 218022 710042 218106 710278
rect 218342 710042 218374 710278
rect 212634 680378 212666 680614
rect 212902 680378 212986 680614
rect 213222 680378 213254 680614
rect 212634 680294 213254 680378
rect 212634 680058 212666 680294
rect 212902 680058 212986 680294
rect 213222 680058 213254 680294
rect 212634 657000 213254 680058
rect 214034 708678 214654 709670
rect 214034 708442 214066 708678
rect 214302 708442 214386 708678
rect 214622 708442 214654 708678
rect 214034 708358 214654 708442
rect 214034 708122 214066 708358
rect 214302 708122 214386 708358
rect 214622 708122 214654 708358
rect 214034 694894 214654 708122
rect 214034 694658 214066 694894
rect 214302 694658 214386 694894
rect 214622 694658 214654 694894
rect 214034 694574 214654 694658
rect 214034 694338 214066 694574
rect 214302 694338 214386 694574
rect 214622 694338 214654 694574
rect 214034 658894 214654 694338
rect 214034 658658 214066 658894
rect 214302 658658 214386 658894
rect 214622 658658 214654 658894
rect 214034 658574 214654 658658
rect 214034 658338 214066 658574
rect 214302 658338 214386 658574
rect 214622 658338 214654 658574
rect 214034 657000 214654 658338
rect 215434 707718 216054 707750
rect 215434 707482 215466 707718
rect 215702 707482 215786 707718
rect 216022 707482 216054 707718
rect 215434 707398 216054 707482
rect 215434 707162 215466 707398
rect 215702 707162 215786 707398
rect 216022 707162 216054 707398
rect 215434 673174 216054 707162
rect 215434 672938 215466 673174
rect 215702 672938 215786 673174
rect 216022 672938 216054 673174
rect 215434 672854 216054 672938
rect 215434 672618 215466 672854
rect 215702 672618 215786 672854
rect 216022 672618 216054 672854
rect 215434 657000 216054 672618
rect 216834 704838 217454 705830
rect 216834 704602 216866 704838
rect 217102 704602 217186 704838
rect 217422 704602 217454 704838
rect 216834 704518 217454 704602
rect 216834 704282 216866 704518
rect 217102 704282 217186 704518
rect 217422 704282 217454 704518
rect 216834 687454 217454 704282
rect 216834 687218 216866 687454
rect 217102 687218 217186 687454
rect 217422 687218 217454 687454
rect 216834 687134 217454 687218
rect 216834 686898 216866 687134
rect 217102 686898 217186 687134
rect 217422 686898 217454 687134
rect 216834 657000 217454 686898
rect 217754 698614 218374 710042
rect 222874 711558 223494 711590
rect 222874 711322 222906 711558
rect 223142 711322 223226 711558
rect 223462 711322 223494 711558
rect 222874 711238 223494 711322
rect 222874 711002 222906 711238
rect 223142 711002 223226 711238
rect 223462 711002 223494 711238
rect 217754 698378 217786 698614
rect 218022 698378 218106 698614
rect 218342 698378 218374 698614
rect 217754 698294 218374 698378
rect 217754 698058 217786 698294
rect 218022 698058 218106 698294
rect 218342 698058 218374 698294
rect 217754 662614 218374 698058
rect 217754 662378 217786 662614
rect 218022 662378 218106 662614
rect 218342 662378 218374 662614
rect 217754 662294 218374 662378
rect 217754 662058 217786 662294
rect 218022 662058 218106 662294
rect 218342 662058 218374 662294
rect 217754 657000 218374 662058
rect 219154 709638 219774 709670
rect 219154 709402 219186 709638
rect 219422 709402 219506 709638
rect 219742 709402 219774 709638
rect 219154 709318 219774 709402
rect 219154 709082 219186 709318
rect 219422 709082 219506 709318
rect 219742 709082 219774 709318
rect 219154 676894 219774 709082
rect 219154 676658 219186 676894
rect 219422 676658 219506 676894
rect 219742 676658 219774 676894
rect 219154 676574 219774 676658
rect 219154 676338 219186 676574
rect 219422 676338 219506 676574
rect 219742 676338 219774 676574
rect 219154 657000 219774 676338
rect 220554 706758 221174 707750
rect 220554 706522 220586 706758
rect 220822 706522 220906 706758
rect 221142 706522 221174 706758
rect 220554 706438 221174 706522
rect 220554 706202 220586 706438
rect 220822 706202 220906 706438
rect 221142 706202 221174 706438
rect 220554 691174 221174 706202
rect 220554 690938 220586 691174
rect 220822 690938 220906 691174
rect 221142 690938 221174 691174
rect 220554 690854 221174 690938
rect 220554 690618 220586 690854
rect 220822 690618 220906 690854
rect 221142 690618 221174 690854
rect 220554 657000 221174 690618
rect 221954 705798 222574 705830
rect 221954 705562 221986 705798
rect 222222 705562 222306 705798
rect 222542 705562 222574 705798
rect 221954 705478 222574 705562
rect 221954 705242 221986 705478
rect 222222 705242 222306 705478
rect 222542 705242 222574 705478
rect 221954 669454 222574 705242
rect 221954 669218 221986 669454
rect 222222 669218 222306 669454
rect 222542 669218 222574 669454
rect 221954 669134 222574 669218
rect 221954 668898 221986 669134
rect 222222 668898 222306 669134
rect 222542 668898 222574 669134
rect 221954 657000 222574 668898
rect 222874 680614 223494 711002
rect 227994 710598 228614 711590
rect 227994 710362 228026 710598
rect 228262 710362 228346 710598
rect 228582 710362 228614 710598
rect 227994 710278 228614 710362
rect 227994 710042 228026 710278
rect 228262 710042 228346 710278
rect 228582 710042 228614 710278
rect 222874 680378 222906 680614
rect 223142 680378 223226 680614
rect 223462 680378 223494 680614
rect 222874 680294 223494 680378
rect 222874 680058 222906 680294
rect 223142 680058 223226 680294
rect 223462 680058 223494 680294
rect 222874 657000 223494 680058
rect 224274 708678 224894 709670
rect 224274 708442 224306 708678
rect 224542 708442 224626 708678
rect 224862 708442 224894 708678
rect 224274 708358 224894 708442
rect 224274 708122 224306 708358
rect 224542 708122 224626 708358
rect 224862 708122 224894 708358
rect 224274 694894 224894 708122
rect 224274 694658 224306 694894
rect 224542 694658 224626 694894
rect 224862 694658 224894 694894
rect 224274 694574 224894 694658
rect 224274 694338 224306 694574
rect 224542 694338 224626 694574
rect 224862 694338 224894 694574
rect 224274 658894 224894 694338
rect 224274 658658 224306 658894
rect 224542 658658 224626 658894
rect 224862 658658 224894 658894
rect 224274 658574 224894 658658
rect 224274 658338 224306 658574
rect 224542 658338 224626 658574
rect 224862 658338 224894 658574
rect 224274 657000 224894 658338
rect 225674 707718 226294 707750
rect 225674 707482 225706 707718
rect 225942 707482 226026 707718
rect 226262 707482 226294 707718
rect 225674 707398 226294 707482
rect 225674 707162 225706 707398
rect 225942 707162 226026 707398
rect 226262 707162 226294 707398
rect 225674 673174 226294 707162
rect 225674 672938 225706 673174
rect 225942 672938 226026 673174
rect 226262 672938 226294 673174
rect 225674 672854 226294 672938
rect 225674 672618 225706 672854
rect 225942 672618 226026 672854
rect 226262 672618 226294 672854
rect 225674 657000 226294 672618
rect 227074 704838 227694 705830
rect 227074 704602 227106 704838
rect 227342 704602 227426 704838
rect 227662 704602 227694 704838
rect 227074 704518 227694 704602
rect 227074 704282 227106 704518
rect 227342 704282 227426 704518
rect 227662 704282 227694 704518
rect 227074 687454 227694 704282
rect 227074 687218 227106 687454
rect 227342 687218 227426 687454
rect 227662 687218 227694 687454
rect 227074 687134 227694 687218
rect 227074 686898 227106 687134
rect 227342 686898 227426 687134
rect 227662 686898 227694 687134
rect 227074 657000 227694 686898
rect 227994 698614 228614 710042
rect 233114 711558 233734 711590
rect 233114 711322 233146 711558
rect 233382 711322 233466 711558
rect 233702 711322 233734 711558
rect 233114 711238 233734 711322
rect 233114 711002 233146 711238
rect 233382 711002 233466 711238
rect 233702 711002 233734 711238
rect 227994 698378 228026 698614
rect 228262 698378 228346 698614
rect 228582 698378 228614 698614
rect 227994 698294 228614 698378
rect 227994 698058 228026 698294
rect 228262 698058 228346 698294
rect 228582 698058 228614 698294
rect 227994 662614 228614 698058
rect 227994 662378 228026 662614
rect 228262 662378 228346 662614
rect 228582 662378 228614 662614
rect 227994 662294 228614 662378
rect 227994 662058 228026 662294
rect 228262 662058 228346 662294
rect 228582 662058 228614 662294
rect 227994 657000 228614 662058
rect 229394 709638 230014 709670
rect 229394 709402 229426 709638
rect 229662 709402 229746 709638
rect 229982 709402 230014 709638
rect 229394 709318 230014 709402
rect 229394 709082 229426 709318
rect 229662 709082 229746 709318
rect 229982 709082 230014 709318
rect 229394 676894 230014 709082
rect 229394 676658 229426 676894
rect 229662 676658 229746 676894
rect 229982 676658 230014 676894
rect 229394 676574 230014 676658
rect 229394 676338 229426 676574
rect 229662 676338 229746 676574
rect 229982 676338 230014 676574
rect 229394 657000 230014 676338
rect 230794 706758 231414 707750
rect 230794 706522 230826 706758
rect 231062 706522 231146 706758
rect 231382 706522 231414 706758
rect 230794 706438 231414 706522
rect 230794 706202 230826 706438
rect 231062 706202 231146 706438
rect 231382 706202 231414 706438
rect 230794 691174 231414 706202
rect 230794 690938 230826 691174
rect 231062 690938 231146 691174
rect 231382 690938 231414 691174
rect 230794 690854 231414 690938
rect 230794 690618 230826 690854
rect 231062 690618 231146 690854
rect 231382 690618 231414 690854
rect 230794 657000 231414 690618
rect 232194 705798 232814 705830
rect 232194 705562 232226 705798
rect 232462 705562 232546 705798
rect 232782 705562 232814 705798
rect 232194 705478 232814 705562
rect 232194 705242 232226 705478
rect 232462 705242 232546 705478
rect 232782 705242 232814 705478
rect 232194 669454 232814 705242
rect 232194 669218 232226 669454
rect 232462 669218 232546 669454
rect 232782 669218 232814 669454
rect 232194 669134 232814 669218
rect 232194 668898 232226 669134
rect 232462 668898 232546 669134
rect 232782 668898 232814 669134
rect 232194 657000 232814 668898
rect 233114 680614 233734 711002
rect 238234 710598 238854 711590
rect 238234 710362 238266 710598
rect 238502 710362 238586 710598
rect 238822 710362 238854 710598
rect 238234 710278 238854 710362
rect 238234 710042 238266 710278
rect 238502 710042 238586 710278
rect 238822 710042 238854 710278
rect 233114 680378 233146 680614
rect 233382 680378 233466 680614
rect 233702 680378 233734 680614
rect 233114 680294 233734 680378
rect 233114 680058 233146 680294
rect 233382 680058 233466 680294
rect 233702 680058 233734 680294
rect 233114 657000 233734 680058
rect 234514 708678 235134 709670
rect 234514 708442 234546 708678
rect 234782 708442 234866 708678
rect 235102 708442 235134 708678
rect 234514 708358 235134 708442
rect 234514 708122 234546 708358
rect 234782 708122 234866 708358
rect 235102 708122 235134 708358
rect 234514 694894 235134 708122
rect 234514 694658 234546 694894
rect 234782 694658 234866 694894
rect 235102 694658 235134 694894
rect 234514 694574 235134 694658
rect 234514 694338 234546 694574
rect 234782 694338 234866 694574
rect 235102 694338 235134 694574
rect 234514 658894 235134 694338
rect 234514 658658 234546 658894
rect 234782 658658 234866 658894
rect 235102 658658 235134 658894
rect 234514 658574 235134 658658
rect 234514 658338 234546 658574
rect 234782 658338 234866 658574
rect 235102 658338 235134 658574
rect 234514 657000 235134 658338
rect 235914 707718 236534 707750
rect 235914 707482 235946 707718
rect 236182 707482 236266 707718
rect 236502 707482 236534 707718
rect 235914 707398 236534 707482
rect 235914 707162 235946 707398
rect 236182 707162 236266 707398
rect 236502 707162 236534 707398
rect 235914 673174 236534 707162
rect 235914 672938 235946 673174
rect 236182 672938 236266 673174
rect 236502 672938 236534 673174
rect 235914 672854 236534 672938
rect 235914 672618 235946 672854
rect 236182 672618 236266 672854
rect 236502 672618 236534 672854
rect 235914 657000 236534 672618
rect 237314 704838 237934 705830
rect 237314 704602 237346 704838
rect 237582 704602 237666 704838
rect 237902 704602 237934 704838
rect 237314 704518 237934 704602
rect 237314 704282 237346 704518
rect 237582 704282 237666 704518
rect 237902 704282 237934 704518
rect 237314 687454 237934 704282
rect 237314 687218 237346 687454
rect 237582 687218 237666 687454
rect 237902 687218 237934 687454
rect 237314 687134 237934 687218
rect 237314 686898 237346 687134
rect 237582 686898 237666 687134
rect 237902 686898 237934 687134
rect 237314 657000 237934 686898
rect 238234 698614 238854 710042
rect 243354 711558 243974 711590
rect 243354 711322 243386 711558
rect 243622 711322 243706 711558
rect 243942 711322 243974 711558
rect 243354 711238 243974 711322
rect 243354 711002 243386 711238
rect 243622 711002 243706 711238
rect 243942 711002 243974 711238
rect 238234 698378 238266 698614
rect 238502 698378 238586 698614
rect 238822 698378 238854 698614
rect 238234 698294 238854 698378
rect 238234 698058 238266 698294
rect 238502 698058 238586 698294
rect 238822 698058 238854 698294
rect 238234 662614 238854 698058
rect 238234 662378 238266 662614
rect 238502 662378 238586 662614
rect 238822 662378 238854 662614
rect 238234 662294 238854 662378
rect 238234 662058 238266 662294
rect 238502 662058 238586 662294
rect 238822 662058 238854 662294
rect 238234 657000 238854 662058
rect 239634 709638 240254 709670
rect 239634 709402 239666 709638
rect 239902 709402 239986 709638
rect 240222 709402 240254 709638
rect 239634 709318 240254 709402
rect 239634 709082 239666 709318
rect 239902 709082 239986 709318
rect 240222 709082 240254 709318
rect 239634 676894 240254 709082
rect 239634 676658 239666 676894
rect 239902 676658 239986 676894
rect 240222 676658 240254 676894
rect 239634 676574 240254 676658
rect 239634 676338 239666 676574
rect 239902 676338 239986 676574
rect 240222 676338 240254 676574
rect 239634 657000 240254 676338
rect 241034 706758 241654 707750
rect 241034 706522 241066 706758
rect 241302 706522 241386 706758
rect 241622 706522 241654 706758
rect 241034 706438 241654 706522
rect 241034 706202 241066 706438
rect 241302 706202 241386 706438
rect 241622 706202 241654 706438
rect 241034 691174 241654 706202
rect 241034 690938 241066 691174
rect 241302 690938 241386 691174
rect 241622 690938 241654 691174
rect 241034 690854 241654 690938
rect 241034 690618 241066 690854
rect 241302 690618 241386 690854
rect 241622 690618 241654 690854
rect 241034 657000 241654 690618
rect 242434 705798 243054 705830
rect 242434 705562 242466 705798
rect 242702 705562 242786 705798
rect 243022 705562 243054 705798
rect 242434 705478 243054 705562
rect 242434 705242 242466 705478
rect 242702 705242 242786 705478
rect 243022 705242 243054 705478
rect 242434 669454 243054 705242
rect 242434 669218 242466 669454
rect 242702 669218 242786 669454
rect 243022 669218 243054 669454
rect 242434 669134 243054 669218
rect 242434 668898 242466 669134
rect 242702 668898 242786 669134
rect 243022 668898 243054 669134
rect 242434 657000 243054 668898
rect 243354 680614 243974 711002
rect 248474 710598 249094 711590
rect 248474 710362 248506 710598
rect 248742 710362 248826 710598
rect 249062 710362 249094 710598
rect 248474 710278 249094 710362
rect 248474 710042 248506 710278
rect 248742 710042 248826 710278
rect 249062 710042 249094 710278
rect 243354 680378 243386 680614
rect 243622 680378 243706 680614
rect 243942 680378 243974 680614
rect 243354 680294 243974 680378
rect 243354 680058 243386 680294
rect 243622 680058 243706 680294
rect 243942 680058 243974 680294
rect 243354 657000 243974 680058
rect 244754 708678 245374 709670
rect 244754 708442 244786 708678
rect 245022 708442 245106 708678
rect 245342 708442 245374 708678
rect 244754 708358 245374 708442
rect 244754 708122 244786 708358
rect 245022 708122 245106 708358
rect 245342 708122 245374 708358
rect 244754 694894 245374 708122
rect 244754 694658 244786 694894
rect 245022 694658 245106 694894
rect 245342 694658 245374 694894
rect 244754 694574 245374 694658
rect 244754 694338 244786 694574
rect 245022 694338 245106 694574
rect 245342 694338 245374 694574
rect 244754 658894 245374 694338
rect 244754 658658 244786 658894
rect 245022 658658 245106 658894
rect 245342 658658 245374 658894
rect 244754 658574 245374 658658
rect 244754 658338 244786 658574
rect 245022 658338 245106 658574
rect 245342 658338 245374 658574
rect 244754 657000 245374 658338
rect 246154 707718 246774 707750
rect 246154 707482 246186 707718
rect 246422 707482 246506 707718
rect 246742 707482 246774 707718
rect 246154 707398 246774 707482
rect 246154 707162 246186 707398
rect 246422 707162 246506 707398
rect 246742 707162 246774 707398
rect 246154 673174 246774 707162
rect 246154 672938 246186 673174
rect 246422 672938 246506 673174
rect 246742 672938 246774 673174
rect 246154 672854 246774 672938
rect 246154 672618 246186 672854
rect 246422 672618 246506 672854
rect 246742 672618 246774 672854
rect 246154 657000 246774 672618
rect 247554 704838 248174 705830
rect 247554 704602 247586 704838
rect 247822 704602 247906 704838
rect 248142 704602 248174 704838
rect 247554 704518 248174 704602
rect 247554 704282 247586 704518
rect 247822 704282 247906 704518
rect 248142 704282 248174 704518
rect 247554 687454 248174 704282
rect 247554 687218 247586 687454
rect 247822 687218 247906 687454
rect 248142 687218 248174 687454
rect 247554 687134 248174 687218
rect 247554 686898 247586 687134
rect 247822 686898 247906 687134
rect 248142 686898 248174 687134
rect 247554 657000 248174 686898
rect 248474 698614 249094 710042
rect 253594 711558 254214 711590
rect 253594 711322 253626 711558
rect 253862 711322 253946 711558
rect 254182 711322 254214 711558
rect 253594 711238 254214 711322
rect 253594 711002 253626 711238
rect 253862 711002 253946 711238
rect 254182 711002 254214 711238
rect 248474 698378 248506 698614
rect 248742 698378 248826 698614
rect 249062 698378 249094 698614
rect 248474 698294 249094 698378
rect 248474 698058 248506 698294
rect 248742 698058 248826 698294
rect 249062 698058 249094 698294
rect 248474 662614 249094 698058
rect 248474 662378 248506 662614
rect 248742 662378 248826 662614
rect 249062 662378 249094 662614
rect 248474 662294 249094 662378
rect 248474 662058 248506 662294
rect 248742 662058 248826 662294
rect 249062 662058 249094 662294
rect 248474 657000 249094 662058
rect 249874 709638 250494 709670
rect 249874 709402 249906 709638
rect 250142 709402 250226 709638
rect 250462 709402 250494 709638
rect 249874 709318 250494 709402
rect 249874 709082 249906 709318
rect 250142 709082 250226 709318
rect 250462 709082 250494 709318
rect 249874 676894 250494 709082
rect 249874 676658 249906 676894
rect 250142 676658 250226 676894
rect 250462 676658 250494 676894
rect 249874 676574 250494 676658
rect 249874 676338 249906 676574
rect 250142 676338 250226 676574
rect 250462 676338 250494 676574
rect 249874 657000 250494 676338
rect 251274 706758 251894 707750
rect 251274 706522 251306 706758
rect 251542 706522 251626 706758
rect 251862 706522 251894 706758
rect 251274 706438 251894 706522
rect 251274 706202 251306 706438
rect 251542 706202 251626 706438
rect 251862 706202 251894 706438
rect 251274 691174 251894 706202
rect 251274 690938 251306 691174
rect 251542 690938 251626 691174
rect 251862 690938 251894 691174
rect 251274 690854 251894 690938
rect 251274 690618 251306 690854
rect 251542 690618 251626 690854
rect 251862 690618 251894 690854
rect 251274 657000 251894 690618
rect 252674 705798 253294 705830
rect 252674 705562 252706 705798
rect 252942 705562 253026 705798
rect 253262 705562 253294 705798
rect 252674 705478 253294 705562
rect 252674 705242 252706 705478
rect 252942 705242 253026 705478
rect 253262 705242 253294 705478
rect 252674 669454 253294 705242
rect 252674 669218 252706 669454
rect 252942 669218 253026 669454
rect 253262 669218 253294 669454
rect 252674 669134 253294 669218
rect 252674 668898 252706 669134
rect 252942 668898 253026 669134
rect 253262 668898 253294 669134
rect 252674 657000 253294 668898
rect 253594 680614 254214 711002
rect 258714 710598 259334 711590
rect 258714 710362 258746 710598
rect 258982 710362 259066 710598
rect 259302 710362 259334 710598
rect 258714 710278 259334 710362
rect 258714 710042 258746 710278
rect 258982 710042 259066 710278
rect 259302 710042 259334 710278
rect 253594 680378 253626 680614
rect 253862 680378 253946 680614
rect 254182 680378 254214 680614
rect 253594 680294 254214 680378
rect 253594 680058 253626 680294
rect 253862 680058 253946 680294
rect 254182 680058 254214 680294
rect 253594 657000 254214 680058
rect 254994 708678 255614 709670
rect 254994 708442 255026 708678
rect 255262 708442 255346 708678
rect 255582 708442 255614 708678
rect 254994 708358 255614 708442
rect 254994 708122 255026 708358
rect 255262 708122 255346 708358
rect 255582 708122 255614 708358
rect 254994 694894 255614 708122
rect 254994 694658 255026 694894
rect 255262 694658 255346 694894
rect 255582 694658 255614 694894
rect 254994 694574 255614 694658
rect 254994 694338 255026 694574
rect 255262 694338 255346 694574
rect 255582 694338 255614 694574
rect 254994 658894 255614 694338
rect 254994 658658 255026 658894
rect 255262 658658 255346 658894
rect 255582 658658 255614 658894
rect 254994 658574 255614 658658
rect 254994 658338 255026 658574
rect 255262 658338 255346 658574
rect 255582 658338 255614 658574
rect 254994 657000 255614 658338
rect 256394 707718 257014 707750
rect 256394 707482 256426 707718
rect 256662 707482 256746 707718
rect 256982 707482 257014 707718
rect 256394 707398 257014 707482
rect 256394 707162 256426 707398
rect 256662 707162 256746 707398
rect 256982 707162 257014 707398
rect 256394 673174 257014 707162
rect 256394 672938 256426 673174
rect 256662 672938 256746 673174
rect 256982 672938 257014 673174
rect 256394 672854 257014 672938
rect 256394 672618 256426 672854
rect 256662 672618 256746 672854
rect 256982 672618 257014 672854
rect 256394 657000 257014 672618
rect 257794 704838 258414 705830
rect 257794 704602 257826 704838
rect 258062 704602 258146 704838
rect 258382 704602 258414 704838
rect 257794 704518 258414 704602
rect 257794 704282 257826 704518
rect 258062 704282 258146 704518
rect 258382 704282 258414 704518
rect 257794 687454 258414 704282
rect 257794 687218 257826 687454
rect 258062 687218 258146 687454
rect 258382 687218 258414 687454
rect 257794 687134 258414 687218
rect 257794 686898 257826 687134
rect 258062 686898 258146 687134
rect 258382 686898 258414 687134
rect 257794 657000 258414 686898
rect 258714 698614 259334 710042
rect 263834 711558 264454 711590
rect 263834 711322 263866 711558
rect 264102 711322 264186 711558
rect 264422 711322 264454 711558
rect 263834 711238 264454 711322
rect 263834 711002 263866 711238
rect 264102 711002 264186 711238
rect 264422 711002 264454 711238
rect 258714 698378 258746 698614
rect 258982 698378 259066 698614
rect 259302 698378 259334 698614
rect 258714 698294 259334 698378
rect 258714 698058 258746 698294
rect 258982 698058 259066 698294
rect 259302 698058 259334 698294
rect 258714 662614 259334 698058
rect 258714 662378 258746 662614
rect 258982 662378 259066 662614
rect 259302 662378 259334 662614
rect 258714 662294 259334 662378
rect 258714 662058 258746 662294
rect 258982 662058 259066 662294
rect 259302 662058 259334 662294
rect 258714 657000 259334 662058
rect 260114 709638 260734 709670
rect 260114 709402 260146 709638
rect 260382 709402 260466 709638
rect 260702 709402 260734 709638
rect 260114 709318 260734 709402
rect 260114 709082 260146 709318
rect 260382 709082 260466 709318
rect 260702 709082 260734 709318
rect 260114 676894 260734 709082
rect 260114 676658 260146 676894
rect 260382 676658 260466 676894
rect 260702 676658 260734 676894
rect 260114 676574 260734 676658
rect 260114 676338 260146 676574
rect 260382 676338 260466 676574
rect 260702 676338 260734 676574
rect 260114 657000 260734 676338
rect 261514 706758 262134 707750
rect 261514 706522 261546 706758
rect 261782 706522 261866 706758
rect 262102 706522 262134 706758
rect 261514 706438 262134 706522
rect 261514 706202 261546 706438
rect 261782 706202 261866 706438
rect 262102 706202 262134 706438
rect 261514 691174 262134 706202
rect 261514 690938 261546 691174
rect 261782 690938 261866 691174
rect 262102 690938 262134 691174
rect 261514 690854 262134 690938
rect 261514 690618 261546 690854
rect 261782 690618 261866 690854
rect 262102 690618 262134 690854
rect 261514 657000 262134 690618
rect 262914 705798 263534 705830
rect 262914 705562 262946 705798
rect 263182 705562 263266 705798
rect 263502 705562 263534 705798
rect 262914 705478 263534 705562
rect 262914 705242 262946 705478
rect 263182 705242 263266 705478
rect 263502 705242 263534 705478
rect 262914 669454 263534 705242
rect 262914 669218 262946 669454
rect 263182 669218 263266 669454
rect 263502 669218 263534 669454
rect 262914 669134 263534 669218
rect 262914 668898 262946 669134
rect 263182 668898 263266 669134
rect 263502 668898 263534 669134
rect 262914 657000 263534 668898
rect 263834 680614 264454 711002
rect 268954 710598 269574 711590
rect 268954 710362 268986 710598
rect 269222 710362 269306 710598
rect 269542 710362 269574 710598
rect 268954 710278 269574 710362
rect 268954 710042 268986 710278
rect 269222 710042 269306 710278
rect 269542 710042 269574 710278
rect 263834 680378 263866 680614
rect 264102 680378 264186 680614
rect 264422 680378 264454 680614
rect 263834 680294 264454 680378
rect 263834 680058 263866 680294
rect 264102 680058 264186 680294
rect 264422 680058 264454 680294
rect 263834 657000 264454 680058
rect 265234 708678 265854 709670
rect 265234 708442 265266 708678
rect 265502 708442 265586 708678
rect 265822 708442 265854 708678
rect 265234 708358 265854 708442
rect 265234 708122 265266 708358
rect 265502 708122 265586 708358
rect 265822 708122 265854 708358
rect 265234 694894 265854 708122
rect 265234 694658 265266 694894
rect 265502 694658 265586 694894
rect 265822 694658 265854 694894
rect 265234 694574 265854 694658
rect 265234 694338 265266 694574
rect 265502 694338 265586 694574
rect 265822 694338 265854 694574
rect 265234 658894 265854 694338
rect 265234 658658 265266 658894
rect 265502 658658 265586 658894
rect 265822 658658 265854 658894
rect 265234 658574 265854 658658
rect 265234 658338 265266 658574
rect 265502 658338 265586 658574
rect 265822 658338 265854 658574
rect 265234 657000 265854 658338
rect 266634 707718 267254 707750
rect 266634 707482 266666 707718
rect 266902 707482 266986 707718
rect 267222 707482 267254 707718
rect 266634 707398 267254 707482
rect 266634 707162 266666 707398
rect 266902 707162 266986 707398
rect 267222 707162 267254 707398
rect 266634 673174 267254 707162
rect 266634 672938 266666 673174
rect 266902 672938 266986 673174
rect 267222 672938 267254 673174
rect 266634 672854 267254 672938
rect 266634 672618 266666 672854
rect 266902 672618 266986 672854
rect 267222 672618 267254 672854
rect 266634 657000 267254 672618
rect 268034 704838 268654 705830
rect 268034 704602 268066 704838
rect 268302 704602 268386 704838
rect 268622 704602 268654 704838
rect 268034 704518 268654 704602
rect 268034 704282 268066 704518
rect 268302 704282 268386 704518
rect 268622 704282 268654 704518
rect 268034 687454 268654 704282
rect 268034 687218 268066 687454
rect 268302 687218 268386 687454
rect 268622 687218 268654 687454
rect 268034 687134 268654 687218
rect 268034 686898 268066 687134
rect 268302 686898 268386 687134
rect 268622 686898 268654 687134
rect 268034 657000 268654 686898
rect 268954 698614 269574 710042
rect 274074 711558 274694 711590
rect 274074 711322 274106 711558
rect 274342 711322 274426 711558
rect 274662 711322 274694 711558
rect 274074 711238 274694 711322
rect 274074 711002 274106 711238
rect 274342 711002 274426 711238
rect 274662 711002 274694 711238
rect 268954 698378 268986 698614
rect 269222 698378 269306 698614
rect 269542 698378 269574 698614
rect 268954 698294 269574 698378
rect 268954 698058 268986 698294
rect 269222 698058 269306 698294
rect 269542 698058 269574 698294
rect 268954 662614 269574 698058
rect 268954 662378 268986 662614
rect 269222 662378 269306 662614
rect 269542 662378 269574 662614
rect 268954 662294 269574 662378
rect 268954 662058 268986 662294
rect 269222 662058 269306 662294
rect 269542 662058 269574 662294
rect 268954 657000 269574 662058
rect 270354 709638 270974 709670
rect 270354 709402 270386 709638
rect 270622 709402 270706 709638
rect 270942 709402 270974 709638
rect 270354 709318 270974 709402
rect 270354 709082 270386 709318
rect 270622 709082 270706 709318
rect 270942 709082 270974 709318
rect 270354 676894 270974 709082
rect 270354 676658 270386 676894
rect 270622 676658 270706 676894
rect 270942 676658 270974 676894
rect 270354 676574 270974 676658
rect 270354 676338 270386 676574
rect 270622 676338 270706 676574
rect 270942 676338 270974 676574
rect 270354 657000 270974 676338
rect 271754 706758 272374 707750
rect 271754 706522 271786 706758
rect 272022 706522 272106 706758
rect 272342 706522 272374 706758
rect 271754 706438 272374 706522
rect 271754 706202 271786 706438
rect 272022 706202 272106 706438
rect 272342 706202 272374 706438
rect 271754 691174 272374 706202
rect 271754 690938 271786 691174
rect 272022 690938 272106 691174
rect 272342 690938 272374 691174
rect 271754 690854 272374 690938
rect 271754 690618 271786 690854
rect 272022 690618 272106 690854
rect 272342 690618 272374 690854
rect 271754 657000 272374 690618
rect 273154 705798 273774 705830
rect 273154 705562 273186 705798
rect 273422 705562 273506 705798
rect 273742 705562 273774 705798
rect 273154 705478 273774 705562
rect 273154 705242 273186 705478
rect 273422 705242 273506 705478
rect 273742 705242 273774 705478
rect 273154 669454 273774 705242
rect 273154 669218 273186 669454
rect 273422 669218 273506 669454
rect 273742 669218 273774 669454
rect 273154 669134 273774 669218
rect 273154 668898 273186 669134
rect 273422 668898 273506 669134
rect 273742 668898 273774 669134
rect 273154 657000 273774 668898
rect 274074 680614 274694 711002
rect 279194 710598 279814 711590
rect 279194 710362 279226 710598
rect 279462 710362 279546 710598
rect 279782 710362 279814 710598
rect 279194 710278 279814 710362
rect 279194 710042 279226 710278
rect 279462 710042 279546 710278
rect 279782 710042 279814 710278
rect 274074 680378 274106 680614
rect 274342 680378 274426 680614
rect 274662 680378 274694 680614
rect 274074 680294 274694 680378
rect 274074 680058 274106 680294
rect 274342 680058 274426 680294
rect 274662 680058 274694 680294
rect 274074 657000 274694 680058
rect 275474 708678 276094 709670
rect 275474 708442 275506 708678
rect 275742 708442 275826 708678
rect 276062 708442 276094 708678
rect 275474 708358 276094 708442
rect 275474 708122 275506 708358
rect 275742 708122 275826 708358
rect 276062 708122 276094 708358
rect 275474 694894 276094 708122
rect 275474 694658 275506 694894
rect 275742 694658 275826 694894
rect 276062 694658 276094 694894
rect 275474 694574 276094 694658
rect 275474 694338 275506 694574
rect 275742 694338 275826 694574
rect 276062 694338 276094 694574
rect 275474 658894 276094 694338
rect 275474 658658 275506 658894
rect 275742 658658 275826 658894
rect 276062 658658 276094 658894
rect 275474 658574 276094 658658
rect 275474 658338 275506 658574
rect 275742 658338 275826 658574
rect 276062 658338 276094 658574
rect 275474 657000 276094 658338
rect 276874 707718 277494 707750
rect 276874 707482 276906 707718
rect 277142 707482 277226 707718
rect 277462 707482 277494 707718
rect 276874 707398 277494 707482
rect 276874 707162 276906 707398
rect 277142 707162 277226 707398
rect 277462 707162 277494 707398
rect 276874 673174 277494 707162
rect 276874 672938 276906 673174
rect 277142 672938 277226 673174
rect 277462 672938 277494 673174
rect 276874 672854 277494 672938
rect 276874 672618 276906 672854
rect 277142 672618 277226 672854
rect 277462 672618 277494 672854
rect 276874 657000 277494 672618
rect 278274 704838 278894 705830
rect 278274 704602 278306 704838
rect 278542 704602 278626 704838
rect 278862 704602 278894 704838
rect 278274 704518 278894 704602
rect 278274 704282 278306 704518
rect 278542 704282 278626 704518
rect 278862 704282 278894 704518
rect 278274 687454 278894 704282
rect 278274 687218 278306 687454
rect 278542 687218 278626 687454
rect 278862 687218 278894 687454
rect 278274 687134 278894 687218
rect 278274 686898 278306 687134
rect 278542 686898 278626 687134
rect 278862 686898 278894 687134
rect 278274 657000 278894 686898
rect 279194 698614 279814 710042
rect 284314 711558 284934 711590
rect 284314 711322 284346 711558
rect 284582 711322 284666 711558
rect 284902 711322 284934 711558
rect 284314 711238 284934 711322
rect 284314 711002 284346 711238
rect 284582 711002 284666 711238
rect 284902 711002 284934 711238
rect 279194 698378 279226 698614
rect 279462 698378 279546 698614
rect 279782 698378 279814 698614
rect 279194 698294 279814 698378
rect 279194 698058 279226 698294
rect 279462 698058 279546 698294
rect 279782 698058 279814 698294
rect 279194 662614 279814 698058
rect 279194 662378 279226 662614
rect 279462 662378 279546 662614
rect 279782 662378 279814 662614
rect 279194 662294 279814 662378
rect 279194 662058 279226 662294
rect 279462 662058 279546 662294
rect 279782 662058 279814 662294
rect 279194 657000 279814 662058
rect 280594 709638 281214 709670
rect 280594 709402 280626 709638
rect 280862 709402 280946 709638
rect 281182 709402 281214 709638
rect 280594 709318 281214 709402
rect 280594 709082 280626 709318
rect 280862 709082 280946 709318
rect 281182 709082 281214 709318
rect 280594 676894 281214 709082
rect 280594 676658 280626 676894
rect 280862 676658 280946 676894
rect 281182 676658 281214 676894
rect 280594 676574 281214 676658
rect 280594 676338 280626 676574
rect 280862 676338 280946 676574
rect 281182 676338 281214 676574
rect 280594 657000 281214 676338
rect 281994 706758 282614 707750
rect 281994 706522 282026 706758
rect 282262 706522 282346 706758
rect 282582 706522 282614 706758
rect 281994 706438 282614 706522
rect 281994 706202 282026 706438
rect 282262 706202 282346 706438
rect 282582 706202 282614 706438
rect 281994 691174 282614 706202
rect 281994 690938 282026 691174
rect 282262 690938 282346 691174
rect 282582 690938 282614 691174
rect 281994 690854 282614 690938
rect 281994 690618 282026 690854
rect 282262 690618 282346 690854
rect 282582 690618 282614 690854
rect 281994 657000 282614 690618
rect 283394 705798 284014 705830
rect 283394 705562 283426 705798
rect 283662 705562 283746 705798
rect 283982 705562 284014 705798
rect 283394 705478 284014 705562
rect 283394 705242 283426 705478
rect 283662 705242 283746 705478
rect 283982 705242 284014 705478
rect 283394 669454 284014 705242
rect 283394 669218 283426 669454
rect 283662 669218 283746 669454
rect 283982 669218 284014 669454
rect 283394 669134 284014 669218
rect 283394 668898 283426 669134
rect 283662 668898 283746 669134
rect 283982 668898 284014 669134
rect 283394 657000 284014 668898
rect 284314 680614 284934 711002
rect 289434 710598 290054 711590
rect 289434 710362 289466 710598
rect 289702 710362 289786 710598
rect 290022 710362 290054 710598
rect 289434 710278 290054 710362
rect 289434 710042 289466 710278
rect 289702 710042 289786 710278
rect 290022 710042 290054 710278
rect 284314 680378 284346 680614
rect 284582 680378 284666 680614
rect 284902 680378 284934 680614
rect 284314 680294 284934 680378
rect 284314 680058 284346 680294
rect 284582 680058 284666 680294
rect 284902 680058 284934 680294
rect 284314 657000 284934 680058
rect 285714 708678 286334 709670
rect 285714 708442 285746 708678
rect 285982 708442 286066 708678
rect 286302 708442 286334 708678
rect 285714 708358 286334 708442
rect 285714 708122 285746 708358
rect 285982 708122 286066 708358
rect 286302 708122 286334 708358
rect 285714 694894 286334 708122
rect 285714 694658 285746 694894
rect 285982 694658 286066 694894
rect 286302 694658 286334 694894
rect 285714 694574 286334 694658
rect 285714 694338 285746 694574
rect 285982 694338 286066 694574
rect 286302 694338 286334 694574
rect 285714 658894 286334 694338
rect 285714 658658 285746 658894
rect 285982 658658 286066 658894
rect 286302 658658 286334 658894
rect 285714 658574 286334 658658
rect 285714 658338 285746 658574
rect 285982 658338 286066 658574
rect 286302 658338 286334 658574
rect 285714 657000 286334 658338
rect 287114 707718 287734 707750
rect 287114 707482 287146 707718
rect 287382 707482 287466 707718
rect 287702 707482 287734 707718
rect 287114 707398 287734 707482
rect 287114 707162 287146 707398
rect 287382 707162 287466 707398
rect 287702 707162 287734 707398
rect 287114 673174 287734 707162
rect 287114 672938 287146 673174
rect 287382 672938 287466 673174
rect 287702 672938 287734 673174
rect 287114 672854 287734 672938
rect 287114 672618 287146 672854
rect 287382 672618 287466 672854
rect 287702 672618 287734 672854
rect 287114 657000 287734 672618
rect 288514 704838 289134 705830
rect 288514 704602 288546 704838
rect 288782 704602 288866 704838
rect 289102 704602 289134 704838
rect 288514 704518 289134 704602
rect 288514 704282 288546 704518
rect 288782 704282 288866 704518
rect 289102 704282 289134 704518
rect 288514 687454 289134 704282
rect 288514 687218 288546 687454
rect 288782 687218 288866 687454
rect 289102 687218 289134 687454
rect 288514 687134 289134 687218
rect 288514 686898 288546 687134
rect 288782 686898 288866 687134
rect 289102 686898 289134 687134
rect 288514 657000 289134 686898
rect 289434 698614 290054 710042
rect 294554 711558 295174 711590
rect 294554 711322 294586 711558
rect 294822 711322 294906 711558
rect 295142 711322 295174 711558
rect 294554 711238 295174 711322
rect 294554 711002 294586 711238
rect 294822 711002 294906 711238
rect 295142 711002 295174 711238
rect 289434 698378 289466 698614
rect 289702 698378 289786 698614
rect 290022 698378 290054 698614
rect 289434 698294 290054 698378
rect 289434 698058 289466 698294
rect 289702 698058 289786 698294
rect 290022 698058 290054 698294
rect 289434 662614 290054 698058
rect 289434 662378 289466 662614
rect 289702 662378 289786 662614
rect 290022 662378 290054 662614
rect 289434 662294 290054 662378
rect 289434 662058 289466 662294
rect 289702 662058 289786 662294
rect 290022 662058 290054 662294
rect 289434 657000 290054 662058
rect 290834 709638 291454 709670
rect 290834 709402 290866 709638
rect 291102 709402 291186 709638
rect 291422 709402 291454 709638
rect 290834 709318 291454 709402
rect 290834 709082 290866 709318
rect 291102 709082 291186 709318
rect 291422 709082 291454 709318
rect 290834 676894 291454 709082
rect 290834 676658 290866 676894
rect 291102 676658 291186 676894
rect 291422 676658 291454 676894
rect 290834 676574 291454 676658
rect 290834 676338 290866 676574
rect 291102 676338 291186 676574
rect 291422 676338 291454 676574
rect 290834 657000 291454 676338
rect 292234 706758 292854 707750
rect 292234 706522 292266 706758
rect 292502 706522 292586 706758
rect 292822 706522 292854 706758
rect 292234 706438 292854 706522
rect 292234 706202 292266 706438
rect 292502 706202 292586 706438
rect 292822 706202 292854 706438
rect 292234 691174 292854 706202
rect 292234 690938 292266 691174
rect 292502 690938 292586 691174
rect 292822 690938 292854 691174
rect 292234 690854 292854 690938
rect 292234 690618 292266 690854
rect 292502 690618 292586 690854
rect 292822 690618 292854 690854
rect 292234 657000 292854 690618
rect 293634 705798 294254 705830
rect 293634 705562 293666 705798
rect 293902 705562 293986 705798
rect 294222 705562 294254 705798
rect 293634 705478 294254 705562
rect 293634 705242 293666 705478
rect 293902 705242 293986 705478
rect 294222 705242 294254 705478
rect 293634 669454 294254 705242
rect 293634 669218 293666 669454
rect 293902 669218 293986 669454
rect 294222 669218 294254 669454
rect 293634 669134 294254 669218
rect 293634 668898 293666 669134
rect 293902 668898 293986 669134
rect 294222 668898 294254 669134
rect 293634 657000 294254 668898
rect 294554 680614 295174 711002
rect 299674 710598 300294 711590
rect 299674 710362 299706 710598
rect 299942 710362 300026 710598
rect 300262 710362 300294 710598
rect 299674 710278 300294 710362
rect 299674 710042 299706 710278
rect 299942 710042 300026 710278
rect 300262 710042 300294 710278
rect 294554 680378 294586 680614
rect 294822 680378 294906 680614
rect 295142 680378 295174 680614
rect 294554 680294 295174 680378
rect 294554 680058 294586 680294
rect 294822 680058 294906 680294
rect 295142 680058 295174 680294
rect 294554 657000 295174 680058
rect 295954 708678 296574 709670
rect 295954 708442 295986 708678
rect 296222 708442 296306 708678
rect 296542 708442 296574 708678
rect 295954 708358 296574 708442
rect 295954 708122 295986 708358
rect 296222 708122 296306 708358
rect 296542 708122 296574 708358
rect 295954 694894 296574 708122
rect 295954 694658 295986 694894
rect 296222 694658 296306 694894
rect 296542 694658 296574 694894
rect 295954 694574 296574 694658
rect 295954 694338 295986 694574
rect 296222 694338 296306 694574
rect 296542 694338 296574 694574
rect 295954 658894 296574 694338
rect 295954 658658 295986 658894
rect 296222 658658 296306 658894
rect 296542 658658 296574 658894
rect 295954 658574 296574 658658
rect 295954 658338 295986 658574
rect 296222 658338 296306 658574
rect 296542 658338 296574 658574
rect 295954 657000 296574 658338
rect 297354 707718 297974 707750
rect 297354 707482 297386 707718
rect 297622 707482 297706 707718
rect 297942 707482 297974 707718
rect 297354 707398 297974 707482
rect 297354 707162 297386 707398
rect 297622 707162 297706 707398
rect 297942 707162 297974 707398
rect 297354 673174 297974 707162
rect 297354 672938 297386 673174
rect 297622 672938 297706 673174
rect 297942 672938 297974 673174
rect 297354 672854 297974 672938
rect 297354 672618 297386 672854
rect 297622 672618 297706 672854
rect 297942 672618 297974 672854
rect 297354 657000 297974 672618
rect 298754 704838 299374 705830
rect 298754 704602 298786 704838
rect 299022 704602 299106 704838
rect 299342 704602 299374 704838
rect 298754 704518 299374 704602
rect 298754 704282 298786 704518
rect 299022 704282 299106 704518
rect 299342 704282 299374 704518
rect 298754 687454 299374 704282
rect 298754 687218 298786 687454
rect 299022 687218 299106 687454
rect 299342 687218 299374 687454
rect 298754 687134 299374 687218
rect 298754 686898 298786 687134
rect 299022 686898 299106 687134
rect 299342 686898 299374 687134
rect 298754 657000 299374 686898
rect 299674 698614 300294 710042
rect 304794 711558 305414 711590
rect 304794 711322 304826 711558
rect 305062 711322 305146 711558
rect 305382 711322 305414 711558
rect 304794 711238 305414 711322
rect 304794 711002 304826 711238
rect 305062 711002 305146 711238
rect 305382 711002 305414 711238
rect 299674 698378 299706 698614
rect 299942 698378 300026 698614
rect 300262 698378 300294 698614
rect 299674 698294 300294 698378
rect 299674 698058 299706 698294
rect 299942 698058 300026 698294
rect 300262 698058 300294 698294
rect 299674 662614 300294 698058
rect 299674 662378 299706 662614
rect 299942 662378 300026 662614
rect 300262 662378 300294 662614
rect 299674 662294 300294 662378
rect 299674 662058 299706 662294
rect 299942 662058 300026 662294
rect 300262 662058 300294 662294
rect 299674 657000 300294 662058
rect 301074 709638 301694 709670
rect 301074 709402 301106 709638
rect 301342 709402 301426 709638
rect 301662 709402 301694 709638
rect 301074 709318 301694 709402
rect 301074 709082 301106 709318
rect 301342 709082 301426 709318
rect 301662 709082 301694 709318
rect 301074 676894 301694 709082
rect 301074 676658 301106 676894
rect 301342 676658 301426 676894
rect 301662 676658 301694 676894
rect 301074 676574 301694 676658
rect 301074 676338 301106 676574
rect 301342 676338 301426 676574
rect 301662 676338 301694 676574
rect 301074 657000 301694 676338
rect 302474 706758 303094 707750
rect 302474 706522 302506 706758
rect 302742 706522 302826 706758
rect 303062 706522 303094 706758
rect 302474 706438 303094 706522
rect 302474 706202 302506 706438
rect 302742 706202 302826 706438
rect 303062 706202 303094 706438
rect 302474 691174 303094 706202
rect 302474 690938 302506 691174
rect 302742 690938 302826 691174
rect 303062 690938 303094 691174
rect 302474 690854 303094 690938
rect 302474 690618 302506 690854
rect 302742 690618 302826 690854
rect 303062 690618 303094 690854
rect 302474 657000 303094 690618
rect 303874 705798 304494 705830
rect 303874 705562 303906 705798
rect 304142 705562 304226 705798
rect 304462 705562 304494 705798
rect 303874 705478 304494 705562
rect 303874 705242 303906 705478
rect 304142 705242 304226 705478
rect 304462 705242 304494 705478
rect 303874 669454 304494 705242
rect 303874 669218 303906 669454
rect 304142 669218 304226 669454
rect 304462 669218 304494 669454
rect 303874 669134 304494 669218
rect 303874 668898 303906 669134
rect 304142 668898 304226 669134
rect 304462 668898 304494 669134
rect 303874 657000 304494 668898
rect 304794 680614 305414 711002
rect 309914 710598 310534 711590
rect 309914 710362 309946 710598
rect 310182 710362 310266 710598
rect 310502 710362 310534 710598
rect 309914 710278 310534 710362
rect 309914 710042 309946 710278
rect 310182 710042 310266 710278
rect 310502 710042 310534 710278
rect 304794 680378 304826 680614
rect 305062 680378 305146 680614
rect 305382 680378 305414 680614
rect 304794 680294 305414 680378
rect 304794 680058 304826 680294
rect 305062 680058 305146 680294
rect 305382 680058 305414 680294
rect 304794 657000 305414 680058
rect 306194 708678 306814 709670
rect 306194 708442 306226 708678
rect 306462 708442 306546 708678
rect 306782 708442 306814 708678
rect 306194 708358 306814 708442
rect 306194 708122 306226 708358
rect 306462 708122 306546 708358
rect 306782 708122 306814 708358
rect 306194 694894 306814 708122
rect 306194 694658 306226 694894
rect 306462 694658 306546 694894
rect 306782 694658 306814 694894
rect 306194 694574 306814 694658
rect 306194 694338 306226 694574
rect 306462 694338 306546 694574
rect 306782 694338 306814 694574
rect 306194 658894 306814 694338
rect 306194 658658 306226 658894
rect 306462 658658 306546 658894
rect 306782 658658 306814 658894
rect 306194 658574 306814 658658
rect 306194 658338 306226 658574
rect 306462 658338 306546 658574
rect 306782 658338 306814 658574
rect 306194 657000 306814 658338
rect 307594 707718 308214 707750
rect 307594 707482 307626 707718
rect 307862 707482 307946 707718
rect 308182 707482 308214 707718
rect 307594 707398 308214 707482
rect 307594 707162 307626 707398
rect 307862 707162 307946 707398
rect 308182 707162 308214 707398
rect 307594 673174 308214 707162
rect 307594 672938 307626 673174
rect 307862 672938 307946 673174
rect 308182 672938 308214 673174
rect 307594 672854 308214 672938
rect 307594 672618 307626 672854
rect 307862 672618 307946 672854
rect 308182 672618 308214 672854
rect 307594 657000 308214 672618
rect 308994 704838 309614 705830
rect 308994 704602 309026 704838
rect 309262 704602 309346 704838
rect 309582 704602 309614 704838
rect 308994 704518 309614 704602
rect 308994 704282 309026 704518
rect 309262 704282 309346 704518
rect 309582 704282 309614 704518
rect 308994 687454 309614 704282
rect 308994 687218 309026 687454
rect 309262 687218 309346 687454
rect 309582 687218 309614 687454
rect 308994 687134 309614 687218
rect 308994 686898 309026 687134
rect 309262 686898 309346 687134
rect 309582 686898 309614 687134
rect 308994 657000 309614 686898
rect 309914 698614 310534 710042
rect 315034 711558 315654 711590
rect 315034 711322 315066 711558
rect 315302 711322 315386 711558
rect 315622 711322 315654 711558
rect 315034 711238 315654 711322
rect 315034 711002 315066 711238
rect 315302 711002 315386 711238
rect 315622 711002 315654 711238
rect 309914 698378 309946 698614
rect 310182 698378 310266 698614
rect 310502 698378 310534 698614
rect 309914 698294 310534 698378
rect 309914 698058 309946 698294
rect 310182 698058 310266 698294
rect 310502 698058 310534 698294
rect 309914 662614 310534 698058
rect 309914 662378 309946 662614
rect 310182 662378 310266 662614
rect 310502 662378 310534 662614
rect 309914 662294 310534 662378
rect 309914 662058 309946 662294
rect 310182 662058 310266 662294
rect 310502 662058 310534 662294
rect 309914 657000 310534 662058
rect 311314 709638 311934 709670
rect 311314 709402 311346 709638
rect 311582 709402 311666 709638
rect 311902 709402 311934 709638
rect 311314 709318 311934 709402
rect 311314 709082 311346 709318
rect 311582 709082 311666 709318
rect 311902 709082 311934 709318
rect 311314 676894 311934 709082
rect 311314 676658 311346 676894
rect 311582 676658 311666 676894
rect 311902 676658 311934 676894
rect 311314 676574 311934 676658
rect 311314 676338 311346 676574
rect 311582 676338 311666 676574
rect 311902 676338 311934 676574
rect 311314 657000 311934 676338
rect 312714 706758 313334 707750
rect 312714 706522 312746 706758
rect 312982 706522 313066 706758
rect 313302 706522 313334 706758
rect 312714 706438 313334 706522
rect 312714 706202 312746 706438
rect 312982 706202 313066 706438
rect 313302 706202 313334 706438
rect 312714 691174 313334 706202
rect 312714 690938 312746 691174
rect 312982 690938 313066 691174
rect 313302 690938 313334 691174
rect 312714 690854 313334 690938
rect 312714 690618 312746 690854
rect 312982 690618 313066 690854
rect 313302 690618 313334 690854
rect 312714 657000 313334 690618
rect 314114 705798 314734 705830
rect 314114 705562 314146 705798
rect 314382 705562 314466 705798
rect 314702 705562 314734 705798
rect 314114 705478 314734 705562
rect 314114 705242 314146 705478
rect 314382 705242 314466 705478
rect 314702 705242 314734 705478
rect 314114 669454 314734 705242
rect 314114 669218 314146 669454
rect 314382 669218 314466 669454
rect 314702 669218 314734 669454
rect 314114 669134 314734 669218
rect 314114 668898 314146 669134
rect 314382 668898 314466 669134
rect 314702 668898 314734 669134
rect 314114 657000 314734 668898
rect 315034 680614 315654 711002
rect 320154 710598 320774 711590
rect 320154 710362 320186 710598
rect 320422 710362 320506 710598
rect 320742 710362 320774 710598
rect 320154 710278 320774 710362
rect 320154 710042 320186 710278
rect 320422 710042 320506 710278
rect 320742 710042 320774 710278
rect 315034 680378 315066 680614
rect 315302 680378 315386 680614
rect 315622 680378 315654 680614
rect 315034 680294 315654 680378
rect 315034 680058 315066 680294
rect 315302 680058 315386 680294
rect 315622 680058 315654 680294
rect 315034 657000 315654 680058
rect 316434 708678 317054 709670
rect 316434 708442 316466 708678
rect 316702 708442 316786 708678
rect 317022 708442 317054 708678
rect 316434 708358 317054 708442
rect 316434 708122 316466 708358
rect 316702 708122 316786 708358
rect 317022 708122 317054 708358
rect 316434 694894 317054 708122
rect 316434 694658 316466 694894
rect 316702 694658 316786 694894
rect 317022 694658 317054 694894
rect 316434 694574 317054 694658
rect 316434 694338 316466 694574
rect 316702 694338 316786 694574
rect 317022 694338 317054 694574
rect 316434 658894 317054 694338
rect 316434 658658 316466 658894
rect 316702 658658 316786 658894
rect 317022 658658 317054 658894
rect 316434 658574 317054 658658
rect 316434 658338 316466 658574
rect 316702 658338 316786 658574
rect 317022 658338 317054 658574
rect 316434 657000 317054 658338
rect 317834 707718 318454 707750
rect 317834 707482 317866 707718
rect 318102 707482 318186 707718
rect 318422 707482 318454 707718
rect 317834 707398 318454 707482
rect 317834 707162 317866 707398
rect 318102 707162 318186 707398
rect 318422 707162 318454 707398
rect 317834 673174 318454 707162
rect 317834 672938 317866 673174
rect 318102 672938 318186 673174
rect 318422 672938 318454 673174
rect 317834 672854 318454 672938
rect 317834 672618 317866 672854
rect 318102 672618 318186 672854
rect 318422 672618 318454 672854
rect 317834 657000 318454 672618
rect 319234 704838 319854 705830
rect 319234 704602 319266 704838
rect 319502 704602 319586 704838
rect 319822 704602 319854 704838
rect 319234 704518 319854 704602
rect 319234 704282 319266 704518
rect 319502 704282 319586 704518
rect 319822 704282 319854 704518
rect 319234 687454 319854 704282
rect 319234 687218 319266 687454
rect 319502 687218 319586 687454
rect 319822 687218 319854 687454
rect 319234 687134 319854 687218
rect 319234 686898 319266 687134
rect 319502 686898 319586 687134
rect 319822 686898 319854 687134
rect 319234 657000 319854 686898
rect 320154 698614 320774 710042
rect 325274 711558 325894 711590
rect 325274 711322 325306 711558
rect 325542 711322 325626 711558
rect 325862 711322 325894 711558
rect 325274 711238 325894 711322
rect 325274 711002 325306 711238
rect 325542 711002 325626 711238
rect 325862 711002 325894 711238
rect 320154 698378 320186 698614
rect 320422 698378 320506 698614
rect 320742 698378 320774 698614
rect 320154 698294 320774 698378
rect 320154 698058 320186 698294
rect 320422 698058 320506 698294
rect 320742 698058 320774 698294
rect 320154 662614 320774 698058
rect 320154 662378 320186 662614
rect 320422 662378 320506 662614
rect 320742 662378 320774 662614
rect 320154 662294 320774 662378
rect 320154 662058 320186 662294
rect 320422 662058 320506 662294
rect 320742 662058 320774 662294
rect 320154 657000 320774 662058
rect 321554 709638 322174 709670
rect 321554 709402 321586 709638
rect 321822 709402 321906 709638
rect 322142 709402 322174 709638
rect 321554 709318 322174 709402
rect 321554 709082 321586 709318
rect 321822 709082 321906 709318
rect 322142 709082 322174 709318
rect 321554 676894 322174 709082
rect 321554 676658 321586 676894
rect 321822 676658 321906 676894
rect 322142 676658 322174 676894
rect 321554 676574 322174 676658
rect 321554 676338 321586 676574
rect 321822 676338 321906 676574
rect 322142 676338 322174 676574
rect 321554 657000 322174 676338
rect 322954 706758 323574 707750
rect 322954 706522 322986 706758
rect 323222 706522 323306 706758
rect 323542 706522 323574 706758
rect 322954 706438 323574 706522
rect 322954 706202 322986 706438
rect 323222 706202 323306 706438
rect 323542 706202 323574 706438
rect 322954 691174 323574 706202
rect 322954 690938 322986 691174
rect 323222 690938 323306 691174
rect 323542 690938 323574 691174
rect 322954 690854 323574 690938
rect 322954 690618 322986 690854
rect 323222 690618 323306 690854
rect 323542 690618 323574 690854
rect 322954 657000 323574 690618
rect 324354 705798 324974 705830
rect 324354 705562 324386 705798
rect 324622 705562 324706 705798
rect 324942 705562 324974 705798
rect 324354 705478 324974 705562
rect 324354 705242 324386 705478
rect 324622 705242 324706 705478
rect 324942 705242 324974 705478
rect 324354 669454 324974 705242
rect 324354 669218 324386 669454
rect 324622 669218 324706 669454
rect 324942 669218 324974 669454
rect 324354 669134 324974 669218
rect 324354 668898 324386 669134
rect 324622 668898 324706 669134
rect 324942 668898 324974 669134
rect 324354 657000 324974 668898
rect 325274 680614 325894 711002
rect 330394 710598 331014 711590
rect 330394 710362 330426 710598
rect 330662 710362 330746 710598
rect 330982 710362 331014 710598
rect 330394 710278 331014 710362
rect 330394 710042 330426 710278
rect 330662 710042 330746 710278
rect 330982 710042 331014 710278
rect 325274 680378 325306 680614
rect 325542 680378 325626 680614
rect 325862 680378 325894 680614
rect 325274 680294 325894 680378
rect 325274 680058 325306 680294
rect 325542 680058 325626 680294
rect 325862 680058 325894 680294
rect 325274 657000 325894 680058
rect 326674 708678 327294 709670
rect 326674 708442 326706 708678
rect 326942 708442 327026 708678
rect 327262 708442 327294 708678
rect 326674 708358 327294 708442
rect 326674 708122 326706 708358
rect 326942 708122 327026 708358
rect 327262 708122 327294 708358
rect 326674 694894 327294 708122
rect 326674 694658 326706 694894
rect 326942 694658 327026 694894
rect 327262 694658 327294 694894
rect 326674 694574 327294 694658
rect 326674 694338 326706 694574
rect 326942 694338 327026 694574
rect 327262 694338 327294 694574
rect 326674 658894 327294 694338
rect 326674 658658 326706 658894
rect 326942 658658 327026 658894
rect 327262 658658 327294 658894
rect 326674 658574 327294 658658
rect 326674 658338 326706 658574
rect 326942 658338 327026 658574
rect 327262 658338 327294 658574
rect 326674 657000 327294 658338
rect 328074 707718 328694 707750
rect 328074 707482 328106 707718
rect 328342 707482 328426 707718
rect 328662 707482 328694 707718
rect 328074 707398 328694 707482
rect 328074 707162 328106 707398
rect 328342 707162 328426 707398
rect 328662 707162 328694 707398
rect 328074 673174 328694 707162
rect 328074 672938 328106 673174
rect 328342 672938 328426 673174
rect 328662 672938 328694 673174
rect 328074 672854 328694 672938
rect 328074 672618 328106 672854
rect 328342 672618 328426 672854
rect 328662 672618 328694 672854
rect 328074 657000 328694 672618
rect 329474 704838 330094 705830
rect 329474 704602 329506 704838
rect 329742 704602 329826 704838
rect 330062 704602 330094 704838
rect 329474 704518 330094 704602
rect 329474 704282 329506 704518
rect 329742 704282 329826 704518
rect 330062 704282 330094 704518
rect 329474 687454 330094 704282
rect 329474 687218 329506 687454
rect 329742 687218 329826 687454
rect 330062 687218 330094 687454
rect 329474 687134 330094 687218
rect 329474 686898 329506 687134
rect 329742 686898 329826 687134
rect 330062 686898 330094 687134
rect 329474 657000 330094 686898
rect 330394 698614 331014 710042
rect 335514 711558 336134 711590
rect 335514 711322 335546 711558
rect 335782 711322 335866 711558
rect 336102 711322 336134 711558
rect 335514 711238 336134 711322
rect 335514 711002 335546 711238
rect 335782 711002 335866 711238
rect 336102 711002 336134 711238
rect 330394 698378 330426 698614
rect 330662 698378 330746 698614
rect 330982 698378 331014 698614
rect 330394 698294 331014 698378
rect 330394 698058 330426 698294
rect 330662 698058 330746 698294
rect 330982 698058 331014 698294
rect 330394 662614 331014 698058
rect 330394 662378 330426 662614
rect 330662 662378 330746 662614
rect 330982 662378 331014 662614
rect 330394 662294 331014 662378
rect 330394 662058 330426 662294
rect 330662 662058 330746 662294
rect 330982 662058 331014 662294
rect 330394 657000 331014 662058
rect 331794 709638 332414 709670
rect 331794 709402 331826 709638
rect 332062 709402 332146 709638
rect 332382 709402 332414 709638
rect 331794 709318 332414 709402
rect 331794 709082 331826 709318
rect 332062 709082 332146 709318
rect 332382 709082 332414 709318
rect 331794 676894 332414 709082
rect 331794 676658 331826 676894
rect 332062 676658 332146 676894
rect 332382 676658 332414 676894
rect 331794 676574 332414 676658
rect 331794 676338 331826 676574
rect 332062 676338 332146 676574
rect 332382 676338 332414 676574
rect 331794 657000 332414 676338
rect 333194 706758 333814 707750
rect 333194 706522 333226 706758
rect 333462 706522 333546 706758
rect 333782 706522 333814 706758
rect 333194 706438 333814 706522
rect 333194 706202 333226 706438
rect 333462 706202 333546 706438
rect 333782 706202 333814 706438
rect 333194 691174 333814 706202
rect 333194 690938 333226 691174
rect 333462 690938 333546 691174
rect 333782 690938 333814 691174
rect 333194 690854 333814 690938
rect 333194 690618 333226 690854
rect 333462 690618 333546 690854
rect 333782 690618 333814 690854
rect 333194 657000 333814 690618
rect 334594 705798 335214 705830
rect 334594 705562 334626 705798
rect 334862 705562 334946 705798
rect 335182 705562 335214 705798
rect 334594 705478 335214 705562
rect 334594 705242 334626 705478
rect 334862 705242 334946 705478
rect 335182 705242 335214 705478
rect 334594 669454 335214 705242
rect 334594 669218 334626 669454
rect 334862 669218 334946 669454
rect 335182 669218 335214 669454
rect 334594 669134 335214 669218
rect 334594 668898 334626 669134
rect 334862 668898 334946 669134
rect 335182 668898 335214 669134
rect 334594 657000 335214 668898
rect 335514 680614 336134 711002
rect 340634 710598 341254 711590
rect 340634 710362 340666 710598
rect 340902 710362 340986 710598
rect 341222 710362 341254 710598
rect 340634 710278 341254 710362
rect 340634 710042 340666 710278
rect 340902 710042 340986 710278
rect 341222 710042 341254 710278
rect 335514 680378 335546 680614
rect 335782 680378 335866 680614
rect 336102 680378 336134 680614
rect 335514 680294 336134 680378
rect 335514 680058 335546 680294
rect 335782 680058 335866 680294
rect 336102 680058 336134 680294
rect 335514 657000 336134 680058
rect 336914 708678 337534 709670
rect 336914 708442 336946 708678
rect 337182 708442 337266 708678
rect 337502 708442 337534 708678
rect 336914 708358 337534 708442
rect 336914 708122 336946 708358
rect 337182 708122 337266 708358
rect 337502 708122 337534 708358
rect 336914 694894 337534 708122
rect 336914 694658 336946 694894
rect 337182 694658 337266 694894
rect 337502 694658 337534 694894
rect 336914 694574 337534 694658
rect 336914 694338 336946 694574
rect 337182 694338 337266 694574
rect 337502 694338 337534 694574
rect 336914 658894 337534 694338
rect 336914 658658 336946 658894
rect 337182 658658 337266 658894
rect 337502 658658 337534 658894
rect 336914 658574 337534 658658
rect 336914 658338 336946 658574
rect 337182 658338 337266 658574
rect 337502 658338 337534 658574
rect 336914 657000 337534 658338
rect 338314 707718 338934 707750
rect 338314 707482 338346 707718
rect 338582 707482 338666 707718
rect 338902 707482 338934 707718
rect 338314 707398 338934 707482
rect 338314 707162 338346 707398
rect 338582 707162 338666 707398
rect 338902 707162 338934 707398
rect 338314 673174 338934 707162
rect 338314 672938 338346 673174
rect 338582 672938 338666 673174
rect 338902 672938 338934 673174
rect 338314 672854 338934 672938
rect 338314 672618 338346 672854
rect 338582 672618 338666 672854
rect 338902 672618 338934 672854
rect 338314 657000 338934 672618
rect 339714 704838 340334 705830
rect 339714 704602 339746 704838
rect 339982 704602 340066 704838
rect 340302 704602 340334 704838
rect 339714 704518 340334 704602
rect 339714 704282 339746 704518
rect 339982 704282 340066 704518
rect 340302 704282 340334 704518
rect 339714 687454 340334 704282
rect 339714 687218 339746 687454
rect 339982 687218 340066 687454
rect 340302 687218 340334 687454
rect 339714 687134 340334 687218
rect 339714 686898 339746 687134
rect 339982 686898 340066 687134
rect 340302 686898 340334 687134
rect 339714 657000 340334 686898
rect 340634 698614 341254 710042
rect 345754 711558 346374 711590
rect 345754 711322 345786 711558
rect 346022 711322 346106 711558
rect 346342 711322 346374 711558
rect 345754 711238 346374 711322
rect 345754 711002 345786 711238
rect 346022 711002 346106 711238
rect 346342 711002 346374 711238
rect 340634 698378 340666 698614
rect 340902 698378 340986 698614
rect 341222 698378 341254 698614
rect 340634 698294 341254 698378
rect 340634 698058 340666 698294
rect 340902 698058 340986 698294
rect 341222 698058 341254 698294
rect 340634 662614 341254 698058
rect 340634 662378 340666 662614
rect 340902 662378 340986 662614
rect 341222 662378 341254 662614
rect 340634 662294 341254 662378
rect 340634 662058 340666 662294
rect 340902 662058 340986 662294
rect 341222 662058 341254 662294
rect 340634 657000 341254 662058
rect 342034 709638 342654 709670
rect 342034 709402 342066 709638
rect 342302 709402 342386 709638
rect 342622 709402 342654 709638
rect 342034 709318 342654 709402
rect 342034 709082 342066 709318
rect 342302 709082 342386 709318
rect 342622 709082 342654 709318
rect 342034 676894 342654 709082
rect 342034 676658 342066 676894
rect 342302 676658 342386 676894
rect 342622 676658 342654 676894
rect 342034 676574 342654 676658
rect 342034 676338 342066 676574
rect 342302 676338 342386 676574
rect 342622 676338 342654 676574
rect 342034 657000 342654 676338
rect 343434 706758 344054 707750
rect 343434 706522 343466 706758
rect 343702 706522 343786 706758
rect 344022 706522 344054 706758
rect 343434 706438 344054 706522
rect 343434 706202 343466 706438
rect 343702 706202 343786 706438
rect 344022 706202 344054 706438
rect 343434 691174 344054 706202
rect 343434 690938 343466 691174
rect 343702 690938 343786 691174
rect 344022 690938 344054 691174
rect 343434 690854 344054 690938
rect 343434 690618 343466 690854
rect 343702 690618 343786 690854
rect 344022 690618 344054 690854
rect 343434 657000 344054 690618
rect 344834 705798 345454 705830
rect 344834 705562 344866 705798
rect 345102 705562 345186 705798
rect 345422 705562 345454 705798
rect 344834 705478 345454 705562
rect 344834 705242 344866 705478
rect 345102 705242 345186 705478
rect 345422 705242 345454 705478
rect 344834 669454 345454 705242
rect 344834 669218 344866 669454
rect 345102 669218 345186 669454
rect 345422 669218 345454 669454
rect 344834 669134 345454 669218
rect 344834 668898 344866 669134
rect 345102 668898 345186 669134
rect 345422 668898 345454 669134
rect 344834 657000 345454 668898
rect 345754 680614 346374 711002
rect 350874 710598 351494 711590
rect 350874 710362 350906 710598
rect 351142 710362 351226 710598
rect 351462 710362 351494 710598
rect 350874 710278 351494 710362
rect 350874 710042 350906 710278
rect 351142 710042 351226 710278
rect 351462 710042 351494 710278
rect 345754 680378 345786 680614
rect 346022 680378 346106 680614
rect 346342 680378 346374 680614
rect 345754 680294 346374 680378
rect 345754 680058 345786 680294
rect 346022 680058 346106 680294
rect 346342 680058 346374 680294
rect 345754 657000 346374 680058
rect 347154 708678 347774 709670
rect 347154 708442 347186 708678
rect 347422 708442 347506 708678
rect 347742 708442 347774 708678
rect 347154 708358 347774 708442
rect 347154 708122 347186 708358
rect 347422 708122 347506 708358
rect 347742 708122 347774 708358
rect 347154 694894 347774 708122
rect 347154 694658 347186 694894
rect 347422 694658 347506 694894
rect 347742 694658 347774 694894
rect 347154 694574 347774 694658
rect 347154 694338 347186 694574
rect 347422 694338 347506 694574
rect 347742 694338 347774 694574
rect 347154 658894 347774 694338
rect 347154 658658 347186 658894
rect 347422 658658 347506 658894
rect 347742 658658 347774 658894
rect 347154 658574 347774 658658
rect 347154 658338 347186 658574
rect 347422 658338 347506 658574
rect 347742 658338 347774 658574
rect 347154 657000 347774 658338
rect 348554 707718 349174 707750
rect 348554 707482 348586 707718
rect 348822 707482 348906 707718
rect 349142 707482 349174 707718
rect 348554 707398 349174 707482
rect 348554 707162 348586 707398
rect 348822 707162 348906 707398
rect 349142 707162 349174 707398
rect 348554 673174 349174 707162
rect 348554 672938 348586 673174
rect 348822 672938 348906 673174
rect 349142 672938 349174 673174
rect 348554 672854 349174 672938
rect 348554 672618 348586 672854
rect 348822 672618 348906 672854
rect 349142 672618 349174 672854
rect 348554 657000 349174 672618
rect 349954 704838 350574 705830
rect 349954 704602 349986 704838
rect 350222 704602 350306 704838
rect 350542 704602 350574 704838
rect 349954 704518 350574 704602
rect 349954 704282 349986 704518
rect 350222 704282 350306 704518
rect 350542 704282 350574 704518
rect 349954 687454 350574 704282
rect 349954 687218 349986 687454
rect 350222 687218 350306 687454
rect 350542 687218 350574 687454
rect 349954 687134 350574 687218
rect 349954 686898 349986 687134
rect 350222 686898 350306 687134
rect 350542 686898 350574 687134
rect 349954 657000 350574 686898
rect 350874 698614 351494 710042
rect 355994 711558 356614 711590
rect 355994 711322 356026 711558
rect 356262 711322 356346 711558
rect 356582 711322 356614 711558
rect 355994 711238 356614 711322
rect 355994 711002 356026 711238
rect 356262 711002 356346 711238
rect 356582 711002 356614 711238
rect 350874 698378 350906 698614
rect 351142 698378 351226 698614
rect 351462 698378 351494 698614
rect 350874 698294 351494 698378
rect 350874 698058 350906 698294
rect 351142 698058 351226 698294
rect 351462 698058 351494 698294
rect 350874 662614 351494 698058
rect 350874 662378 350906 662614
rect 351142 662378 351226 662614
rect 351462 662378 351494 662614
rect 350874 662294 351494 662378
rect 350874 662058 350906 662294
rect 351142 662058 351226 662294
rect 351462 662058 351494 662294
rect 350874 657000 351494 662058
rect 352274 709638 352894 709670
rect 352274 709402 352306 709638
rect 352542 709402 352626 709638
rect 352862 709402 352894 709638
rect 352274 709318 352894 709402
rect 352274 709082 352306 709318
rect 352542 709082 352626 709318
rect 352862 709082 352894 709318
rect 352274 676894 352894 709082
rect 352274 676658 352306 676894
rect 352542 676658 352626 676894
rect 352862 676658 352894 676894
rect 352274 676574 352894 676658
rect 352274 676338 352306 676574
rect 352542 676338 352626 676574
rect 352862 676338 352894 676574
rect 352274 657000 352894 676338
rect 353674 706758 354294 707750
rect 353674 706522 353706 706758
rect 353942 706522 354026 706758
rect 354262 706522 354294 706758
rect 353674 706438 354294 706522
rect 353674 706202 353706 706438
rect 353942 706202 354026 706438
rect 354262 706202 354294 706438
rect 353674 691174 354294 706202
rect 353674 690938 353706 691174
rect 353942 690938 354026 691174
rect 354262 690938 354294 691174
rect 353674 690854 354294 690938
rect 353674 690618 353706 690854
rect 353942 690618 354026 690854
rect 354262 690618 354294 690854
rect 353674 657000 354294 690618
rect 355074 705798 355694 705830
rect 355074 705562 355106 705798
rect 355342 705562 355426 705798
rect 355662 705562 355694 705798
rect 355074 705478 355694 705562
rect 355074 705242 355106 705478
rect 355342 705242 355426 705478
rect 355662 705242 355694 705478
rect 355074 669454 355694 705242
rect 355074 669218 355106 669454
rect 355342 669218 355426 669454
rect 355662 669218 355694 669454
rect 355074 669134 355694 669218
rect 355074 668898 355106 669134
rect 355342 668898 355426 669134
rect 355662 668898 355694 669134
rect 355074 657000 355694 668898
rect 355994 680614 356614 711002
rect 361114 710598 361734 711590
rect 361114 710362 361146 710598
rect 361382 710362 361466 710598
rect 361702 710362 361734 710598
rect 361114 710278 361734 710362
rect 361114 710042 361146 710278
rect 361382 710042 361466 710278
rect 361702 710042 361734 710278
rect 355994 680378 356026 680614
rect 356262 680378 356346 680614
rect 356582 680378 356614 680614
rect 355994 680294 356614 680378
rect 355994 680058 356026 680294
rect 356262 680058 356346 680294
rect 356582 680058 356614 680294
rect 355994 657000 356614 680058
rect 357394 708678 358014 709670
rect 357394 708442 357426 708678
rect 357662 708442 357746 708678
rect 357982 708442 358014 708678
rect 357394 708358 358014 708442
rect 357394 708122 357426 708358
rect 357662 708122 357746 708358
rect 357982 708122 358014 708358
rect 357394 694894 358014 708122
rect 357394 694658 357426 694894
rect 357662 694658 357746 694894
rect 357982 694658 358014 694894
rect 357394 694574 358014 694658
rect 357394 694338 357426 694574
rect 357662 694338 357746 694574
rect 357982 694338 358014 694574
rect 357394 658894 358014 694338
rect 357394 658658 357426 658894
rect 357662 658658 357746 658894
rect 357982 658658 358014 658894
rect 357394 658574 358014 658658
rect 357394 658338 357426 658574
rect 357662 658338 357746 658574
rect 357982 658338 358014 658574
rect 357394 657000 358014 658338
rect 358794 707718 359414 707750
rect 358794 707482 358826 707718
rect 359062 707482 359146 707718
rect 359382 707482 359414 707718
rect 358794 707398 359414 707482
rect 358794 707162 358826 707398
rect 359062 707162 359146 707398
rect 359382 707162 359414 707398
rect 358794 673174 359414 707162
rect 358794 672938 358826 673174
rect 359062 672938 359146 673174
rect 359382 672938 359414 673174
rect 358794 672854 359414 672938
rect 358794 672618 358826 672854
rect 359062 672618 359146 672854
rect 359382 672618 359414 672854
rect 358794 657000 359414 672618
rect 360194 704838 360814 705830
rect 360194 704602 360226 704838
rect 360462 704602 360546 704838
rect 360782 704602 360814 704838
rect 360194 704518 360814 704602
rect 360194 704282 360226 704518
rect 360462 704282 360546 704518
rect 360782 704282 360814 704518
rect 360194 687454 360814 704282
rect 360194 687218 360226 687454
rect 360462 687218 360546 687454
rect 360782 687218 360814 687454
rect 360194 687134 360814 687218
rect 360194 686898 360226 687134
rect 360462 686898 360546 687134
rect 360782 686898 360814 687134
rect 360194 657000 360814 686898
rect 361114 698614 361734 710042
rect 366234 711558 366854 711590
rect 366234 711322 366266 711558
rect 366502 711322 366586 711558
rect 366822 711322 366854 711558
rect 366234 711238 366854 711322
rect 366234 711002 366266 711238
rect 366502 711002 366586 711238
rect 366822 711002 366854 711238
rect 361114 698378 361146 698614
rect 361382 698378 361466 698614
rect 361702 698378 361734 698614
rect 361114 698294 361734 698378
rect 361114 698058 361146 698294
rect 361382 698058 361466 698294
rect 361702 698058 361734 698294
rect 361114 662614 361734 698058
rect 361114 662378 361146 662614
rect 361382 662378 361466 662614
rect 361702 662378 361734 662614
rect 361114 662294 361734 662378
rect 361114 662058 361146 662294
rect 361382 662058 361466 662294
rect 361702 662058 361734 662294
rect 361114 657000 361734 662058
rect 362514 709638 363134 709670
rect 362514 709402 362546 709638
rect 362782 709402 362866 709638
rect 363102 709402 363134 709638
rect 362514 709318 363134 709402
rect 362514 709082 362546 709318
rect 362782 709082 362866 709318
rect 363102 709082 363134 709318
rect 362514 676894 363134 709082
rect 362514 676658 362546 676894
rect 362782 676658 362866 676894
rect 363102 676658 363134 676894
rect 362514 676574 363134 676658
rect 362514 676338 362546 676574
rect 362782 676338 362866 676574
rect 363102 676338 363134 676574
rect 362514 657000 363134 676338
rect 363914 706758 364534 707750
rect 363914 706522 363946 706758
rect 364182 706522 364266 706758
rect 364502 706522 364534 706758
rect 363914 706438 364534 706522
rect 363914 706202 363946 706438
rect 364182 706202 364266 706438
rect 364502 706202 364534 706438
rect 363914 691174 364534 706202
rect 363914 690938 363946 691174
rect 364182 690938 364266 691174
rect 364502 690938 364534 691174
rect 363914 690854 364534 690938
rect 363914 690618 363946 690854
rect 364182 690618 364266 690854
rect 364502 690618 364534 690854
rect 363914 657000 364534 690618
rect 365314 705798 365934 705830
rect 365314 705562 365346 705798
rect 365582 705562 365666 705798
rect 365902 705562 365934 705798
rect 365314 705478 365934 705562
rect 365314 705242 365346 705478
rect 365582 705242 365666 705478
rect 365902 705242 365934 705478
rect 365314 669454 365934 705242
rect 365314 669218 365346 669454
rect 365582 669218 365666 669454
rect 365902 669218 365934 669454
rect 365314 669134 365934 669218
rect 365314 668898 365346 669134
rect 365582 668898 365666 669134
rect 365902 668898 365934 669134
rect 365314 657000 365934 668898
rect 366234 680614 366854 711002
rect 371354 710598 371974 711590
rect 371354 710362 371386 710598
rect 371622 710362 371706 710598
rect 371942 710362 371974 710598
rect 371354 710278 371974 710362
rect 371354 710042 371386 710278
rect 371622 710042 371706 710278
rect 371942 710042 371974 710278
rect 366234 680378 366266 680614
rect 366502 680378 366586 680614
rect 366822 680378 366854 680614
rect 366234 680294 366854 680378
rect 366234 680058 366266 680294
rect 366502 680058 366586 680294
rect 366822 680058 366854 680294
rect 366234 657000 366854 680058
rect 367634 708678 368254 709670
rect 367634 708442 367666 708678
rect 367902 708442 367986 708678
rect 368222 708442 368254 708678
rect 367634 708358 368254 708442
rect 367634 708122 367666 708358
rect 367902 708122 367986 708358
rect 368222 708122 368254 708358
rect 367634 694894 368254 708122
rect 367634 694658 367666 694894
rect 367902 694658 367986 694894
rect 368222 694658 368254 694894
rect 367634 694574 368254 694658
rect 367634 694338 367666 694574
rect 367902 694338 367986 694574
rect 368222 694338 368254 694574
rect 367634 658894 368254 694338
rect 367634 658658 367666 658894
rect 367902 658658 367986 658894
rect 368222 658658 368254 658894
rect 367634 658574 368254 658658
rect 367634 658338 367666 658574
rect 367902 658338 367986 658574
rect 368222 658338 368254 658574
rect 367634 657000 368254 658338
rect 369034 707718 369654 707750
rect 369034 707482 369066 707718
rect 369302 707482 369386 707718
rect 369622 707482 369654 707718
rect 369034 707398 369654 707482
rect 369034 707162 369066 707398
rect 369302 707162 369386 707398
rect 369622 707162 369654 707398
rect 369034 673174 369654 707162
rect 369034 672938 369066 673174
rect 369302 672938 369386 673174
rect 369622 672938 369654 673174
rect 369034 672854 369654 672938
rect 369034 672618 369066 672854
rect 369302 672618 369386 672854
rect 369622 672618 369654 672854
rect 369034 657000 369654 672618
rect 370434 704838 371054 705830
rect 370434 704602 370466 704838
rect 370702 704602 370786 704838
rect 371022 704602 371054 704838
rect 370434 704518 371054 704602
rect 370434 704282 370466 704518
rect 370702 704282 370786 704518
rect 371022 704282 371054 704518
rect 370434 687454 371054 704282
rect 370434 687218 370466 687454
rect 370702 687218 370786 687454
rect 371022 687218 371054 687454
rect 370434 687134 371054 687218
rect 370434 686898 370466 687134
rect 370702 686898 370786 687134
rect 371022 686898 371054 687134
rect 370434 657000 371054 686898
rect 371354 698614 371974 710042
rect 376474 711558 377094 711590
rect 376474 711322 376506 711558
rect 376742 711322 376826 711558
rect 377062 711322 377094 711558
rect 376474 711238 377094 711322
rect 376474 711002 376506 711238
rect 376742 711002 376826 711238
rect 377062 711002 377094 711238
rect 371354 698378 371386 698614
rect 371622 698378 371706 698614
rect 371942 698378 371974 698614
rect 371354 698294 371974 698378
rect 371354 698058 371386 698294
rect 371622 698058 371706 698294
rect 371942 698058 371974 698294
rect 371354 662614 371974 698058
rect 371354 662378 371386 662614
rect 371622 662378 371706 662614
rect 371942 662378 371974 662614
rect 371354 662294 371974 662378
rect 371354 662058 371386 662294
rect 371622 662058 371706 662294
rect 371942 662058 371974 662294
rect 371354 657000 371974 662058
rect 372754 709638 373374 709670
rect 372754 709402 372786 709638
rect 373022 709402 373106 709638
rect 373342 709402 373374 709638
rect 372754 709318 373374 709402
rect 372754 709082 372786 709318
rect 373022 709082 373106 709318
rect 373342 709082 373374 709318
rect 372754 676894 373374 709082
rect 372754 676658 372786 676894
rect 373022 676658 373106 676894
rect 373342 676658 373374 676894
rect 372754 676574 373374 676658
rect 372754 676338 372786 676574
rect 373022 676338 373106 676574
rect 373342 676338 373374 676574
rect 372754 657000 373374 676338
rect 374154 706758 374774 707750
rect 374154 706522 374186 706758
rect 374422 706522 374506 706758
rect 374742 706522 374774 706758
rect 374154 706438 374774 706522
rect 374154 706202 374186 706438
rect 374422 706202 374506 706438
rect 374742 706202 374774 706438
rect 374154 691174 374774 706202
rect 374154 690938 374186 691174
rect 374422 690938 374506 691174
rect 374742 690938 374774 691174
rect 374154 690854 374774 690938
rect 374154 690618 374186 690854
rect 374422 690618 374506 690854
rect 374742 690618 374774 690854
rect 374154 657000 374774 690618
rect 375554 705798 376174 705830
rect 375554 705562 375586 705798
rect 375822 705562 375906 705798
rect 376142 705562 376174 705798
rect 375554 705478 376174 705562
rect 375554 705242 375586 705478
rect 375822 705242 375906 705478
rect 376142 705242 376174 705478
rect 375554 669454 376174 705242
rect 375554 669218 375586 669454
rect 375822 669218 375906 669454
rect 376142 669218 376174 669454
rect 375554 669134 376174 669218
rect 375554 668898 375586 669134
rect 375822 668898 375906 669134
rect 376142 668898 376174 669134
rect 375554 657000 376174 668898
rect 376474 680614 377094 711002
rect 381594 710598 382214 711590
rect 381594 710362 381626 710598
rect 381862 710362 381946 710598
rect 382182 710362 382214 710598
rect 381594 710278 382214 710362
rect 381594 710042 381626 710278
rect 381862 710042 381946 710278
rect 382182 710042 382214 710278
rect 376474 680378 376506 680614
rect 376742 680378 376826 680614
rect 377062 680378 377094 680614
rect 376474 680294 377094 680378
rect 376474 680058 376506 680294
rect 376742 680058 376826 680294
rect 377062 680058 377094 680294
rect 376474 657000 377094 680058
rect 377874 708678 378494 709670
rect 377874 708442 377906 708678
rect 378142 708442 378226 708678
rect 378462 708442 378494 708678
rect 377874 708358 378494 708442
rect 377874 708122 377906 708358
rect 378142 708122 378226 708358
rect 378462 708122 378494 708358
rect 377874 694894 378494 708122
rect 377874 694658 377906 694894
rect 378142 694658 378226 694894
rect 378462 694658 378494 694894
rect 377874 694574 378494 694658
rect 377874 694338 377906 694574
rect 378142 694338 378226 694574
rect 378462 694338 378494 694574
rect 377874 658894 378494 694338
rect 377874 658658 377906 658894
rect 378142 658658 378226 658894
rect 378462 658658 378494 658894
rect 377874 658574 378494 658658
rect 377874 658338 377906 658574
rect 378142 658338 378226 658574
rect 378462 658338 378494 658574
rect 377874 657000 378494 658338
rect 379274 707718 379894 707750
rect 379274 707482 379306 707718
rect 379542 707482 379626 707718
rect 379862 707482 379894 707718
rect 379274 707398 379894 707482
rect 379274 707162 379306 707398
rect 379542 707162 379626 707398
rect 379862 707162 379894 707398
rect 379274 673174 379894 707162
rect 379274 672938 379306 673174
rect 379542 672938 379626 673174
rect 379862 672938 379894 673174
rect 379274 672854 379894 672938
rect 379274 672618 379306 672854
rect 379542 672618 379626 672854
rect 379862 672618 379894 672854
rect 379274 657000 379894 672618
rect 380674 704838 381294 705830
rect 380674 704602 380706 704838
rect 380942 704602 381026 704838
rect 381262 704602 381294 704838
rect 380674 704518 381294 704602
rect 380674 704282 380706 704518
rect 380942 704282 381026 704518
rect 381262 704282 381294 704518
rect 380674 687454 381294 704282
rect 380674 687218 380706 687454
rect 380942 687218 381026 687454
rect 381262 687218 381294 687454
rect 380674 687134 381294 687218
rect 380674 686898 380706 687134
rect 380942 686898 381026 687134
rect 381262 686898 381294 687134
rect 380674 657000 381294 686898
rect 381594 698614 382214 710042
rect 386714 711558 387334 711590
rect 386714 711322 386746 711558
rect 386982 711322 387066 711558
rect 387302 711322 387334 711558
rect 386714 711238 387334 711322
rect 386714 711002 386746 711238
rect 386982 711002 387066 711238
rect 387302 711002 387334 711238
rect 381594 698378 381626 698614
rect 381862 698378 381946 698614
rect 382182 698378 382214 698614
rect 381594 698294 382214 698378
rect 381594 698058 381626 698294
rect 381862 698058 381946 698294
rect 382182 698058 382214 698294
rect 381594 662614 382214 698058
rect 381594 662378 381626 662614
rect 381862 662378 381946 662614
rect 382182 662378 382214 662614
rect 381594 662294 382214 662378
rect 381594 662058 381626 662294
rect 381862 662058 381946 662294
rect 382182 662058 382214 662294
rect 381594 657000 382214 662058
rect 382994 709638 383614 709670
rect 382994 709402 383026 709638
rect 383262 709402 383346 709638
rect 383582 709402 383614 709638
rect 382994 709318 383614 709402
rect 382994 709082 383026 709318
rect 383262 709082 383346 709318
rect 383582 709082 383614 709318
rect 382994 676894 383614 709082
rect 382994 676658 383026 676894
rect 383262 676658 383346 676894
rect 383582 676658 383614 676894
rect 382994 676574 383614 676658
rect 382994 676338 383026 676574
rect 383262 676338 383346 676574
rect 383582 676338 383614 676574
rect 382994 657000 383614 676338
rect 384394 706758 385014 707750
rect 384394 706522 384426 706758
rect 384662 706522 384746 706758
rect 384982 706522 385014 706758
rect 384394 706438 385014 706522
rect 384394 706202 384426 706438
rect 384662 706202 384746 706438
rect 384982 706202 385014 706438
rect 384394 691174 385014 706202
rect 384394 690938 384426 691174
rect 384662 690938 384746 691174
rect 384982 690938 385014 691174
rect 384394 690854 385014 690938
rect 384394 690618 384426 690854
rect 384662 690618 384746 690854
rect 384982 690618 385014 690854
rect 384394 657000 385014 690618
rect 385794 705798 386414 705830
rect 385794 705562 385826 705798
rect 386062 705562 386146 705798
rect 386382 705562 386414 705798
rect 385794 705478 386414 705562
rect 385794 705242 385826 705478
rect 386062 705242 386146 705478
rect 386382 705242 386414 705478
rect 385794 669454 386414 705242
rect 385794 669218 385826 669454
rect 386062 669218 386146 669454
rect 386382 669218 386414 669454
rect 385794 669134 386414 669218
rect 385794 668898 385826 669134
rect 386062 668898 386146 669134
rect 386382 668898 386414 669134
rect 385794 657000 386414 668898
rect 386714 680614 387334 711002
rect 391834 710598 392454 711590
rect 391834 710362 391866 710598
rect 392102 710362 392186 710598
rect 392422 710362 392454 710598
rect 391834 710278 392454 710362
rect 391834 710042 391866 710278
rect 392102 710042 392186 710278
rect 392422 710042 392454 710278
rect 386714 680378 386746 680614
rect 386982 680378 387066 680614
rect 387302 680378 387334 680614
rect 386714 680294 387334 680378
rect 386714 680058 386746 680294
rect 386982 680058 387066 680294
rect 387302 680058 387334 680294
rect 386714 657000 387334 680058
rect 388114 708678 388734 709670
rect 388114 708442 388146 708678
rect 388382 708442 388466 708678
rect 388702 708442 388734 708678
rect 388114 708358 388734 708442
rect 388114 708122 388146 708358
rect 388382 708122 388466 708358
rect 388702 708122 388734 708358
rect 388114 694894 388734 708122
rect 388114 694658 388146 694894
rect 388382 694658 388466 694894
rect 388702 694658 388734 694894
rect 388114 694574 388734 694658
rect 388114 694338 388146 694574
rect 388382 694338 388466 694574
rect 388702 694338 388734 694574
rect 388114 658894 388734 694338
rect 388114 658658 388146 658894
rect 388382 658658 388466 658894
rect 388702 658658 388734 658894
rect 388114 658574 388734 658658
rect 388114 658338 388146 658574
rect 388382 658338 388466 658574
rect 388702 658338 388734 658574
rect 388114 657000 388734 658338
rect 389514 707718 390134 707750
rect 389514 707482 389546 707718
rect 389782 707482 389866 707718
rect 390102 707482 390134 707718
rect 389514 707398 390134 707482
rect 389514 707162 389546 707398
rect 389782 707162 389866 707398
rect 390102 707162 390134 707398
rect 389514 673174 390134 707162
rect 389514 672938 389546 673174
rect 389782 672938 389866 673174
rect 390102 672938 390134 673174
rect 389514 672854 390134 672938
rect 389514 672618 389546 672854
rect 389782 672618 389866 672854
rect 390102 672618 390134 672854
rect 389514 657000 390134 672618
rect 390914 704838 391534 705830
rect 390914 704602 390946 704838
rect 391182 704602 391266 704838
rect 391502 704602 391534 704838
rect 390914 704518 391534 704602
rect 390914 704282 390946 704518
rect 391182 704282 391266 704518
rect 391502 704282 391534 704518
rect 390914 687454 391534 704282
rect 390914 687218 390946 687454
rect 391182 687218 391266 687454
rect 391502 687218 391534 687454
rect 390914 687134 391534 687218
rect 390914 686898 390946 687134
rect 391182 686898 391266 687134
rect 391502 686898 391534 687134
rect 390914 657000 391534 686898
rect 391834 698614 392454 710042
rect 396954 711558 397574 711590
rect 396954 711322 396986 711558
rect 397222 711322 397306 711558
rect 397542 711322 397574 711558
rect 396954 711238 397574 711322
rect 396954 711002 396986 711238
rect 397222 711002 397306 711238
rect 397542 711002 397574 711238
rect 391834 698378 391866 698614
rect 392102 698378 392186 698614
rect 392422 698378 392454 698614
rect 391834 698294 392454 698378
rect 391834 698058 391866 698294
rect 392102 698058 392186 698294
rect 392422 698058 392454 698294
rect 391834 662614 392454 698058
rect 391834 662378 391866 662614
rect 392102 662378 392186 662614
rect 392422 662378 392454 662614
rect 391834 662294 392454 662378
rect 391834 662058 391866 662294
rect 392102 662058 392186 662294
rect 392422 662058 392454 662294
rect 391834 657000 392454 662058
rect 393234 709638 393854 709670
rect 393234 709402 393266 709638
rect 393502 709402 393586 709638
rect 393822 709402 393854 709638
rect 393234 709318 393854 709402
rect 393234 709082 393266 709318
rect 393502 709082 393586 709318
rect 393822 709082 393854 709318
rect 393234 676894 393854 709082
rect 393234 676658 393266 676894
rect 393502 676658 393586 676894
rect 393822 676658 393854 676894
rect 393234 676574 393854 676658
rect 393234 676338 393266 676574
rect 393502 676338 393586 676574
rect 393822 676338 393854 676574
rect 393234 657000 393854 676338
rect 394634 706758 395254 707750
rect 394634 706522 394666 706758
rect 394902 706522 394986 706758
rect 395222 706522 395254 706758
rect 394634 706438 395254 706522
rect 394634 706202 394666 706438
rect 394902 706202 394986 706438
rect 395222 706202 395254 706438
rect 394634 691174 395254 706202
rect 394634 690938 394666 691174
rect 394902 690938 394986 691174
rect 395222 690938 395254 691174
rect 394634 690854 395254 690938
rect 394634 690618 394666 690854
rect 394902 690618 394986 690854
rect 395222 690618 395254 690854
rect 394634 657000 395254 690618
rect 396034 705798 396654 705830
rect 396034 705562 396066 705798
rect 396302 705562 396386 705798
rect 396622 705562 396654 705798
rect 396034 705478 396654 705562
rect 396034 705242 396066 705478
rect 396302 705242 396386 705478
rect 396622 705242 396654 705478
rect 396034 669454 396654 705242
rect 396034 669218 396066 669454
rect 396302 669218 396386 669454
rect 396622 669218 396654 669454
rect 396034 669134 396654 669218
rect 396034 668898 396066 669134
rect 396302 668898 396386 669134
rect 396622 668898 396654 669134
rect 396034 657000 396654 668898
rect 396954 680614 397574 711002
rect 402074 710598 402694 711590
rect 402074 710362 402106 710598
rect 402342 710362 402426 710598
rect 402662 710362 402694 710598
rect 402074 710278 402694 710362
rect 402074 710042 402106 710278
rect 402342 710042 402426 710278
rect 402662 710042 402694 710278
rect 396954 680378 396986 680614
rect 397222 680378 397306 680614
rect 397542 680378 397574 680614
rect 396954 680294 397574 680378
rect 396954 680058 396986 680294
rect 397222 680058 397306 680294
rect 397542 680058 397574 680294
rect 396954 657000 397574 680058
rect 398354 708678 398974 709670
rect 398354 708442 398386 708678
rect 398622 708442 398706 708678
rect 398942 708442 398974 708678
rect 398354 708358 398974 708442
rect 398354 708122 398386 708358
rect 398622 708122 398706 708358
rect 398942 708122 398974 708358
rect 398354 694894 398974 708122
rect 398354 694658 398386 694894
rect 398622 694658 398706 694894
rect 398942 694658 398974 694894
rect 398354 694574 398974 694658
rect 398354 694338 398386 694574
rect 398622 694338 398706 694574
rect 398942 694338 398974 694574
rect 398354 658894 398974 694338
rect 398354 658658 398386 658894
rect 398622 658658 398706 658894
rect 398942 658658 398974 658894
rect 398354 658574 398974 658658
rect 398354 658338 398386 658574
rect 398622 658338 398706 658574
rect 398942 658338 398974 658574
rect 398354 657000 398974 658338
rect 399754 707718 400374 707750
rect 399754 707482 399786 707718
rect 400022 707482 400106 707718
rect 400342 707482 400374 707718
rect 399754 707398 400374 707482
rect 399754 707162 399786 707398
rect 400022 707162 400106 707398
rect 400342 707162 400374 707398
rect 399754 673174 400374 707162
rect 399754 672938 399786 673174
rect 400022 672938 400106 673174
rect 400342 672938 400374 673174
rect 399754 672854 400374 672938
rect 399754 672618 399786 672854
rect 400022 672618 400106 672854
rect 400342 672618 400374 672854
rect 399754 657000 400374 672618
rect 401154 704838 401774 705830
rect 401154 704602 401186 704838
rect 401422 704602 401506 704838
rect 401742 704602 401774 704838
rect 401154 704518 401774 704602
rect 401154 704282 401186 704518
rect 401422 704282 401506 704518
rect 401742 704282 401774 704518
rect 401154 687454 401774 704282
rect 401154 687218 401186 687454
rect 401422 687218 401506 687454
rect 401742 687218 401774 687454
rect 401154 687134 401774 687218
rect 401154 686898 401186 687134
rect 401422 686898 401506 687134
rect 401742 686898 401774 687134
rect 401154 657000 401774 686898
rect 402074 698614 402694 710042
rect 407194 711558 407814 711590
rect 407194 711322 407226 711558
rect 407462 711322 407546 711558
rect 407782 711322 407814 711558
rect 407194 711238 407814 711322
rect 407194 711002 407226 711238
rect 407462 711002 407546 711238
rect 407782 711002 407814 711238
rect 402074 698378 402106 698614
rect 402342 698378 402426 698614
rect 402662 698378 402694 698614
rect 402074 698294 402694 698378
rect 402074 698058 402106 698294
rect 402342 698058 402426 698294
rect 402662 698058 402694 698294
rect 402074 662614 402694 698058
rect 402074 662378 402106 662614
rect 402342 662378 402426 662614
rect 402662 662378 402694 662614
rect 402074 662294 402694 662378
rect 402074 662058 402106 662294
rect 402342 662058 402426 662294
rect 402662 662058 402694 662294
rect 402074 657000 402694 662058
rect 403474 709638 404094 709670
rect 403474 709402 403506 709638
rect 403742 709402 403826 709638
rect 404062 709402 404094 709638
rect 403474 709318 404094 709402
rect 403474 709082 403506 709318
rect 403742 709082 403826 709318
rect 404062 709082 404094 709318
rect 403474 676894 404094 709082
rect 403474 676658 403506 676894
rect 403742 676658 403826 676894
rect 404062 676658 404094 676894
rect 403474 676574 404094 676658
rect 403474 676338 403506 676574
rect 403742 676338 403826 676574
rect 404062 676338 404094 676574
rect 403474 657000 404094 676338
rect 404874 706758 405494 707750
rect 404874 706522 404906 706758
rect 405142 706522 405226 706758
rect 405462 706522 405494 706758
rect 404874 706438 405494 706522
rect 404874 706202 404906 706438
rect 405142 706202 405226 706438
rect 405462 706202 405494 706438
rect 404874 691174 405494 706202
rect 404874 690938 404906 691174
rect 405142 690938 405226 691174
rect 405462 690938 405494 691174
rect 404874 690854 405494 690938
rect 404874 690618 404906 690854
rect 405142 690618 405226 690854
rect 405462 690618 405494 690854
rect 404874 657000 405494 690618
rect 406274 705798 406894 705830
rect 406274 705562 406306 705798
rect 406542 705562 406626 705798
rect 406862 705562 406894 705798
rect 406274 705478 406894 705562
rect 406274 705242 406306 705478
rect 406542 705242 406626 705478
rect 406862 705242 406894 705478
rect 406274 669454 406894 705242
rect 406274 669218 406306 669454
rect 406542 669218 406626 669454
rect 406862 669218 406894 669454
rect 406274 669134 406894 669218
rect 406274 668898 406306 669134
rect 406542 668898 406626 669134
rect 406862 668898 406894 669134
rect 406274 657000 406894 668898
rect 407194 680614 407814 711002
rect 412314 710598 412934 711590
rect 412314 710362 412346 710598
rect 412582 710362 412666 710598
rect 412902 710362 412934 710598
rect 412314 710278 412934 710362
rect 412314 710042 412346 710278
rect 412582 710042 412666 710278
rect 412902 710042 412934 710278
rect 407194 680378 407226 680614
rect 407462 680378 407546 680614
rect 407782 680378 407814 680614
rect 407194 680294 407814 680378
rect 407194 680058 407226 680294
rect 407462 680058 407546 680294
rect 407782 680058 407814 680294
rect 407194 657000 407814 680058
rect 408594 708678 409214 709670
rect 408594 708442 408626 708678
rect 408862 708442 408946 708678
rect 409182 708442 409214 708678
rect 408594 708358 409214 708442
rect 408594 708122 408626 708358
rect 408862 708122 408946 708358
rect 409182 708122 409214 708358
rect 408594 694894 409214 708122
rect 408594 694658 408626 694894
rect 408862 694658 408946 694894
rect 409182 694658 409214 694894
rect 408594 694574 409214 694658
rect 408594 694338 408626 694574
rect 408862 694338 408946 694574
rect 409182 694338 409214 694574
rect 408594 658894 409214 694338
rect 408594 658658 408626 658894
rect 408862 658658 408946 658894
rect 409182 658658 409214 658894
rect 408594 658574 409214 658658
rect 408594 658338 408626 658574
rect 408862 658338 408946 658574
rect 409182 658338 409214 658574
rect 408594 657000 409214 658338
rect 409994 707718 410614 707750
rect 409994 707482 410026 707718
rect 410262 707482 410346 707718
rect 410582 707482 410614 707718
rect 409994 707398 410614 707482
rect 409994 707162 410026 707398
rect 410262 707162 410346 707398
rect 410582 707162 410614 707398
rect 409994 673174 410614 707162
rect 409994 672938 410026 673174
rect 410262 672938 410346 673174
rect 410582 672938 410614 673174
rect 409994 672854 410614 672938
rect 409994 672618 410026 672854
rect 410262 672618 410346 672854
rect 410582 672618 410614 672854
rect 409994 657000 410614 672618
rect 411394 704838 412014 705830
rect 411394 704602 411426 704838
rect 411662 704602 411746 704838
rect 411982 704602 412014 704838
rect 411394 704518 412014 704602
rect 411394 704282 411426 704518
rect 411662 704282 411746 704518
rect 411982 704282 412014 704518
rect 411394 687454 412014 704282
rect 411394 687218 411426 687454
rect 411662 687218 411746 687454
rect 411982 687218 412014 687454
rect 411394 687134 412014 687218
rect 411394 686898 411426 687134
rect 411662 686898 411746 687134
rect 411982 686898 412014 687134
rect 411394 657000 412014 686898
rect 412314 698614 412934 710042
rect 417434 711558 418054 711590
rect 417434 711322 417466 711558
rect 417702 711322 417786 711558
rect 418022 711322 418054 711558
rect 417434 711238 418054 711322
rect 417434 711002 417466 711238
rect 417702 711002 417786 711238
rect 418022 711002 418054 711238
rect 412314 698378 412346 698614
rect 412582 698378 412666 698614
rect 412902 698378 412934 698614
rect 412314 698294 412934 698378
rect 412314 698058 412346 698294
rect 412582 698058 412666 698294
rect 412902 698058 412934 698294
rect 412314 662614 412934 698058
rect 412314 662378 412346 662614
rect 412582 662378 412666 662614
rect 412902 662378 412934 662614
rect 412314 662294 412934 662378
rect 412314 662058 412346 662294
rect 412582 662058 412666 662294
rect 412902 662058 412934 662294
rect 412314 657000 412934 662058
rect 413714 709638 414334 709670
rect 413714 709402 413746 709638
rect 413982 709402 414066 709638
rect 414302 709402 414334 709638
rect 413714 709318 414334 709402
rect 413714 709082 413746 709318
rect 413982 709082 414066 709318
rect 414302 709082 414334 709318
rect 413714 676894 414334 709082
rect 413714 676658 413746 676894
rect 413982 676658 414066 676894
rect 414302 676658 414334 676894
rect 413714 676574 414334 676658
rect 413714 676338 413746 676574
rect 413982 676338 414066 676574
rect 414302 676338 414334 676574
rect 413714 657000 414334 676338
rect 415114 706758 415734 707750
rect 415114 706522 415146 706758
rect 415382 706522 415466 706758
rect 415702 706522 415734 706758
rect 415114 706438 415734 706522
rect 415114 706202 415146 706438
rect 415382 706202 415466 706438
rect 415702 706202 415734 706438
rect 415114 691174 415734 706202
rect 415114 690938 415146 691174
rect 415382 690938 415466 691174
rect 415702 690938 415734 691174
rect 415114 690854 415734 690938
rect 415114 690618 415146 690854
rect 415382 690618 415466 690854
rect 415702 690618 415734 690854
rect 415114 657000 415734 690618
rect 416514 705798 417134 705830
rect 416514 705562 416546 705798
rect 416782 705562 416866 705798
rect 417102 705562 417134 705798
rect 416514 705478 417134 705562
rect 416514 705242 416546 705478
rect 416782 705242 416866 705478
rect 417102 705242 417134 705478
rect 416514 669454 417134 705242
rect 416514 669218 416546 669454
rect 416782 669218 416866 669454
rect 417102 669218 417134 669454
rect 416514 669134 417134 669218
rect 416514 668898 416546 669134
rect 416782 668898 416866 669134
rect 417102 668898 417134 669134
rect 416514 657000 417134 668898
rect 417434 680614 418054 711002
rect 422554 710598 423174 711590
rect 422554 710362 422586 710598
rect 422822 710362 422906 710598
rect 423142 710362 423174 710598
rect 422554 710278 423174 710362
rect 422554 710042 422586 710278
rect 422822 710042 422906 710278
rect 423142 710042 423174 710278
rect 417434 680378 417466 680614
rect 417702 680378 417786 680614
rect 418022 680378 418054 680614
rect 417434 680294 418054 680378
rect 417434 680058 417466 680294
rect 417702 680058 417786 680294
rect 418022 680058 418054 680294
rect 417434 657000 418054 680058
rect 418834 708678 419454 709670
rect 418834 708442 418866 708678
rect 419102 708442 419186 708678
rect 419422 708442 419454 708678
rect 418834 708358 419454 708442
rect 418834 708122 418866 708358
rect 419102 708122 419186 708358
rect 419422 708122 419454 708358
rect 418834 694894 419454 708122
rect 418834 694658 418866 694894
rect 419102 694658 419186 694894
rect 419422 694658 419454 694894
rect 418834 694574 419454 694658
rect 418834 694338 418866 694574
rect 419102 694338 419186 694574
rect 419422 694338 419454 694574
rect 418834 658894 419454 694338
rect 418834 658658 418866 658894
rect 419102 658658 419186 658894
rect 419422 658658 419454 658894
rect 418834 658574 419454 658658
rect 418834 658338 418866 658574
rect 419102 658338 419186 658574
rect 419422 658338 419454 658574
rect 418834 657000 419454 658338
rect 420234 707718 420854 707750
rect 420234 707482 420266 707718
rect 420502 707482 420586 707718
rect 420822 707482 420854 707718
rect 420234 707398 420854 707482
rect 420234 707162 420266 707398
rect 420502 707162 420586 707398
rect 420822 707162 420854 707398
rect 420234 673174 420854 707162
rect 420234 672938 420266 673174
rect 420502 672938 420586 673174
rect 420822 672938 420854 673174
rect 420234 672854 420854 672938
rect 420234 672618 420266 672854
rect 420502 672618 420586 672854
rect 420822 672618 420854 672854
rect 420234 657000 420854 672618
rect 421634 704838 422254 705830
rect 421634 704602 421666 704838
rect 421902 704602 421986 704838
rect 422222 704602 422254 704838
rect 421634 704518 422254 704602
rect 421634 704282 421666 704518
rect 421902 704282 421986 704518
rect 422222 704282 422254 704518
rect 421634 687454 422254 704282
rect 421634 687218 421666 687454
rect 421902 687218 421986 687454
rect 422222 687218 422254 687454
rect 421634 687134 422254 687218
rect 421634 686898 421666 687134
rect 421902 686898 421986 687134
rect 422222 686898 422254 687134
rect 421634 657000 422254 686898
rect 422554 698614 423174 710042
rect 427674 711558 428294 711590
rect 427674 711322 427706 711558
rect 427942 711322 428026 711558
rect 428262 711322 428294 711558
rect 427674 711238 428294 711322
rect 427674 711002 427706 711238
rect 427942 711002 428026 711238
rect 428262 711002 428294 711238
rect 422554 698378 422586 698614
rect 422822 698378 422906 698614
rect 423142 698378 423174 698614
rect 422554 698294 423174 698378
rect 422554 698058 422586 698294
rect 422822 698058 422906 698294
rect 423142 698058 423174 698294
rect 422554 662614 423174 698058
rect 422554 662378 422586 662614
rect 422822 662378 422906 662614
rect 423142 662378 423174 662614
rect 422554 662294 423174 662378
rect 422554 662058 422586 662294
rect 422822 662058 422906 662294
rect 423142 662058 423174 662294
rect 422554 657000 423174 662058
rect 423954 709638 424574 709670
rect 423954 709402 423986 709638
rect 424222 709402 424306 709638
rect 424542 709402 424574 709638
rect 423954 709318 424574 709402
rect 423954 709082 423986 709318
rect 424222 709082 424306 709318
rect 424542 709082 424574 709318
rect 423954 676894 424574 709082
rect 423954 676658 423986 676894
rect 424222 676658 424306 676894
rect 424542 676658 424574 676894
rect 423954 676574 424574 676658
rect 423954 676338 423986 676574
rect 424222 676338 424306 676574
rect 424542 676338 424574 676574
rect 423954 657000 424574 676338
rect 425354 706758 425974 707750
rect 425354 706522 425386 706758
rect 425622 706522 425706 706758
rect 425942 706522 425974 706758
rect 425354 706438 425974 706522
rect 425354 706202 425386 706438
rect 425622 706202 425706 706438
rect 425942 706202 425974 706438
rect 425354 691174 425974 706202
rect 425354 690938 425386 691174
rect 425622 690938 425706 691174
rect 425942 690938 425974 691174
rect 425354 690854 425974 690938
rect 425354 690618 425386 690854
rect 425622 690618 425706 690854
rect 425942 690618 425974 690854
rect 425354 657000 425974 690618
rect 426754 705798 427374 705830
rect 426754 705562 426786 705798
rect 427022 705562 427106 705798
rect 427342 705562 427374 705798
rect 426754 705478 427374 705562
rect 426754 705242 426786 705478
rect 427022 705242 427106 705478
rect 427342 705242 427374 705478
rect 426754 669454 427374 705242
rect 426754 669218 426786 669454
rect 427022 669218 427106 669454
rect 427342 669218 427374 669454
rect 426754 669134 427374 669218
rect 426754 668898 426786 669134
rect 427022 668898 427106 669134
rect 427342 668898 427374 669134
rect 426754 657000 427374 668898
rect 427674 680614 428294 711002
rect 432794 710598 433414 711590
rect 432794 710362 432826 710598
rect 433062 710362 433146 710598
rect 433382 710362 433414 710598
rect 432794 710278 433414 710362
rect 432794 710042 432826 710278
rect 433062 710042 433146 710278
rect 433382 710042 433414 710278
rect 427674 680378 427706 680614
rect 427942 680378 428026 680614
rect 428262 680378 428294 680614
rect 427674 680294 428294 680378
rect 427674 680058 427706 680294
rect 427942 680058 428026 680294
rect 428262 680058 428294 680294
rect 427674 657000 428294 680058
rect 429074 708678 429694 709670
rect 429074 708442 429106 708678
rect 429342 708442 429426 708678
rect 429662 708442 429694 708678
rect 429074 708358 429694 708442
rect 429074 708122 429106 708358
rect 429342 708122 429426 708358
rect 429662 708122 429694 708358
rect 429074 694894 429694 708122
rect 429074 694658 429106 694894
rect 429342 694658 429426 694894
rect 429662 694658 429694 694894
rect 429074 694574 429694 694658
rect 429074 694338 429106 694574
rect 429342 694338 429426 694574
rect 429662 694338 429694 694574
rect 429074 658894 429694 694338
rect 429074 658658 429106 658894
rect 429342 658658 429426 658894
rect 429662 658658 429694 658894
rect 429074 658574 429694 658658
rect 429074 658338 429106 658574
rect 429342 658338 429426 658574
rect 429662 658338 429694 658574
rect 429074 657000 429694 658338
rect 430474 707718 431094 707750
rect 430474 707482 430506 707718
rect 430742 707482 430826 707718
rect 431062 707482 431094 707718
rect 430474 707398 431094 707482
rect 430474 707162 430506 707398
rect 430742 707162 430826 707398
rect 431062 707162 431094 707398
rect 430474 673174 431094 707162
rect 430474 672938 430506 673174
rect 430742 672938 430826 673174
rect 431062 672938 431094 673174
rect 430474 672854 431094 672938
rect 430474 672618 430506 672854
rect 430742 672618 430826 672854
rect 431062 672618 431094 672854
rect 430474 657000 431094 672618
rect 431874 704838 432494 705830
rect 431874 704602 431906 704838
rect 432142 704602 432226 704838
rect 432462 704602 432494 704838
rect 431874 704518 432494 704602
rect 431874 704282 431906 704518
rect 432142 704282 432226 704518
rect 432462 704282 432494 704518
rect 431874 687454 432494 704282
rect 431874 687218 431906 687454
rect 432142 687218 432226 687454
rect 432462 687218 432494 687454
rect 431874 687134 432494 687218
rect 431874 686898 431906 687134
rect 432142 686898 432226 687134
rect 432462 686898 432494 687134
rect 431874 657000 432494 686898
rect 432794 698614 433414 710042
rect 437914 711558 438534 711590
rect 437914 711322 437946 711558
rect 438182 711322 438266 711558
rect 438502 711322 438534 711558
rect 437914 711238 438534 711322
rect 437914 711002 437946 711238
rect 438182 711002 438266 711238
rect 438502 711002 438534 711238
rect 432794 698378 432826 698614
rect 433062 698378 433146 698614
rect 433382 698378 433414 698614
rect 432794 698294 433414 698378
rect 432794 698058 432826 698294
rect 433062 698058 433146 698294
rect 433382 698058 433414 698294
rect 432794 662614 433414 698058
rect 432794 662378 432826 662614
rect 433062 662378 433146 662614
rect 433382 662378 433414 662614
rect 432794 662294 433414 662378
rect 432794 662058 432826 662294
rect 433062 662058 433146 662294
rect 433382 662058 433414 662294
rect 432794 657000 433414 662058
rect 434194 709638 434814 709670
rect 434194 709402 434226 709638
rect 434462 709402 434546 709638
rect 434782 709402 434814 709638
rect 434194 709318 434814 709402
rect 434194 709082 434226 709318
rect 434462 709082 434546 709318
rect 434782 709082 434814 709318
rect 434194 676894 434814 709082
rect 434194 676658 434226 676894
rect 434462 676658 434546 676894
rect 434782 676658 434814 676894
rect 434194 676574 434814 676658
rect 434194 676338 434226 676574
rect 434462 676338 434546 676574
rect 434782 676338 434814 676574
rect 434194 657000 434814 676338
rect 435594 706758 436214 707750
rect 435594 706522 435626 706758
rect 435862 706522 435946 706758
rect 436182 706522 436214 706758
rect 435594 706438 436214 706522
rect 435594 706202 435626 706438
rect 435862 706202 435946 706438
rect 436182 706202 436214 706438
rect 435594 691174 436214 706202
rect 435594 690938 435626 691174
rect 435862 690938 435946 691174
rect 436182 690938 436214 691174
rect 435594 690854 436214 690938
rect 435594 690618 435626 690854
rect 435862 690618 435946 690854
rect 436182 690618 436214 690854
rect 435594 657000 436214 690618
rect 436994 705798 437614 705830
rect 436994 705562 437026 705798
rect 437262 705562 437346 705798
rect 437582 705562 437614 705798
rect 436994 705478 437614 705562
rect 436994 705242 437026 705478
rect 437262 705242 437346 705478
rect 437582 705242 437614 705478
rect 436994 669454 437614 705242
rect 436994 669218 437026 669454
rect 437262 669218 437346 669454
rect 437582 669218 437614 669454
rect 436994 669134 437614 669218
rect 436994 668898 437026 669134
rect 437262 668898 437346 669134
rect 437582 668898 437614 669134
rect 436994 657000 437614 668898
rect 437914 680614 438534 711002
rect 443034 710598 443654 711590
rect 443034 710362 443066 710598
rect 443302 710362 443386 710598
rect 443622 710362 443654 710598
rect 443034 710278 443654 710362
rect 443034 710042 443066 710278
rect 443302 710042 443386 710278
rect 443622 710042 443654 710278
rect 437914 680378 437946 680614
rect 438182 680378 438266 680614
rect 438502 680378 438534 680614
rect 437914 680294 438534 680378
rect 437914 680058 437946 680294
rect 438182 680058 438266 680294
rect 438502 680058 438534 680294
rect 437914 657000 438534 680058
rect 439314 708678 439934 709670
rect 439314 708442 439346 708678
rect 439582 708442 439666 708678
rect 439902 708442 439934 708678
rect 439314 708358 439934 708442
rect 439314 708122 439346 708358
rect 439582 708122 439666 708358
rect 439902 708122 439934 708358
rect 439314 694894 439934 708122
rect 439314 694658 439346 694894
rect 439582 694658 439666 694894
rect 439902 694658 439934 694894
rect 439314 694574 439934 694658
rect 439314 694338 439346 694574
rect 439582 694338 439666 694574
rect 439902 694338 439934 694574
rect 439314 658894 439934 694338
rect 439314 658658 439346 658894
rect 439582 658658 439666 658894
rect 439902 658658 439934 658894
rect 439314 658574 439934 658658
rect 439314 658338 439346 658574
rect 439582 658338 439666 658574
rect 439902 658338 439934 658574
rect 439314 657000 439934 658338
rect 440714 707718 441334 707750
rect 440714 707482 440746 707718
rect 440982 707482 441066 707718
rect 441302 707482 441334 707718
rect 440714 707398 441334 707482
rect 440714 707162 440746 707398
rect 440982 707162 441066 707398
rect 441302 707162 441334 707398
rect 440714 673174 441334 707162
rect 440714 672938 440746 673174
rect 440982 672938 441066 673174
rect 441302 672938 441334 673174
rect 440714 672854 441334 672938
rect 440714 672618 440746 672854
rect 440982 672618 441066 672854
rect 441302 672618 441334 672854
rect 440714 657000 441334 672618
rect 442114 704838 442734 705830
rect 442114 704602 442146 704838
rect 442382 704602 442466 704838
rect 442702 704602 442734 704838
rect 442114 704518 442734 704602
rect 442114 704282 442146 704518
rect 442382 704282 442466 704518
rect 442702 704282 442734 704518
rect 442114 687454 442734 704282
rect 442114 687218 442146 687454
rect 442382 687218 442466 687454
rect 442702 687218 442734 687454
rect 442114 687134 442734 687218
rect 442114 686898 442146 687134
rect 442382 686898 442466 687134
rect 442702 686898 442734 687134
rect 442114 657000 442734 686898
rect 443034 698614 443654 710042
rect 448154 711558 448774 711590
rect 448154 711322 448186 711558
rect 448422 711322 448506 711558
rect 448742 711322 448774 711558
rect 448154 711238 448774 711322
rect 448154 711002 448186 711238
rect 448422 711002 448506 711238
rect 448742 711002 448774 711238
rect 443034 698378 443066 698614
rect 443302 698378 443386 698614
rect 443622 698378 443654 698614
rect 443034 698294 443654 698378
rect 443034 698058 443066 698294
rect 443302 698058 443386 698294
rect 443622 698058 443654 698294
rect 443034 662614 443654 698058
rect 443034 662378 443066 662614
rect 443302 662378 443386 662614
rect 443622 662378 443654 662614
rect 443034 662294 443654 662378
rect 443034 662058 443066 662294
rect 443302 662058 443386 662294
rect 443622 662058 443654 662294
rect 443034 657000 443654 662058
rect 444434 709638 445054 709670
rect 444434 709402 444466 709638
rect 444702 709402 444786 709638
rect 445022 709402 445054 709638
rect 444434 709318 445054 709402
rect 444434 709082 444466 709318
rect 444702 709082 444786 709318
rect 445022 709082 445054 709318
rect 444434 676894 445054 709082
rect 444434 676658 444466 676894
rect 444702 676658 444786 676894
rect 445022 676658 445054 676894
rect 444434 676574 445054 676658
rect 444434 676338 444466 676574
rect 444702 676338 444786 676574
rect 445022 676338 445054 676574
rect 444434 657000 445054 676338
rect 445834 706758 446454 707750
rect 445834 706522 445866 706758
rect 446102 706522 446186 706758
rect 446422 706522 446454 706758
rect 445834 706438 446454 706522
rect 445834 706202 445866 706438
rect 446102 706202 446186 706438
rect 446422 706202 446454 706438
rect 445834 691174 446454 706202
rect 445834 690938 445866 691174
rect 446102 690938 446186 691174
rect 446422 690938 446454 691174
rect 445834 690854 446454 690938
rect 445834 690618 445866 690854
rect 446102 690618 446186 690854
rect 446422 690618 446454 690854
rect 445834 657000 446454 690618
rect 447234 705798 447854 705830
rect 447234 705562 447266 705798
rect 447502 705562 447586 705798
rect 447822 705562 447854 705798
rect 447234 705478 447854 705562
rect 447234 705242 447266 705478
rect 447502 705242 447586 705478
rect 447822 705242 447854 705478
rect 447234 669454 447854 705242
rect 447234 669218 447266 669454
rect 447502 669218 447586 669454
rect 447822 669218 447854 669454
rect 447234 669134 447854 669218
rect 447234 668898 447266 669134
rect 447502 668898 447586 669134
rect 447822 668898 447854 669134
rect 447234 657000 447854 668898
rect 448154 680614 448774 711002
rect 453274 710598 453894 711590
rect 453274 710362 453306 710598
rect 453542 710362 453626 710598
rect 453862 710362 453894 710598
rect 453274 710278 453894 710362
rect 453274 710042 453306 710278
rect 453542 710042 453626 710278
rect 453862 710042 453894 710278
rect 448154 680378 448186 680614
rect 448422 680378 448506 680614
rect 448742 680378 448774 680614
rect 448154 680294 448774 680378
rect 448154 680058 448186 680294
rect 448422 680058 448506 680294
rect 448742 680058 448774 680294
rect 448154 657000 448774 680058
rect 449554 708678 450174 709670
rect 449554 708442 449586 708678
rect 449822 708442 449906 708678
rect 450142 708442 450174 708678
rect 449554 708358 450174 708442
rect 449554 708122 449586 708358
rect 449822 708122 449906 708358
rect 450142 708122 450174 708358
rect 449554 694894 450174 708122
rect 449554 694658 449586 694894
rect 449822 694658 449906 694894
rect 450142 694658 450174 694894
rect 449554 694574 450174 694658
rect 449554 694338 449586 694574
rect 449822 694338 449906 694574
rect 450142 694338 450174 694574
rect 449554 658894 450174 694338
rect 449554 658658 449586 658894
rect 449822 658658 449906 658894
rect 450142 658658 450174 658894
rect 449554 658574 450174 658658
rect 449554 658338 449586 658574
rect 449822 658338 449906 658574
rect 450142 658338 450174 658574
rect 449554 657000 450174 658338
rect 450954 707718 451574 707750
rect 450954 707482 450986 707718
rect 451222 707482 451306 707718
rect 451542 707482 451574 707718
rect 450954 707398 451574 707482
rect 450954 707162 450986 707398
rect 451222 707162 451306 707398
rect 451542 707162 451574 707398
rect 450954 673174 451574 707162
rect 450954 672938 450986 673174
rect 451222 672938 451306 673174
rect 451542 672938 451574 673174
rect 450954 672854 451574 672938
rect 450954 672618 450986 672854
rect 451222 672618 451306 672854
rect 451542 672618 451574 672854
rect 450954 657000 451574 672618
rect 452354 704838 452974 705830
rect 452354 704602 452386 704838
rect 452622 704602 452706 704838
rect 452942 704602 452974 704838
rect 452354 704518 452974 704602
rect 452354 704282 452386 704518
rect 452622 704282 452706 704518
rect 452942 704282 452974 704518
rect 452354 687454 452974 704282
rect 452354 687218 452386 687454
rect 452622 687218 452706 687454
rect 452942 687218 452974 687454
rect 452354 687134 452974 687218
rect 452354 686898 452386 687134
rect 452622 686898 452706 687134
rect 452942 686898 452974 687134
rect 452354 657000 452974 686898
rect 453274 698614 453894 710042
rect 458394 711558 459014 711590
rect 458394 711322 458426 711558
rect 458662 711322 458746 711558
rect 458982 711322 459014 711558
rect 458394 711238 459014 711322
rect 458394 711002 458426 711238
rect 458662 711002 458746 711238
rect 458982 711002 459014 711238
rect 453274 698378 453306 698614
rect 453542 698378 453626 698614
rect 453862 698378 453894 698614
rect 453274 698294 453894 698378
rect 453274 698058 453306 698294
rect 453542 698058 453626 698294
rect 453862 698058 453894 698294
rect 453274 662614 453894 698058
rect 453274 662378 453306 662614
rect 453542 662378 453626 662614
rect 453862 662378 453894 662614
rect 453274 662294 453894 662378
rect 453274 662058 453306 662294
rect 453542 662058 453626 662294
rect 453862 662058 453894 662294
rect 453274 657000 453894 662058
rect 454674 709638 455294 709670
rect 454674 709402 454706 709638
rect 454942 709402 455026 709638
rect 455262 709402 455294 709638
rect 454674 709318 455294 709402
rect 454674 709082 454706 709318
rect 454942 709082 455026 709318
rect 455262 709082 455294 709318
rect 454674 676894 455294 709082
rect 454674 676658 454706 676894
rect 454942 676658 455026 676894
rect 455262 676658 455294 676894
rect 454674 676574 455294 676658
rect 454674 676338 454706 676574
rect 454942 676338 455026 676574
rect 455262 676338 455294 676574
rect 454674 657000 455294 676338
rect 456074 706758 456694 707750
rect 456074 706522 456106 706758
rect 456342 706522 456426 706758
rect 456662 706522 456694 706758
rect 456074 706438 456694 706522
rect 456074 706202 456106 706438
rect 456342 706202 456426 706438
rect 456662 706202 456694 706438
rect 456074 691174 456694 706202
rect 456074 690938 456106 691174
rect 456342 690938 456426 691174
rect 456662 690938 456694 691174
rect 456074 690854 456694 690938
rect 456074 690618 456106 690854
rect 456342 690618 456426 690854
rect 456662 690618 456694 690854
rect 456074 657000 456694 690618
rect 457474 705798 458094 705830
rect 457474 705562 457506 705798
rect 457742 705562 457826 705798
rect 458062 705562 458094 705798
rect 457474 705478 458094 705562
rect 457474 705242 457506 705478
rect 457742 705242 457826 705478
rect 458062 705242 458094 705478
rect 457474 669454 458094 705242
rect 457474 669218 457506 669454
rect 457742 669218 457826 669454
rect 458062 669218 458094 669454
rect 457474 669134 458094 669218
rect 457474 668898 457506 669134
rect 457742 668898 457826 669134
rect 458062 668898 458094 669134
rect 457474 657000 458094 668898
rect 458394 680614 459014 711002
rect 463514 710598 464134 711590
rect 463514 710362 463546 710598
rect 463782 710362 463866 710598
rect 464102 710362 464134 710598
rect 463514 710278 464134 710362
rect 463514 710042 463546 710278
rect 463782 710042 463866 710278
rect 464102 710042 464134 710278
rect 458394 680378 458426 680614
rect 458662 680378 458746 680614
rect 458982 680378 459014 680614
rect 458394 680294 459014 680378
rect 458394 680058 458426 680294
rect 458662 680058 458746 680294
rect 458982 680058 459014 680294
rect 458394 657000 459014 680058
rect 459794 708678 460414 709670
rect 459794 708442 459826 708678
rect 460062 708442 460146 708678
rect 460382 708442 460414 708678
rect 459794 708358 460414 708442
rect 459794 708122 459826 708358
rect 460062 708122 460146 708358
rect 460382 708122 460414 708358
rect 459794 694894 460414 708122
rect 459794 694658 459826 694894
rect 460062 694658 460146 694894
rect 460382 694658 460414 694894
rect 459794 694574 460414 694658
rect 459794 694338 459826 694574
rect 460062 694338 460146 694574
rect 460382 694338 460414 694574
rect 459794 658894 460414 694338
rect 459794 658658 459826 658894
rect 460062 658658 460146 658894
rect 460382 658658 460414 658894
rect 459794 658574 460414 658658
rect 459794 658338 459826 658574
rect 460062 658338 460146 658574
rect 460382 658338 460414 658574
rect 459794 657000 460414 658338
rect 461194 707718 461814 707750
rect 461194 707482 461226 707718
rect 461462 707482 461546 707718
rect 461782 707482 461814 707718
rect 461194 707398 461814 707482
rect 461194 707162 461226 707398
rect 461462 707162 461546 707398
rect 461782 707162 461814 707398
rect 461194 673174 461814 707162
rect 461194 672938 461226 673174
rect 461462 672938 461546 673174
rect 461782 672938 461814 673174
rect 461194 672854 461814 672938
rect 461194 672618 461226 672854
rect 461462 672618 461546 672854
rect 461782 672618 461814 672854
rect 461194 657000 461814 672618
rect 462594 704838 463214 705830
rect 462594 704602 462626 704838
rect 462862 704602 462946 704838
rect 463182 704602 463214 704838
rect 462594 704518 463214 704602
rect 462594 704282 462626 704518
rect 462862 704282 462946 704518
rect 463182 704282 463214 704518
rect 462594 687454 463214 704282
rect 462594 687218 462626 687454
rect 462862 687218 462946 687454
rect 463182 687218 463214 687454
rect 462594 687134 463214 687218
rect 462594 686898 462626 687134
rect 462862 686898 462946 687134
rect 463182 686898 463214 687134
rect 462594 657000 463214 686898
rect 463514 698614 464134 710042
rect 468634 711558 469254 711590
rect 468634 711322 468666 711558
rect 468902 711322 468986 711558
rect 469222 711322 469254 711558
rect 468634 711238 469254 711322
rect 468634 711002 468666 711238
rect 468902 711002 468986 711238
rect 469222 711002 469254 711238
rect 463514 698378 463546 698614
rect 463782 698378 463866 698614
rect 464102 698378 464134 698614
rect 463514 698294 464134 698378
rect 463514 698058 463546 698294
rect 463782 698058 463866 698294
rect 464102 698058 464134 698294
rect 463514 662614 464134 698058
rect 463514 662378 463546 662614
rect 463782 662378 463866 662614
rect 464102 662378 464134 662614
rect 463514 662294 464134 662378
rect 463514 662058 463546 662294
rect 463782 662058 463866 662294
rect 464102 662058 464134 662294
rect 463514 657000 464134 662058
rect 464914 709638 465534 709670
rect 464914 709402 464946 709638
rect 465182 709402 465266 709638
rect 465502 709402 465534 709638
rect 464914 709318 465534 709402
rect 464914 709082 464946 709318
rect 465182 709082 465266 709318
rect 465502 709082 465534 709318
rect 464914 676894 465534 709082
rect 464914 676658 464946 676894
rect 465182 676658 465266 676894
rect 465502 676658 465534 676894
rect 464914 676574 465534 676658
rect 464914 676338 464946 676574
rect 465182 676338 465266 676574
rect 465502 676338 465534 676574
rect 464914 657000 465534 676338
rect 466314 706758 466934 707750
rect 466314 706522 466346 706758
rect 466582 706522 466666 706758
rect 466902 706522 466934 706758
rect 466314 706438 466934 706522
rect 466314 706202 466346 706438
rect 466582 706202 466666 706438
rect 466902 706202 466934 706438
rect 466314 691174 466934 706202
rect 466314 690938 466346 691174
rect 466582 690938 466666 691174
rect 466902 690938 466934 691174
rect 466314 690854 466934 690938
rect 466314 690618 466346 690854
rect 466582 690618 466666 690854
rect 466902 690618 466934 690854
rect 466314 657000 466934 690618
rect 467714 705798 468334 705830
rect 467714 705562 467746 705798
rect 467982 705562 468066 705798
rect 468302 705562 468334 705798
rect 467714 705478 468334 705562
rect 467714 705242 467746 705478
rect 467982 705242 468066 705478
rect 468302 705242 468334 705478
rect 467714 669454 468334 705242
rect 467714 669218 467746 669454
rect 467982 669218 468066 669454
rect 468302 669218 468334 669454
rect 467714 669134 468334 669218
rect 467714 668898 467746 669134
rect 467982 668898 468066 669134
rect 468302 668898 468334 669134
rect 467714 657000 468334 668898
rect 468634 680614 469254 711002
rect 473754 710598 474374 711590
rect 473754 710362 473786 710598
rect 474022 710362 474106 710598
rect 474342 710362 474374 710598
rect 473754 710278 474374 710362
rect 473754 710042 473786 710278
rect 474022 710042 474106 710278
rect 474342 710042 474374 710278
rect 468634 680378 468666 680614
rect 468902 680378 468986 680614
rect 469222 680378 469254 680614
rect 468634 680294 469254 680378
rect 468634 680058 468666 680294
rect 468902 680058 468986 680294
rect 469222 680058 469254 680294
rect 468634 657000 469254 680058
rect 470034 708678 470654 709670
rect 470034 708442 470066 708678
rect 470302 708442 470386 708678
rect 470622 708442 470654 708678
rect 470034 708358 470654 708442
rect 470034 708122 470066 708358
rect 470302 708122 470386 708358
rect 470622 708122 470654 708358
rect 470034 694894 470654 708122
rect 470034 694658 470066 694894
rect 470302 694658 470386 694894
rect 470622 694658 470654 694894
rect 470034 694574 470654 694658
rect 470034 694338 470066 694574
rect 470302 694338 470386 694574
rect 470622 694338 470654 694574
rect 470034 658894 470654 694338
rect 470034 658658 470066 658894
rect 470302 658658 470386 658894
rect 470622 658658 470654 658894
rect 470034 658574 470654 658658
rect 470034 658338 470066 658574
rect 470302 658338 470386 658574
rect 470622 658338 470654 658574
rect 470034 657000 470654 658338
rect 471434 707718 472054 707750
rect 471434 707482 471466 707718
rect 471702 707482 471786 707718
rect 472022 707482 472054 707718
rect 471434 707398 472054 707482
rect 471434 707162 471466 707398
rect 471702 707162 471786 707398
rect 472022 707162 472054 707398
rect 471434 673174 472054 707162
rect 471434 672938 471466 673174
rect 471702 672938 471786 673174
rect 472022 672938 472054 673174
rect 471434 672854 472054 672938
rect 471434 672618 471466 672854
rect 471702 672618 471786 672854
rect 472022 672618 472054 672854
rect 471434 657000 472054 672618
rect 472834 704838 473454 705830
rect 472834 704602 472866 704838
rect 473102 704602 473186 704838
rect 473422 704602 473454 704838
rect 472834 704518 473454 704602
rect 472834 704282 472866 704518
rect 473102 704282 473186 704518
rect 473422 704282 473454 704518
rect 472834 687454 473454 704282
rect 472834 687218 472866 687454
rect 473102 687218 473186 687454
rect 473422 687218 473454 687454
rect 472834 687134 473454 687218
rect 472834 686898 472866 687134
rect 473102 686898 473186 687134
rect 473422 686898 473454 687134
rect 472834 657000 473454 686898
rect 473754 698614 474374 710042
rect 478874 711558 479494 711590
rect 478874 711322 478906 711558
rect 479142 711322 479226 711558
rect 479462 711322 479494 711558
rect 478874 711238 479494 711322
rect 478874 711002 478906 711238
rect 479142 711002 479226 711238
rect 479462 711002 479494 711238
rect 473754 698378 473786 698614
rect 474022 698378 474106 698614
rect 474342 698378 474374 698614
rect 473754 698294 474374 698378
rect 473754 698058 473786 698294
rect 474022 698058 474106 698294
rect 474342 698058 474374 698294
rect 473754 662614 474374 698058
rect 473754 662378 473786 662614
rect 474022 662378 474106 662614
rect 474342 662378 474374 662614
rect 473754 662294 474374 662378
rect 473754 662058 473786 662294
rect 474022 662058 474106 662294
rect 474342 662058 474374 662294
rect 473754 657000 474374 662058
rect 475154 709638 475774 709670
rect 475154 709402 475186 709638
rect 475422 709402 475506 709638
rect 475742 709402 475774 709638
rect 475154 709318 475774 709402
rect 475154 709082 475186 709318
rect 475422 709082 475506 709318
rect 475742 709082 475774 709318
rect 475154 676894 475774 709082
rect 475154 676658 475186 676894
rect 475422 676658 475506 676894
rect 475742 676658 475774 676894
rect 475154 676574 475774 676658
rect 475154 676338 475186 676574
rect 475422 676338 475506 676574
rect 475742 676338 475774 676574
rect 475154 657000 475774 676338
rect 476554 706758 477174 707750
rect 476554 706522 476586 706758
rect 476822 706522 476906 706758
rect 477142 706522 477174 706758
rect 476554 706438 477174 706522
rect 476554 706202 476586 706438
rect 476822 706202 476906 706438
rect 477142 706202 477174 706438
rect 476554 691174 477174 706202
rect 476554 690938 476586 691174
rect 476822 690938 476906 691174
rect 477142 690938 477174 691174
rect 476554 690854 477174 690938
rect 476554 690618 476586 690854
rect 476822 690618 476906 690854
rect 477142 690618 477174 690854
rect 476554 657000 477174 690618
rect 477954 705798 478574 705830
rect 477954 705562 477986 705798
rect 478222 705562 478306 705798
rect 478542 705562 478574 705798
rect 477954 705478 478574 705562
rect 477954 705242 477986 705478
rect 478222 705242 478306 705478
rect 478542 705242 478574 705478
rect 477954 669454 478574 705242
rect 477954 669218 477986 669454
rect 478222 669218 478306 669454
rect 478542 669218 478574 669454
rect 477954 669134 478574 669218
rect 477954 668898 477986 669134
rect 478222 668898 478306 669134
rect 478542 668898 478574 669134
rect 477954 657000 478574 668898
rect 478874 680614 479494 711002
rect 483994 710598 484614 711590
rect 483994 710362 484026 710598
rect 484262 710362 484346 710598
rect 484582 710362 484614 710598
rect 483994 710278 484614 710362
rect 483994 710042 484026 710278
rect 484262 710042 484346 710278
rect 484582 710042 484614 710278
rect 478874 680378 478906 680614
rect 479142 680378 479226 680614
rect 479462 680378 479494 680614
rect 478874 680294 479494 680378
rect 478874 680058 478906 680294
rect 479142 680058 479226 680294
rect 479462 680058 479494 680294
rect 478874 657000 479494 680058
rect 480274 708678 480894 709670
rect 480274 708442 480306 708678
rect 480542 708442 480626 708678
rect 480862 708442 480894 708678
rect 480274 708358 480894 708442
rect 480274 708122 480306 708358
rect 480542 708122 480626 708358
rect 480862 708122 480894 708358
rect 480274 694894 480894 708122
rect 480274 694658 480306 694894
rect 480542 694658 480626 694894
rect 480862 694658 480894 694894
rect 480274 694574 480894 694658
rect 480274 694338 480306 694574
rect 480542 694338 480626 694574
rect 480862 694338 480894 694574
rect 480274 658894 480894 694338
rect 480274 658658 480306 658894
rect 480542 658658 480626 658894
rect 480862 658658 480894 658894
rect 480274 658574 480894 658658
rect 480274 658338 480306 658574
rect 480542 658338 480626 658574
rect 480862 658338 480894 658574
rect 480274 657000 480894 658338
rect 481674 707718 482294 707750
rect 481674 707482 481706 707718
rect 481942 707482 482026 707718
rect 482262 707482 482294 707718
rect 481674 707398 482294 707482
rect 481674 707162 481706 707398
rect 481942 707162 482026 707398
rect 482262 707162 482294 707398
rect 481674 673174 482294 707162
rect 481674 672938 481706 673174
rect 481942 672938 482026 673174
rect 482262 672938 482294 673174
rect 481674 672854 482294 672938
rect 481674 672618 481706 672854
rect 481942 672618 482026 672854
rect 482262 672618 482294 672854
rect 481674 657000 482294 672618
rect 483074 704838 483694 705830
rect 483074 704602 483106 704838
rect 483342 704602 483426 704838
rect 483662 704602 483694 704838
rect 483074 704518 483694 704602
rect 483074 704282 483106 704518
rect 483342 704282 483426 704518
rect 483662 704282 483694 704518
rect 483074 687454 483694 704282
rect 483074 687218 483106 687454
rect 483342 687218 483426 687454
rect 483662 687218 483694 687454
rect 483074 687134 483694 687218
rect 483074 686898 483106 687134
rect 483342 686898 483426 687134
rect 483662 686898 483694 687134
rect 483074 657000 483694 686898
rect 483994 698614 484614 710042
rect 489114 711558 489734 711590
rect 489114 711322 489146 711558
rect 489382 711322 489466 711558
rect 489702 711322 489734 711558
rect 489114 711238 489734 711322
rect 489114 711002 489146 711238
rect 489382 711002 489466 711238
rect 489702 711002 489734 711238
rect 483994 698378 484026 698614
rect 484262 698378 484346 698614
rect 484582 698378 484614 698614
rect 483994 698294 484614 698378
rect 483994 698058 484026 698294
rect 484262 698058 484346 698294
rect 484582 698058 484614 698294
rect 483994 662614 484614 698058
rect 483994 662378 484026 662614
rect 484262 662378 484346 662614
rect 484582 662378 484614 662614
rect 483994 662294 484614 662378
rect 483994 662058 484026 662294
rect 484262 662058 484346 662294
rect 484582 662058 484614 662294
rect 483994 657000 484614 662058
rect 485394 709638 486014 709670
rect 485394 709402 485426 709638
rect 485662 709402 485746 709638
rect 485982 709402 486014 709638
rect 485394 709318 486014 709402
rect 485394 709082 485426 709318
rect 485662 709082 485746 709318
rect 485982 709082 486014 709318
rect 485394 676894 486014 709082
rect 485394 676658 485426 676894
rect 485662 676658 485746 676894
rect 485982 676658 486014 676894
rect 485394 676574 486014 676658
rect 485394 676338 485426 676574
rect 485662 676338 485746 676574
rect 485982 676338 486014 676574
rect 485394 657000 486014 676338
rect 486794 706758 487414 707750
rect 486794 706522 486826 706758
rect 487062 706522 487146 706758
rect 487382 706522 487414 706758
rect 486794 706438 487414 706522
rect 486794 706202 486826 706438
rect 487062 706202 487146 706438
rect 487382 706202 487414 706438
rect 486794 691174 487414 706202
rect 486794 690938 486826 691174
rect 487062 690938 487146 691174
rect 487382 690938 487414 691174
rect 486794 690854 487414 690938
rect 486794 690618 486826 690854
rect 487062 690618 487146 690854
rect 487382 690618 487414 690854
rect 486794 657000 487414 690618
rect 488194 705798 488814 705830
rect 488194 705562 488226 705798
rect 488462 705562 488546 705798
rect 488782 705562 488814 705798
rect 488194 705478 488814 705562
rect 488194 705242 488226 705478
rect 488462 705242 488546 705478
rect 488782 705242 488814 705478
rect 488194 669454 488814 705242
rect 488194 669218 488226 669454
rect 488462 669218 488546 669454
rect 488782 669218 488814 669454
rect 488194 669134 488814 669218
rect 488194 668898 488226 669134
rect 488462 668898 488546 669134
rect 488782 668898 488814 669134
rect 488194 657000 488814 668898
rect 489114 680614 489734 711002
rect 494234 710598 494854 711590
rect 494234 710362 494266 710598
rect 494502 710362 494586 710598
rect 494822 710362 494854 710598
rect 494234 710278 494854 710362
rect 494234 710042 494266 710278
rect 494502 710042 494586 710278
rect 494822 710042 494854 710278
rect 489114 680378 489146 680614
rect 489382 680378 489466 680614
rect 489702 680378 489734 680614
rect 489114 680294 489734 680378
rect 489114 680058 489146 680294
rect 489382 680058 489466 680294
rect 489702 680058 489734 680294
rect 489114 657000 489734 680058
rect 490514 708678 491134 709670
rect 490514 708442 490546 708678
rect 490782 708442 490866 708678
rect 491102 708442 491134 708678
rect 490514 708358 491134 708442
rect 490514 708122 490546 708358
rect 490782 708122 490866 708358
rect 491102 708122 491134 708358
rect 490514 694894 491134 708122
rect 490514 694658 490546 694894
rect 490782 694658 490866 694894
rect 491102 694658 491134 694894
rect 490514 694574 491134 694658
rect 490514 694338 490546 694574
rect 490782 694338 490866 694574
rect 491102 694338 491134 694574
rect 490514 658894 491134 694338
rect 490514 658658 490546 658894
rect 490782 658658 490866 658894
rect 491102 658658 491134 658894
rect 490514 658574 491134 658658
rect 490514 658338 490546 658574
rect 490782 658338 490866 658574
rect 491102 658338 491134 658574
rect 490514 657000 491134 658338
rect 491914 707718 492534 707750
rect 491914 707482 491946 707718
rect 492182 707482 492266 707718
rect 492502 707482 492534 707718
rect 491914 707398 492534 707482
rect 491914 707162 491946 707398
rect 492182 707162 492266 707398
rect 492502 707162 492534 707398
rect 491914 673174 492534 707162
rect 491914 672938 491946 673174
rect 492182 672938 492266 673174
rect 492502 672938 492534 673174
rect 491914 672854 492534 672938
rect 491914 672618 491946 672854
rect 492182 672618 492266 672854
rect 492502 672618 492534 672854
rect 491914 657000 492534 672618
rect 493314 704838 493934 705830
rect 493314 704602 493346 704838
rect 493582 704602 493666 704838
rect 493902 704602 493934 704838
rect 493314 704518 493934 704602
rect 493314 704282 493346 704518
rect 493582 704282 493666 704518
rect 493902 704282 493934 704518
rect 493314 687454 493934 704282
rect 493314 687218 493346 687454
rect 493582 687218 493666 687454
rect 493902 687218 493934 687454
rect 493314 687134 493934 687218
rect 493314 686898 493346 687134
rect 493582 686898 493666 687134
rect 493902 686898 493934 687134
rect 493314 657000 493934 686898
rect 494234 698614 494854 710042
rect 499354 711558 499974 711590
rect 499354 711322 499386 711558
rect 499622 711322 499706 711558
rect 499942 711322 499974 711558
rect 499354 711238 499974 711322
rect 499354 711002 499386 711238
rect 499622 711002 499706 711238
rect 499942 711002 499974 711238
rect 494234 698378 494266 698614
rect 494502 698378 494586 698614
rect 494822 698378 494854 698614
rect 494234 698294 494854 698378
rect 494234 698058 494266 698294
rect 494502 698058 494586 698294
rect 494822 698058 494854 698294
rect 494234 662614 494854 698058
rect 494234 662378 494266 662614
rect 494502 662378 494586 662614
rect 494822 662378 494854 662614
rect 494234 662294 494854 662378
rect 494234 662058 494266 662294
rect 494502 662058 494586 662294
rect 494822 662058 494854 662294
rect 494234 657000 494854 662058
rect 495634 709638 496254 709670
rect 495634 709402 495666 709638
rect 495902 709402 495986 709638
rect 496222 709402 496254 709638
rect 495634 709318 496254 709402
rect 495634 709082 495666 709318
rect 495902 709082 495986 709318
rect 496222 709082 496254 709318
rect 495634 676894 496254 709082
rect 495634 676658 495666 676894
rect 495902 676658 495986 676894
rect 496222 676658 496254 676894
rect 495634 676574 496254 676658
rect 495634 676338 495666 676574
rect 495902 676338 495986 676574
rect 496222 676338 496254 676574
rect 495634 657000 496254 676338
rect 497034 706758 497654 707750
rect 497034 706522 497066 706758
rect 497302 706522 497386 706758
rect 497622 706522 497654 706758
rect 497034 706438 497654 706522
rect 497034 706202 497066 706438
rect 497302 706202 497386 706438
rect 497622 706202 497654 706438
rect 497034 691174 497654 706202
rect 497034 690938 497066 691174
rect 497302 690938 497386 691174
rect 497622 690938 497654 691174
rect 497034 690854 497654 690938
rect 497034 690618 497066 690854
rect 497302 690618 497386 690854
rect 497622 690618 497654 690854
rect 497034 657000 497654 690618
rect 498434 705798 499054 705830
rect 498434 705562 498466 705798
rect 498702 705562 498786 705798
rect 499022 705562 499054 705798
rect 498434 705478 499054 705562
rect 498434 705242 498466 705478
rect 498702 705242 498786 705478
rect 499022 705242 499054 705478
rect 498434 669454 499054 705242
rect 498434 669218 498466 669454
rect 498702 669218 498786 669454
rect 499022 669218 499054 669454
rect 498434 669134 499054 669218
rect 498434 668898 498466 669134
rect 498702 668898 498786 669134
rect 499022 668898 499054 669134
rect 498434 657000 499054 668898
rect 499354 680614 499974 711002
rect 504474 710598 505094 711590
rect 504474 710362 504506 710598
rect 504742 710362 504826 710598
rect 505062 710362 505094 710598
rect 504474 710278 505094 710362
rect 504474 710042 504506 710278
rect 504742 710042 504826 710278
rect 505062 710042 505094 710278
rect 499354 680378 499386 680614
rect 499622 680378 499706 680614
rect 499942 680378 499974 680614
rect 499354 680294 499974 680378
rect 499354 680058 499386 680294
rect 499622 680058 499706 680294
rect 499942 680058 499974 680294
rect 499354 657000 499974 680058
rect 500754 708678 501374 709670
rect 500754 708442 500786 708678
rect 501022 708442 501106 708678
rect 501342 708442 501374 708678
rect 500754 708358 501374 708442
rect 500754 708122 500786 708358
rect 501022 708122 501106 708358
rect 501342 708122 501374 708358
rect 500754 694894 501374 708122
rect 500754 694658 500786 694894
rect 501022 694658 501106 694894
rect 501342 694658 501374 694894
rect 500754 694574 501374 694658
rect 500754 694338 500786 694574
rect 501022 694338 501106 694574
rect 501342 694338 501374 694574
rect 500754 658894 501374 694338
rect 500754 658658 500786 658894
rect 501022 658658 501106 658894
rect 501342 658658 501374 658894
rect 500754 658574 501374 658658
rect 500754 658338 500786 658574
rect 501022 658338 501106 658574
rect 501342 658338 501374 658574
rect 500754 657000 501374 658338
rect 502154 707718 502774 707750
rect 502154 707482 502186 707718
rect 502422 707482 502506 707718
rect 502742 707482 502774 707718
rect 502154 707398 502774 707482
rect 502154 707162 502186 707398
rect 502422 707162 502506 707398
rect 502742 707162 502774 707398
rect 502154 673174 502774 707162
rect 502154 672938 502186 673174
rect 502422 672938 502506 673174
rect 502742 672938 502774 673174
rect 502154 672854 502774 672938
rect 502154 672618 502186 672854
rect 502422 672618 502506 672854
rect 502742 672618 502774 672854
rect 502154 657000 502774 672618
rect 503554 704838 504174 705830
rect 503554 704602 503586 704838
rect 503822 704602 503906 704838
rect 504142 704602 504174 704838
rect 503554 704518 504174 704602
rect 503554 704282 503586 704518
rect 503822 704282 503906 704518
rect 504142 704282 504174 704518
rect 503554 687454 504174 704282
rect 503554 687218 503586 687454
rect 503822 687218 503906 687454
rect 504142 687218 504174 687454
rect 503554 687134 504174 687218
rect 503554 686898 503586 687134
rect 503822 686898 503906 687134
rect 504142 686898 504174 687134
rect 503554 657000 504174 686898
rect 504474 698614 505094 710042
rect 509594 711558 510214 711590
rect 509594 711322 509626 711558
rect 509862 711322 509946 711558
rect 510182 711322 510214 711558
rect 509594 711238 510214 711322
rect 509594 711002 509626 711238
rect 509862 711002 509946 711238
rect 510182 711002 510214 711238
rect 504474 698378 504506 698614
rect 504742 698378 504826 698614
rect 505062 698378 505094 698614
rect 504474 698294 505094 698378
rect 504474 698058 504506 698294
rect 504742 698058 504826 698294
rect 505062 698058 505094 698294
rect 504474 662614 505094 698058
rect 504474 662378 504506 662614
rect 504742 662378 504826 662614
rect 505062 662378 505094 662614
rect 504474 662294 505094 662378
rect 504474 662058 504506 662294
rect 504742 662058 504826 662294
rect 505062 662058 505094 662294
rect 504474 657000 505094 662058
rect 505874 709638 506494 709670
rect 505874 709402 505906 709638
rect 506142 709402 506226 709638
rect 506462 709402 506494 709638
rect 505874 709318 506494 709402
rect 505874 709082 505906 709318
rect 506142 709082 506226 709318
rect 506462 709082 506494 709318
rect 505874 676894 506494 709082
rect 505874 676658 505906 676894
rect 506142 676658 506226 676894
rect 506462 676658 506494 676894
rect 505874 676574 506494 676658
rect 505874 676338 505906 676574
rect 506142 676338 506226 676574
rect 506462 676338 506494 676574
rect 505874 657000 506494 676338
rect 507274 706758 507894 707750
rect 507274 706522 507306 706758
rect 507542 706522 507626 706758
rect 507862 706522 507894 706758
rect 507274 706438 507894 706522
rect 507274 706202 507306 706438
rect 507542 706202 507626 706438
rect 507862 706202 507894 706438
rect 507274 691174 507894 706202
rect 507274 690938 507306 691174
rect 507542 690938 507626 691174
rect 507862 690938 507894 691174
rect 507274 690854 507894 690938
rect 507274 690618 507306 690854
rect 507542 690618 507626 690854
rect 507862 690618 507894 690854
rect 507274 657000 507894 690618
rect 508674 705798 509294 705830
rect 508674 705562 508706 705798
rect 508942 705562 509026 705798
rect 509262 705562 509294 705798
rect 508674 705478 509294 705562
rect 508674 705242 508706 705478
rect 508942 705242 509026 705478
rect 509262 705242 509294 705478
rect 508674 669454 509294 705242
rect 508674 669218 508706 669454
rect 508942 669218 509026 669454
rect 509262 669218 509294 669454
rect 508674 669134 509294 669218
rect 508674 668898 508706 669134
rect 508942 668898 509026 669134
rect 509262 668898 509294 669134
rect 508674 657000 509294 668898
rect 509594 680614 510214 711002
rect 514714 710598 515334 711590
rect 514714 710362 514746 710598
rect 514982 710362 515066 710598
rect 515302 710362 515334 710598
rect 514714 710278 515334 710362
rect 514714 710042 514746 710278
rect 514982 710042 515066 710278
rect 515302 710042 515334 710278
rect 509594 680378 509626 680614
rect 509862 680378 509946 680614
rect 510182 680378 510214 680614
rect 509594 680294 510214 680378
rect 509594 680058 509626 680294
rect 509862 680058 509946 680294
rect 510182 680058 510214 680294
rect 509594 657000 510214 680058
rect 510994 708678 511614 709670
rect 510994 708442 511026 708678
rect 511262 708442 511346 708678
rect 511582 708442 511614 708678
rect 510994 708358 511614 708442
rect 510994 708122 511026 708358
rect 511262 708122 511346 708358
rect 511582 708122 511614 708358
rect 510994 694894 511614 708122
rect 510994 694658 511026 694894
rect 511262 694658 511346 694894
rect 511582 694658 511614 694894
rect 510994 694574 511614 694658
rect 510994 694338 511026 694574
rect 511262 694338 511346 694574
rect 511582 694338 511614 694574
rect 510994 658894 511614 694338
rect 510994 658658 511026 658894
rect 511262 658658 511346 658894
rect 511582 658658 511614 658894
rect 510994 658574 511614 658658
rect 510994 658338 511026 658574
rect 511262 658338 511346 658574
rect 511582 658338 511614 658574
rect 510994 657000 511614 658338
rect 512394 707718 513014 707750
rect 512394 707482 512426 707718
rect 512662 707482 512746 707718
rect 512982 707482 513014 707718
rect 512394 707398 513014 707482
rect 512394 707162 512426 707398
rect 512662 707162 512746 707398
rect 512982 707162 513014 707398
rect 512394 673174 513014 707162
rect 512394 672938 512426 673174
rect 512662 672938 512746 673174
rect 512982 672938 513014 673174
rect 512394 672854 513014 672938
rect 512394 672618 512426 672854
rect 512662 672618 512746 672854
rect 512982 672618 513014 672854
rect 512394 657000 513014 672618
rect 513794 704838 514414 705830
rect 513794 704602 513826 704838
rect 514062 704602 514146 704838
rect 514382 704602 514414 704838
rect 513794 704518 514414 704602
rect 513794 704282 513826 704518
rect 514062 704282 514146 704518
rect 514382 704282 514414 704518
rect 513794 687454 514414 704282
rect 513794 687218 513826 687454
rect 514062 687218 514146 687454
rect 514382 687218 514414 687454
rect 513794 687134 514414 687218
rect 513794 686898 513826 687134
rect 514062 686898 514146 687134
rect 514382 686898 514414 687134
rect 513794 657000 514414 686898
rect 514714 698614 515334 710042
rect 519834 711558 520454 711590
rect 519834 711322 519866 711558
rect 520102 711322 520186 711558
rect 520422 711322 520454 711558
rect 519834 711238 520454 711322
rect 519834 711002 519866 711238
rect 520102 711002 520186 711238
rect 520422 711002 520454 711238
rect 514714 698378 514746 698614
rect 514982 698378 515066 698614
rect 515302 698378 515334 698614
rect 514714 698294 515334 698378
rect 514714 698058 514746 698294
rect 514982 698058 515066 698294
rect 515302 698058 515334 698294
rect 514714 662614 515334 698058
rect 514714 662378 514746 662614
rect 514982 662378 515066 662614
rect 515302 662378 515334 662614
rect 514714 662294 515334 662378
rect 514714 662058 514746 662294
rect 514982 662058 515066 662294
rect 515302 662058 515334 662294
rect 514714 657000 515334 662058
rect 516114 709638 516734 709670
rect 516114 709402 516146 709638
rect 516382 709402 516466 709638
rect 516702 709402 516734 709638
rect 516114 709318 516734 709402
rect 516114 709082 516146 709318
rect 516382 709082 516466 709318
rect 516702 709082 516734 709318
rect 516114 676894 516734 709082
rect 516114 676658 516146 676894
rect 516382 676658 516466 676894
rect 516702 676658 516734 676894
rect 516114 676574 516734 676658
rect 516114 676338 516146 676574
rect 516382 676338 516466 676574
rect 516702 676338 516734 676574
rect 516114 657000 516734 676338
rect 517514 706758 518134 707750
rect 517514 706522 517546 706758
rect 517782 706522 517866 706758
rect 518102 706522 518134 706758
rect 517514 706438 518134 706522
rect 517514 706202 517546 706438
rect 517782 706202 517866 706438
rect 518102 706202 518134 706438
rect 517514 691174 518134 706202
rect 517514 690938 517546 691174
rect 517782 690938 517866 691174
rect 518102 690938 518134 691174
rect 517514 690854 518134 690938
rect 517514 690618 517546 690854
rect 517782 690618 517866 690854
rect 518102 690618 518134 690854
rect 517514 657000 518134 690618
rect 518914 705798 519534 705830
rect 518914 705562 518946 705798
rect 519182 705562 519266 705798
rect 519502 705562 519534 705798
rect 518914 705478 519534 705562
rect 518914 705242 518946 705478
rect 519182 705242 519266 705478
rect 519502 705242 519534 705478
rect 518914 669454 519534 705242
rect 518914 669218 518946 669454
rect 519182 669218 519266 669454
rect 519502 669218 519534 669454
rect 518914 669134 519534 669218
rect 518914 668898 518946 669134
rect 519182 668898 519266 669134
rect 519502 668898 519534 669134
rect 518914 657000 519534 668898
rect 519834 680614 520454 711002
rect 524954 710598 525574 711590
rect 524954 710362 524986 710598
rect 525222 710362 525306 710598
rect 525542 710362 525574 710598
rect 524954 710278 525574 710362
rect 524954 710042 524986 710278
rect 525222 710042 525306 710278
rect 525542 710042 525574 710278
rect 519834 680378 519866 680614
rect 520102 680378 520186 680614
rect 520422 680378 520454 680614
rect 519834 680294 520454 680378
rect 519834 680058 519866 680294
rect 520102 680058 520186 680294
rect 520422 680058 520454 680294
rect 519834 657000 520454 680058
rect 521234 708678 521854 709670
rect 521234 708442 521266 708678
rect 521502 708442 521586 708678
rect 521822 708442 521854 708678
rect 521234 708358 521854 708442
rect 521234 708122 521266 708358
rect 521502 708122 521586 708358
rect 521822 708122 521854 708358
rect 521234 694894 521854 708122
rect 521234 694658 521266 694894
rect 521502 694658 521586 694894
rect 521822 694658 521854 694894
rect 521234 694574 521854 694658
rect 521234 694338 521266 694574
rect 521502 694338 521586 694574
rect 521822 694338 521854 694574
rect 521234 658894 521854 694338
rect 521234 658658 521266 658894
rect 521502 658658 521586 658894
rect 521822 658658 521854 658894
rect 521234 658574 521854 658658
rect 521234 658338 521266 658574
rect 521502 658338 521586 658574
rect 521822 658338 521854 658574
rect 521234 657000 521854 658338
rect 522634 707718 523254 707750
rect 522634 707482 522666 707718
rect 522902 707482 522986 707718
rect 523222 707482 523254 707718
rect 522634 707398 523254 707482
rect 522634 707162 522666 707398
rect 522902 707162 522986 707398
rect 523222 707162 523254 707398
rect 522634 673174 523254 707162
rect 522634 672938 522666 673174
rect 522902 672938 522986 673174
rect 523222 672938 523254 673174
rect 522634 672854 523254 672938
rect 522634 672618 522666 672854
rect 522902 672618 522986 672854
rect 523222 672618 523254 672854
rect 522634 657000 523254 672618
rect 524034 704838 524654 705830
rect 524034 704602 524066 704838
rect 524302 704602 524386 704838
rect 524622 704602 524654 704838
rect 524034 704518 524654 704602
rect 524034 704282 524066 704518
rect 524302 704282 524386 704518
rect 524622 704282 524654 704518
rect 524034 687454 524654 704282
rect 524034 687218 524066 687454
rect 524302 687218 524386 687454
rect 524622 687218 524654 687454
rect 524034 687134 524654 687218
rect 524034 686898 524066 687134
rect 524302 686898 524386 687134
rect 524622 686898 524654 687134
rect 524034 657000 524654 686898
rect 524954 698614 525574 710042
rect 530074 711558 530694 711590
rect 530074 711322 530106 711558
rect 530342 711322 530426 711558
rect 530662 711322 530694 711558
rect 530074 711238 530694 711322
rect 530074 711002 530106 711238
rect 530342 711002 530426 711238
rect 530662 711002 530694 711238
rect 524954 698378 524986 698614
rect 525222 698378 525306 698614
rect 525542 698378 525574 698614
rect 524954 698294 525574 698378
rect 524954 698058 524986 698294
rect 525222 698058 525306 698294
rect 525542 698058 525574 698294
rect 524954 662614 525574 698058
rect 524954 662378 524986 662614
rect 525222 662378 525306 662614
rect 525542 662378 525574 662614
rect 524954 662294 525574 662378
rect 524954 662058 524986 662294
rect 525222 662058 525306 662294
rect 525542 662058 525574 662294
rect 524954 657000 525574 662058
rect 526354 709638 526974 709670
rect 526354 709402 526386 709638
rect 526622 709402 526706 709638
rect 526942 709402 526974 709638
rect 526354 709318 526974 709402
rect 526354 709082 526386 709318
rect 526622 709082 526706 709318
rect 526942 709082 526974 709318
rect 526354 676894 526974 709082
rect 526354 676658 526386 676894
rect 526622 676658 526706 676894
rect 526942 676658 526974 676894
rect 526354 676574 526974 676658
rect 526354 676338 526386 676574
rect 526622 676338 526706 676574
rect 526942 676338 526974 676574
rect 526354 657000 526974 676338
rect 527754 706758 528374 707750
rect 527754 706522 527786 706758
rect 528022 706522 528106 706758
rect 528342 706522 528374 706758
rect 527754 706438 528374 706522
rect 527754 706202 527786 706438
rect 528022 706202 528106 706438
rect 528342 706202 528374 706438
rect 527754 691174 528374 706202
rect 527754 690938 527786 691174
rect 528022 690938 528106 691174
rect 528342 690938 528374 691174
rect 527754 690854 528374 690938
rect 527754 690618 527786 690854
rect 528022 690618 528106 690854
rect 528342 690618 528374 690854
rect 527754 657000 528374 690618
rect 529154 705798 529774 705830
rect 529154 705562 529186 705798
rect 529422 705562 529506 705798
rect 529742 705562 529774 705798
rect 529154 705478 529774 705562
rect 529154 705242 529186 705478
rect 529422 705242 529506 705478
rect 529742 705242 529774 705478
rect 529154 669454 529774 705242
rect 529154 669218 529186 669454
rect 529422 669218 529506 669454
rect 529742 669218 529774 669454
rect 529154 669134 529774 669218
rect 529154 668898 529186 669134
rect 529422 668898 529506 669134
rect 529742 668898 529774 669134
rect 529154 657000 529774 668898
rect 530074 680614 530694 711002
rect 535194 710598 535814 711590
rect 535194 710362 535226 710598
rect 535462 710362 535546 710598
rect 535782 710362 535814 710598
rect 535194 710278 535814 710362
rect 535194 710042 535226 710278
rect 535462 710042 535546 710278
rect 535782 710042 535814 710278
rect 530074 680378 530106 680614
rect 530342 680378 530426 680614
rect 530662 680378 530694 680614
rect 530074 680294 530694 680378
rect 530074 680058 530106 680294
rect 530342 680058 530426 680294
rect 530662 680058 530694 680294
rect 530074 657000 530694 680058
rect 531474 708678 532094 709670
rect 531474 708442 531506 708678
rect 531742 708442 531826 708678
rect 532062 708442 532094 708678
rect 531474 708358 532094 708442
rect 531474 708122 531506 708358
rect 531742 708122 531826 708358
rect 532062 708122 532094 708358
rect 531474 694894 532094 708122
rect 531474 694658 531506 694894
rect 531742 694658 531826 694894
rect 532062 694658 532094 694894
rect 531474 694574 532094 694658
rect 531474 694338 531506 694574
rect 531742 694338 531826 694574
rect 532062 694338 532094 694574
rect 531474 658894 532094 694338
rect 531474 658658 531506 658894
rect 531742 658658 531826 658894
rect 532062 658658 532094 658894
rect 531474 658574 532094 658658
rect 531474 658338 531506 658574
rect 531742 658338 531826 658574
rect 532062 658338 532094 658574
rect 531474 657000 532094 658338
rect 532874 707718 533494 707750
rect 532874 707482 532906 707718
rect 533142 707482 533226 707718
rect 533462 707482 533494 707718
rect 532874 707398 533494 707482
rect 532874 707162 532906 707398
rect 533142 707162 533226 707398
rect 533462 707162 533494 707398
rect 532874 673174 533494 707162
rect 532874 672938 532906 673174
rect 533142 672938 533226 673174
rect 533462 672938 533494 673174
rect 532874 672854 533494 672938
rect 532874 672618 532906 672854
rect 533142 672618 533226 672854
rect 533462 672618 533494 672854
rect 532874 657000 533494 672618
rect 534274 704838 534894 705830
rect 534274 704602 534306 704838
rect 534542 704602 534626 704838
rect 534862 704602 534894 704838
rect 534274 704518 534894 704602
rect 534274 704282 534306 704518
rect 534542 704282 534626 704518
rect 534862 704282 534894 704518
rect 534274 687454 534894 704282
rect 534274 687218 534306 687454
rect 534542 687218 534626 687454
rect 534862 687218 534894 687454
rect 534274 687134 534894 687218
rect 534274 686898 534306 687134
rect 534542 686898 534626 687134
rect 534862 686898 534894 687134
rect 534274 657000 534894 686898
rect 535194 698614 535814 710042
rect 540314 711558 540934 711590
rect 540314 711322 540346 711558
rect 540582 711322 540666 711558
rect 540902 711322 540934 711558
rect 540314 711238 540934 711322
rect 540314 711002 540346 711238
rect 540582 711002 540666 711238
rect 540902 711002 540934 711238
rect 535194 698378 535226 698614
rect 535462 698378 535546 698614
rect 535782 698378 535814 698614
rect 535194 698294 535814 698378
rect 535194 698058 535226 698294
rect 535462 698058 535546 698294
rect 535782 698058 535814 698294
rect 535194 662614 535814 698058
rect 535194 662378 535226 662614
rect 535462 662378 535546 662614
rect 535782 662378 535814 662614
rect 535194 662294 535814 662378
rect 535194 662058 535226 662294
rect 535462 662058 535546 662294
rect 535782 662058 535814 662294
rect 535194 657000 535814 662058
rect 536594 709638 537214 709670
rect 536594 709402 536626 709638
rect 536862 709402 536946 709638
rect 537182 709402 537214 709638
rect 536594 709318 537214 709402
rect 536594 709082 536626 709318
rect 536862 709082 536946 709318
rect 537182 709082 537214 709318
rect 536594 676894 537214 709082
rect 536594 676658 536626 676894
rect 536862 676658 536946 676894
rect 537182 676658 537214 676894
rect 536594 676574 537214 676658
rect 536594 676338 536626 676574
rect 536862 676338 536946 676574
rect 537182 676338 537214 676574
rect 536594 657000 537214 676338
rect 537994 706758 538614 707750
rect 537994 706522 538026 706758
rect 538262 706522 538346 706758
rect 538582 706522 538614 706758
rect 537994 706438 538614 706522
rect 537994 706202 538026 706438
rect 538262 706202 538346 706438
rect 538582 706202 538614 706438
rect 537994 691174 538614 706202
rect 537994 690938 538026 691174
rect 538262 690938 538346 691174
rect 538582 690938 538614 691174
rect 537994 690854 538614 690938
rect 537994 690618 538026 690854
rect 538262 690618 538346 690854
rect 538582 690618 538614 690854
rect 537994 657000 538614 690618
rect 539394 705798 540014 705830
rect 539394 705562 539426 705798
rect 539662 705562 539746 705798
rect 539982 705562 540014 705798
rect 539394 705478 540014 705562
rect 539394 705242 539426 705478
rect 539662 705242 539746 705478
rect 539982 705242 540014 705478
rect 539394 669454 540014 705242
rect 539394 669218 539426 669454
rect 539662 669218 539746 669454
rect 539982 669218 540014 669454
rect 539394 669134 540014 669218
rect 539394 668898 539426 669134
rect 539662 668898 539746 669134
rect 539982 668898 540014 669134
rect 539394 657000 540014 668898
rect 540314 680614 540934 711002
rect 545434 710598 546054 711590
rect 545434 710362 545466 710598
rect 545702 710362 545786 710598
rect 546022 710362 546054 710598
rect 545434 710278 546054 710362
rect 545434 710042 545466 710278
rect 545702 710042 545786 710278
rect 546022 710042 546054 710278
rect 540314 680378 540346 680614
rect 540582 680378 540666 680614
rect 540902 680378 540934 680614
rect 540314 680294 540934 680378
rect 540314 680058 540346 680294
rect 540582 680058 540666 680294
rect 540902 680058 540934 680294
rect 540314 657000 540934 680058
rect 541714 708678 542334 709670
rect 541714 708442 541746 708678
rect 541982 708442 542066 708678
rect 542302 708442 542334 708678
rect 541714 708358 542334 708442
rect 541714 708122 541746 708358
rect 541982 708122 542066 708358
rect 542302 708122 542334 708358
rect 541714 694894 542334 708122
rect 541714 694658 541746 694894
rect 541982 694658 542066 694894
rect 542302 694658 542334 694894
rect 541714 694574 542334 694658
rect 541714 694338 541746 694574
rect 541982 694338 542066 694574
rect 542302 694338 542334 694574
rect 541714 658894 542334 694338
rect 541714 658658 541746 658894
rect 541982 658658 542066 658894
rect 542302 658658 542334 658894
rect 541714 658574 542334 658658
rect 541714 658338 541746 658574
rect 541982 658338 542066 658574
rect 542302 658338 542334 658574
rect 15754 654938 15786 655174
rect 16022 654938 16106 655174
rect 16342 654938 16374 655174
rect 15754 654854 16374 654938
rect 15754 654618 15786 654854
rect 16022 654618 16106 654854
rect 16342 654618 16374 654854
rect 15754 619174 16374 654618
rect 23288 651454 23608 651486
rect 23288 651218 23330 651454
rect 23566 651218 23608 651454
rect 23288 651134 23608 651218
rect 23288 650898 23330 651134
rect 23566 650898 23608 651134
rect 23288 650866 23608 650898
rect 33528 651454 33848 651486
rect 33528 651218 33570 651454
rect 33806 651218 33848 651454
rect 33528 651134 33848 651218
rect 33528 650898 33570 651134
rect 33806 650898 33848 651134
rect 33528 650866 33848 650898
rect 43768 651454 44088 651486
rect 43768 651218 43810 651454
rect 44046 651218 44088 651454
rect 43768 651134 44088 651218
rect 43768 650898 43810 651134
rect 44046 650898 44088 651134
rect 43768 650866 44088 650898
rect 54008 651454 54328 651486
rect 54008 651218 54050 651454
rect 54286 651218 54328 651454
rect 54008 651134 54328 651218
rect 54008 650898 54050 651134
rect 54286 650898 54328 651134
rect 54008 650866 54328 650898
rect 64248 651454 64568 651486
rect 64248 651218 64290 651454
rect 64526 651218 64568 651454
rect 64248 651134 64568 651218
rect 64248 650898 64290 651134
rect 64526 650898 64568 651134
rect 64248 650866 64568 650898
rect 74488 651454 74808 651486
rect 74488 651218 74530 651454
rect 74766 651218 74808 651454
rect 74488 651134 74808 651218
rect 74488 650898 74530 651134
rect 74766 650898 74808 651134
rect 74488 650866 74808 650898
rect 84728 651454 85048 651486
rect 84728 651218 84770 651454
rect 85006 651218 85048 651454
rect 84728 651134 85048 651218
rect 84728 650898 84770 651134
rect 85006 650898 85048 651134
rect 84728 650866 85048 650898
rect 94968 651454 95288 651486
rect 94968 651218 95010 651454
rect 95246 651218 95288 651454
rect 94968 651134 95288 651218
rect 94968 650898 95010 651134
rect 95246 650898 95288 651134
rect 94968 650866 95288 650898
rect 105208 651454 105528 651486
rect 105208 651218 105250 651454
rect 105486 651218 105528 651454
rect 105208 651134 105528 651218
rect 105208 650898 105250 651134
rect 105486 650898 105528 651134
rect 105208 650866 105528 650898
rect 115448 651454 115768 651486
rect 115448 651218 115490 651454
rect 115726 651218 115768 651454
rect 115448 651134 115768 651218
rect 115448 650898 115490 651134
rect 115726 650898 115768 651134
rect 115448 650866 115768 650898
rect 125688 651454 126008 651486
rect 125688 651218 125730 651454
rect 125966 651218 126008 651454
rect 125688 651134 126008 651218
rect 125688 650898 125730 651134
rect 125966 650898 126008 651134
rect 125688 650866 126008 650898
rect 135928 651454 136248 651486
rect 135928 651218 135970 651454
rect 136206 651218 136248 651454
rect 135928 651134 136248 651218
rect 135928 650898 135970 651134
rect 136206 650898 136248 651134
rect 135928 650866 136248 650898
rect 146168 651454 146488 651486
rect 146168 651218 146210 651454
rect 146446 651218 146488 651454
rect 146168 651134 146488 651218
rect 146168 650898 146210 651134
rect 146446 650898 146488 651134
rect 146168 650866 146488 650898
rect 156408 651454 156728 651486
rect 156408 651218 156450 651454
rect 156686 651218 156728 651454
rect 156408 651134 156728 651218
rect 156408 650898 156450 651134
rect 156686 650898 156728 651134
rect 156408 650866 156728 650898
rect 166648 651454 166968 651486
rect 166648 651218 166690 651454
rect 166926 651218 166968 651454
rect 166648 651134 166968 651218
rect 166648 650898 166690 651134
rect 166926 650898 166968 651134
rect 166648 650866 166968 650898
rect 176888 651454 177208 651486
rect 176888 651218 176930 651454
rect 177166 651218 177208 651454
rect 176888 651134 177208 651218
rect 176888 650898 176930 651134
rect 177166 650898 177208 651134
rect 176888 650866 177208 650898
rect 187128 651454 187448 651486
rect 187128 651218 187170 651454
rect 187406 651218 187448 651454
rect 187128 651134 187448 651218
rect 187128 650898 187170 651134
rect 187406 650898 187448 651134
rect 187128 650866 187448 650898
rect 197368 651454 197688 651486
rect 197368 651218 197410 651454
rect 197646 651218 197688 651454
rect 197368 651134 197688 651218
rect 197368 650898 197410 651134
rect 197646 650898 197688 651134
rect 197368 650866 197688 650898
rect 207608 651454 207928 651486
rect 207608 651218 207650 651454
rect 207886 651218 207928 651454
rect 207608 651134 207928 651218
rect 207608 650898 207650 651134
rect 207886 650898 207928 651134
rect 207608 650866 207928 650898
rect 217848 651454 218168 651486
rect 217848 651218 217890 651454
rect 218126 651218 218168 651454
rect 217848 651134 218168 651218
rect 217848 650898 217890 651134
rect 218126 650898 218168 651134
rect 217848 650866 218168 650898
rect 228088 651454 228408 651486
rect 228088 651218 228130 651454
rect 228366 651218 228408 651454
rect 228088 651134 228408 651218
rect 228088 650898 228130 651134
rect 228366 650898 228408 651134
rect 228088 650866 228408 650898
rect 238328 651454 238648 651486
rect 238328 651218 238370 651454
rect 238606 651218 238648 651454
rect 238328 651134 238648 651218
rect 238328 650898 238370 651134
rect 238606 650898 238648 651134
rect 238328 650866 238648 650898
rect 248568 651454 248888 651486
rect 248568 651218 248610 651454
rect 248846 651218 248888 651454
rect 248568 651134 248888 651218
rect 248568 650898 248610 651134
rect 248846 650898 248888 651134
rect 248568 650866 248888 650898
rect 258808 651454 259128 651486
rect 258808 651218 258850 651454
rect 259086 651218 259128 651454
rect 258808 651134 259128 651218
rect 258808 650898 258850 651134
rect 259086 650898 259128 651134
rect 258808 650866 259128 650898
rect 269048 651454 269368 651486
rect 269048 651218 269090 651454
rect 269326 651218 269368 651454
rect 269048 651134 269368 651218
rect 269048 650898 269090 651134
rect 269326 650898 269368 651134
rect 269048 650866 269368 650898
rect 279288 651454 279608 651486
rect 279288 651218 279330 651454
rect 279566 651218 279608 651454
rect 279288 651134 279608 651218
rect 279288 650898 279330 651134
rect 279566 650898 279608 651134
rect 279288 650866 279608 650898
rect 289528 651454 289848 651486
rect 289528 651218 289570 651454
rect 289806 651218 289848 651454
rect 289528 651134 289848 651218
rect 289528 650898 289570 651134
rect 289806 650898 289848 651134
rect 289528 650866 289848 650898
rect 299768 651454 300088 651486
rect 299768 651218 299810 651454
rect 300046 651218 300088 651454
rect 299768 651134 300088 651218
rect 299768 650898 299810 651134
rect 300046 650898 300088 651134
rect 299768 650866 300088 650898
rect 310008 651454 310328 651486
rect 310008 651218 310050 651454
rect 310286 651218 310328 651454
rect 310008 651134 310328 651218
rect 310008 650898 310050 651134
rect 310286 650898 310328 651134
rect 310008 650866 310328 650898
rect 320248 651454 320568 651486
rect 320248 651218 320290 651454
rect 320526 651218 320568 651454
rect 320248 651134 320568 651218
rect 320248 650898 320290 651134
rect 320526 650898 320568 651134
rect 320248 650866 320568 650898
rect 330488 651454 330808 651486
rect 330488 651218 330530 651454
rect 330766 651218 330808 651454
rect 330488 651134 330808 651218
rect 330488 650898 330530 651134
rect 330766 650898 330808 651134
rect 330488 650866 330808 650898
rect 340728 651454 341048 651486
rect 340728 651218 340770 651454
rect 341006 651218 341048 651454
rect 340728 651134 341048 651218
rect 340728 650898 340770 651134
rect 341006 650898 341048 651134
rect 340728 650866 341048 650898
rect 350968 651454 351288 651486
rect 350968 651218 351010 651454
rect 351246 651218 351288 651454
rect 350968 651134 351288 651218
rect 350968 650898 351010 651134
rect 351246 650898 351288 651134
rect 350968 650866 351288 650898
rect 361208 651454 361528 651486
rect 361208 651218 361250 651454
rect 361486 651218 361528 651454
rect 361208 651134 361528 651218
rect 361208 650898 361250 651134
rect 361486 650898 361528 651134
rect 361208 650866 361528 650898
rect 371448 651454 371768 651486
rect 371448 651218 371490 651454
rect 371726 651218 371768 651454
rect 371448 651134 371768 651218
rect 371448 650898 371490 651134
rect 371726 650898 371768 651134
rect 371448 650866 371768 650898
rect 381688 651454 382008 651486
rect 381688 651218 381730 651454
rect 381966 651218 382008 651454
rect 381688 651134 382008 651218
rect 381688 650898 381730 651134
rect 381966 650898 382008 651134
rect 381688 650866 382008 650898
rect 391928 651454 392248 651486
rect 391928 651218 391970 651454
rect 392206 651218 392248 651454
rect 391928 651134 392248 651218
rect 391928 650898 391970 651134
rect 392206 650898 392248 651134
rect 391928 650866 392248 650898
rect 402168 651454 402488 651486
rect 402168 651218 402210 651454
rect 402446 651218 402488 651454
rect 402168 651134 402488 651218
rect 402168 650898 402210 651134
rect 402446 650898 402488 651134
rect 402168 650866 402488 650898
rect 412408 651454 412728 651486
rect 412408 651218 412450 651454
rect 412686 651218 412728 651454
rect 412408 651134 412728 651218
rect 412408 650898 412450 651134
rect 412686 650898 412728 651134
rect 412408 650866 412728 650898
rect 422648 651454 422968 651486
rect 422648 651218 422690 651454
rect 422926 651218 422968 651454
rect 422648 651134 422968 651218
rect 422648 650898 422690 651134
rect 422926 650898 422968 651134
rect 422648 650866 422968 650898
rect 432888 651454 433208 651486
rect 432888 651218 432930 651454
rect 433166 651218 433208 651454
rect 432888 651134 433208 651218
rect 432888 650898 432930 651134
rect 433166 650898 433208 651134
rect 432888 650866 433208 650898
rect 443128 651454 443448 651486
rect 443128 651218 443170 651454
rect 443406 651218 443448 651454
rect 443128 651134 443448 651218
rect 443128 650898 443170 651134
rect 443406 650898 443448 651134
rect 443128 650866 443448 650898
rect 453368 651454 453688 651486
rect 453368 651218 453410 651454
rect 453646 651218 453688 651454
rect 453368 651134 453688 651218
rect 453368 650898 453410 651134
rect 453646 650898 453688 651134
rect 453368 650866 453688 650898
rect 463608 651454 463928 651486
rect 463608 651218 463650 651454
rect 463886 651218 463928 651454
rect 463608 651134 463928 651218
rect 463608 650898 463650 651134
rect 463886 650898 463928 651134
rect 463608 650866 463928 650898
rect 473848 651454 474168 651486
rect 473848 651218 473890 651454
rect 474126 651218 474168 651454
rect 473848 651134 474168 651218
rect 473848 650898 473890 651134
rect 474126 650898 474168 651134
rect 473848 650866 474168 650898
rect 484088 651454 484408 651486
rect 484088 651218 484130 651454
rect 484366 651218 484408 651454
rect 484088 651134 484408 651218
rect 484088 650898 484130 651134
rect 484366 650898 484408 651134
rect 484088 650866 484408 650898
rect 494328 651454 494648 651486
rect 494328 651218 494370 651454
rect 494606 651218 494648 651454
rect 494328 651134 494648 651218
rect 494328 650898 494370 651134
rect 494606 650898 494648 651134
rect 494328 650866 494648 650898
rect 504568 651454 504888 651486
rect 504568 651218 504610 651454
rect 504846 651218 504888 651454
rect 504568 651134 504888 651218
rect 504568 650898 504610 651134
rect 504846 650898 504888 651134
rect 504568 650866 504888 650898
rect 514808 651454 515128 651486
rect 514808 651218 514850 651454
rect 515086 651218 515128 651454
rect 514808 651134 515128 651218
rect 514808 650898 514850 651134
rect 515086 650898 515128 651134
rect 514808 650866 515128 650898
rect 525048 651454 525368 651486
rect 525048 651218 525090 651454
rect 525326 651218 525368 651454
rect 525048 651134 525368 651218
rect 525048 650898 525090 651134
rect 525326 650898 525368 651134
rect 525048 650866 525368 650898
rect 535288 651454 535608 651486
rect 535288 651218 535330 651454
rect 535566 651218 535608 651454
rect 535288 651134 535608 651218
rect 535288 650898 535330 651134
rect 535566 650898 535608 651134
rect 535288 650866 535608 650898
rect 28408 633454 28728 633486
rect 28408 633218 28450 633454
rect 28686 633218 28728 633454
rect 28408 633134 28728 633218
rect 28408 632898 28450 633134
rect 28686 632898 28728 633134
rect 28408 632866 28728 632898
rect 38648 633454 38968 633486
rect 38648 633218 38690 633454
rect 38926 633218 38968 633454
rect 38648 633134 38968 633218
rect 38648 632898 38690 633134
rect 38926 632898 38968 633134
rect 38648 632866 38968 632898
rect 48888 633454 49208 633486
rect 48888 633218 48930 633454
rect 49166 633218 49208 633454
rect 48888 633134 49208 633218
rect 48888 632898 48930 633134
rect 49166 632898 49208 633134
rect 48888 632866 49208 632898
rect 59128 633454 59448 633486
rect 59128 633218 59170 633454
rect 59406 633218 59448 633454
rect 59128 633134 59448 633218
rect 59128 632898 59170 633134
rect 59406 632898 59448 633134
rect 59128 632866 59448 632898
rect 69368 633454 69688 633486
rect 69368 633218 69410 633454
rect 69646 633218 69688 633454
rect 69368 633134 69688 633218
rect 69368 632898 69410 633134
rect 69646 632898 69688 633134
rect 69368 632866 69688 632898
rect 79608 633454 79928 633486
rect 79608 633218 79650 633454
rect 79886 633218 79928 633454
rect 79608 633134 79928 633218
rect 79608 632898 79650 633134
rect 79886 632898 79928 633134
rect 79608 632866 79928 632898
rect 89848 633454 90168 633486
rect 89848 633218 89890 633454
rect 90126 633218 90168 633454
rect 89848 633134 90168 633218
rect 89848 632898 89890 633134
rect 90126 632898 90168 633134
rect 89848 632866 90168 632898
rect 100088 633454 100408 633486
rect 100088 633218 100130 633454
rect 100366 633218 100408 633454
rect 100088 633134 100408 633218
rect 100088 632898 100130 633134
rect 100366 632898 100408 633134
rect 100088 632866 100408 632898
rect 110328 633454 110648 633486
rect 110328 633218 110370 633454
rect 110606 633218 110648 633454
rect 110328 633134 110648 633218
rect 110328 632898 110370 633134
rect 110606 632898 110648 633134
rect 110328 632866 110648 632898
rect 120568 633454 120888 633486
rect 120568 633218 120610 633454
rect 120846 633218 120888 633454
rect 120568 633134 120888 633218
rect 120568 632898 120610 633134
rect 120846 632898 120888 633134
rect 120568 632866 120888 632898
rect 130808 633454 131128 633486
rect 130808 633218 130850 633454
rect 131086 633218 131128 633454
rect 130808 633134 131128 633218
rect 130808 632898 130850 633134
rect 131086 632898 131128 633134
rect 130808 632866 131128 632898
rect 141048 633454 141368 633486
rect 141048 633218 141090 633454
rect 141326 633218 141368 633454
rect 141048 633134 141368 633218
rect 141048 632898 141090 633134
rect 141326 632898 141368 633134
rect 141048 632866 141368 632898
rect 151288 633454 151608 633486
rect 151288 633218 151330 633454
rect 151566 633218 151608 633454
rect 151288 633134 151608 633218
rect 151288 632898 151330 633134
rect 151566 632898 151608 633134
rect 151288 632866 151608 632898
rect 161528 633454 161848 633486
rect 161528 633218 161570 633454
rect 161806 633218 161848 633454
rect 161528 633134 161848 633218
rect 161528 632898 161570 633134
rect 161806 632898 161848 633134
rect 161528 632866 161848 632898
rect 171768 633454 172088 633486
rect 171768 633218 171810 633454
rect 172046 633218 172088 633454
rect 171768 633134 172088 633218
rect 171768 632898 171810 633134
rect 172046 632898 172088 633134
rect 171768 632866 172088 632898
rect 182008 633454 182328 633486
rect 182008 633218 182050 633454
rect 182286 633218 182328 633454
rect 182008 633134 182328 633218
rect 182008 632898 182050 633134
rect 182286 632898 182328 633134
rect 182008 632866 182328 632898
rect 192248 633454 192568 633486
rect 192248 633218 192290 633454
rect 192526 633218 192568 633454
rect 192248 633134 192568 633218
rect 192248 632898 192290 633134
rect 192526 632898 192568 633134
rect 192248 632866 192568 632898
rect 202488 633454 202808 633486
rect 202488 633218 202530 633454
rect 202766 633218 202808 633454
rect 202488 633134 202808 633218
rect 202488 632898 202530 633134
rect 202766 632898 202808 633134
rect 202488 632866 202808 632898
rect 212728 633454 213048 633486
rect 212728 633218 212770 633454
rect 213006 633218 213048 633454
rect 212728 633134 213048 633218
rect 212728 632898 212770 633134
rect 213006 632898 213048 633134
rect 212728 632866 213048 632898
rect 222968 633454 223288 633486
rect 222968 633218 223010 633454
rect 223246 633218 223288 633454
rect 222968 633134 223288 633218
rect 222968 632898 223010 633134
rect 223246 632898 223288 633134
rect 222968 632866 223288 632898
rect 233208 633454 233528 633486
rect 233208 633218 233250 633454
rect 233486 633218 233528 633454
rect 233208 633134 233528 633218
rect 233208 632898 233250 633134
rect 233486 632898 233528 633134
rect 233208 632866 233528 632898
rect 243448 633454 243768 633486
rect 243448 633218 243490 633454
rect 243726 633218 243768 633454
rect 243448 633134 243768 633218
rect 243448 632898 243490 633134
rect 243726 632898 243768 633134
rect 243448 632866 243768 632898
rect 253688 633454 254008 633486
rect 253688 633218 253730 633454
rect 253966 633218 254008 633454
rect 253688 633134 254008 633218
rect 253688 632898 253730 633134
rect 253966 632898 254008 633134
rect 253688 632866 254008 632898
rect 263928 633454 264248 633486
rect 263928 633218 263970 633454
rect 264206 633218 264248 633454
rect 263928 633134 264248 633218
rect 263928 632898 263970 633134
rect 264206 632898 264248 633134
rect 263928 632866 264248 632898
rect 274168 633454 274488 633486
rect 274168 633218 274210 633454
rect 274446 633218 274488 633454
rect 274168 633134 274488 633218
rect 274168 632898 274210 633134
rect 274446 632898 274488 633134
rect 274168 632866 274488 632898
rect 284408 633454 284728 633486
rect 284408 633218 284450 633454
rect 284686 633218 284728 633454
rect 284408 633134 284728 633218
rect 284408 632898 284450 633134
rect 284686 632898 284728 633134
rect 284408 632866 284728 632898
rect 294648 633454 294968 633486
rect 294648 633218 294690 633454
rect 294926 633218 294968 633454
rect 294648 633134 294968 633218
rect 294648 632898 294690 633134
rect 294926 632898 294968 633134
rect 294648 632866 294968 632898
rect 304888 633454 305208 633486
rect 304888 633218 304930 633454
rect 305166 633218 305208 633454
rect 304888 633134 305208 633218
rect 304888 632898 304930 633134
rect 305166 632898 305208 633134
rect 304888 632866 305208 632898
rect 315128 633454 315448 633486
rect 315128 633218 315170 633454
rect 315406 633218 315448 633454
rect 315128 633134 315448 633218
rect 315128 632898 315170 633134
rect 315406 632898 315448 633134
rect 315128 632866 315448 632898
rect 325368 633454 325688 633486
rect 325368 633218 325410 633454
rect 325646 633218 325688 633454
rect 325368 633134 325688 633218
rect 325368 632898 325410 633134
rect 325646 632898 325688 633134
rect 325368 632866 325688 632898
rect 335608 633454 335928 633486
rect 335608 633218 335650 633454
rect 335886 633218 335928 633454
rect 335608 633134 335928 633218
rect 335608 632898 335650 633134
rect 335886 632898 335928 633134
rect 335608 632866 335928 632898
rect 345848 633454 346168 633486
rect 345848 633218 345890 633454
rect 346126 633218 346168 633454
rect 345848 633134 346168 633218
rect 345848 632898 345890 633134
rect 346126 632898 346168 633134
rect 345848 632866 346168 632898
rect 356088 633454 356408 633486
rect 356088 633218 356130 633454
rect 356366 633218 356408 633454
rect 356088 633134 356408 633218
rect 356088 632898 356130 633134
rect 356366 632898 356408 633134
rect 356088 632866 356408 632898
rect 366328 633454 366648 633486
rect 366328 633218 366370 633454
rect 366606 633218 366648 633454
rect 366328 633134 366648 633218
rect 366328 632898 366370 633134
rect 366606 632898 366648 633134
rect 366328 632866 366648 632898
rect 376568 633454 376888 633486
rect 376568 633218 376610 633454
rect 376846 633218 376888 633454
rect 376568 633134 376888 633218
rect 376568 632898 376610 633134
rect 376846 632898 376888 633134
rect 376568 632866 376888 632898
rect 386808 633454 387128 633486
rect 386808 633218 386850 633454
rect 387086 633218 387128 633454
rect 386808 633134 387128 633218
rect 386808 632898 386850 633134
rect 387086 632898 387128 633134
rect 386808 632866 387128 632898
rect 397048 633454 397368 633486
rect 397048 633218 397090 633454
rect 397326 633218 397368 633454
rect 397048 633134 397368 633218
rect 397048 632898 397090 633134
rect 397326 632898 397368 633134
rect 397048 632866 397368 632898
rect 407288 633454 407608 633486
rect 407288 633218 407330 633454
rect 407566 633218 407608 633454
rect 407288 633134 407608 633218
rect 407288 632898 407330 633134
rect 407566 632898 407608 633134
rect 407288 632866 407608 632898
rect 417528 633454 417848 633486
rect 417528 633218 417570 633454
rect 417806 633218 417848 633454
rect 417528 633134 417848 633218
rect 417528 632898 417570 633134
rect 417806 632898 417848 633134
rect 417528 632866 417848 632898
rect 427768 633454 428088 633486
rect 427768 633218 427810 633454
rect 428046 633218 428088 633454
rect 427768 633134 428088 633218
rect 427768 632898 427810 633134
rect 428046 632898 428088 633134
rect 427768 632866 428088 632898
rect 438008 633454 438328 633486
rect 438008 633218 438050 633454
rect 438286 633218 438328 633454
rect 438008 633134 438328 633218
rect 438008 632898 438050 633134
rect 438286 632898 438328 633134
rect 438008 632866 438328 632898
rect 448248 633454 448568 633486
rect 448248 633218 448290 633454
rect 448526 633218 448568 633454
rect 448248 633134 448568 633218
rect 448248 632898 448290 633134
rect 448526 632898 448568 633134
rect 448248 632866 448568 632898
rect 458488 633454 458808 633486
rect 458488 633218 458530 633454
rect 458766 633218 458808 633454
rect 458488 633134 458808 633218
rect 458488 632898 458530 633134
rect 458766 632898 458808 633134
rect 458488 632866 458808 632898
rect 468728 633454 469048 633486
rect 468728 633218 468770 633454
rect 469006 633218 469048 633454
rect 468728 633134 469048 633218
rect 468728 632898 468770 633134
rect 469006 632898 469048 633134
rect 468728 632866 469048 632898
rect 478968 633454 479288 633486
rect 478968 633218 479010 633454
rect 479246 633218 479288 633454
rect 478968 633134 479288 633218
rect 478968 632898 479010 633134
rect 479246 632898 479288 633134
rect 478968 632866 479288 632898
rect 489208 633454 489528 633486
rect 489208 633218 489250 633454
rect 489486 633218 489528 633454
rect 489208 633134 489528 633218
rect 489208 632898 489250 633134
rect 489486 632898 489528 633134
rect 489208 632866 489528 632898
rect 499448 633454 499768 633486
rect 499448 633218 499490 633454
rect 499726 633218 499768 633454
rect 499448 633134 499768 633218
rect 499448 632898 499490 633134
rect 499726 632898 499768 633134
rect 499448 632866 499768 632898
rect 509688 633454 510008 633486
rect 509688 633218 509730 633454
rect 509966 633218 510008 633454
rect 509688 633134 510008 633218
rect 509688 632898 509730 633134
rect 509966 632898 510008 633134
rect 509688 632866 510008 632898
rect 519928 633454 520248 633486
rect 519928 633218 519970 633454
rect 520206 633218 520248 633454
rect 519928 633134 520248 633218
rect 519928 632898 519970 633134
rect 520206 632898 520248 633134
rect 519928 632866 520248 632898
rect 530168 633454 530488 633486
rect 530168 633218 530210 633454
rect 530446 633218 530488 633454
rect 530168 633134 530488 633218
rect 530168 632898 530210 633134
rect 530446 632898 530488 633134
rect 530168 632866 530488 632898
rect 15754 618938 15786 619174
rect 16022 618938 16106 619174
rect 16342 618938 16374 619174
rect 15754 618854 16374 618938
rect 15754 618618 15786 618854
rect 16022 618618 16106 618854
rect 16342 618618 16374 618854
rect 15754 583174 16374 618618
rect 541714 622894 542334 658338
rect 541714 622658 541746 622894
rect 541982 622658 542066 622894
rect 542302 622658 542334 622894
rect 541714 622574 542334 622658
rect 541714 622338 541746 622574
rect 541982 622338 542066 622574
rect 542302 622338 542334 622574
rect 23288 615454 23608 615486
rect 23288 615218 23330 615454
rect 23566 615218 23608 615454
rect 23288 615134 23608 615218
rect 23288 614898 23330 615134
rect 23566 614898 23608 615134
rect 23288 614866 23608 614898
rect 33528 615454 33848 615486
rect 33528 615218 33570 615454
rect 33806 615218 33848 615454
rect 33528 615134 33848 615218
rect 33528 614898 33570 615134
rect 33806 614898 33848 615134
rect 33528 614866 33848 614898
rect 43768 615454 44088 615486
rect 43768 615218 43810 615454
rect 44046 615218 44088 615454
rect 43768 615134 44088 615218
rect 43768 614898 43810 615134
rect 44046 614898 44088 615134
rect 43768 614866 44088 614898
rect 54008 615454 54328 615486
rect 54008 615218 54050 615454
rect 54286 615218 54328 615454
rect 54008 615134 54328 615218
rect 54008 614898 54050 615134
rect 54286 614898 54328 615134
rect 54008 614866 54328 614898
rect 64248 615454 64568 615486
rect 64248 615218 64290 615454
rect 64526 615218 64568 615454
rect 64248 615134 64568 615218
rect 64248 614898 64290 615134
rect 64526 614898 64568 615134
rect 64248 614866 64568 614898
rect 74488 615454 74808 615486
rect 74488 615218 74530 615454
rect 74766 615218 74808 615454
rect 74488 615134 74808 615218
rect 74488 614898 74530 615134
rect 74766 614898 74808 615134
rect 74488 614866 74808 614898
rect 84728 615454 85048 615486
rect 84728 615218 84770 615454
rect 85006 615218 85048 615454
rect 84728 615134 85048 615218
rect 84728 614898 84770 615134
rect 85006 614898 85048 615134
rect 84728 614866 85048 614898
rect 94968 615454 95288 615486
rect 94968 615218 95010 615454
rect 95246 615218 95288 615454
rect 94968 615134 95288 615218
rect 94968 614898 95010 615134
rect 95246 614898 95288 615134
rect 94968 614866 95288 614898
rect 105208 615454 105528 615486
rect 105208 615218 105250 615454
rect 105486 615218 105528 615454
rect 105208 615134 105528 615218
rect 105208 614898 105250 615134
rect 105486 614898 105528 615134
rect 105208 614866 105528 614898
rect 115448 615454 115768 615486
rect 115448 615218 115490 615454
rect 115726 615218 115768 615454
rect 115448 615134 115768 615218
rect 115448 614898 115490 615134
rect 115726 614898 115768 615134
rect 115448 614866 115768 614898
rect 125688 615454 126008 615486
rect 125688 615218 125730 615454
rect 125966 615218 126008 615454
rect 125688 615134 126008 615218
rect 125688 614898 125730 615134
rect 125966 614898 126008 615134
rect 125688 614866 126008 614898
rect 135928 615454 136248 615486
rect 135928 615218 135970 615454
rect 136206 615218 136248 615454
rect 135928 615134 136248 615218
rect 135928 614898 135970 615134
rect 136206 614898 136248 615134
rect 135928 614866 136248 614898
rect 146168 615454 146488 615486
rect 146168 615218 146210 615454
rect 146446 615218 146488 615454
rect 146168 615134 146488 615218
rect 146168 614898 146210 615134
rect 146446 614898 146488 615134
rect 146168 614866 146488 614898
rect 156408 615454 156728 615486
rect 156408 615218 156450 615454
rect 156686 615218 156728 615454
rect 156408 615134 156728 615218
rect 156408 614898 156450 615134
rect 156686 614898 156728 615134
rect 156408 614866 156728 614898
rect 166648 615454 166968 615486
rect 166648 615218 166690 615454
rect 166926 615218 166968 615454
rect 166648 615134 166968 615218
rect 166648 614898 166690 615134
rect 166926 614898 166968 615134
rect 166648 614866 166968 614898
rect 176888 615454 177208 615486
rect 176888 615218 176930 615454
rect 177166 615218 177208 615454
rect 176888 615134 177208 615218
rect 176888 614898 176930 615134
rect 177166 614898 177208 615134
rect 176888 614866 177208 614898
rect 187128 615454 187448 615486
rect 187128 615218 187170 615454
rect 187406 615218 187448 615454
rect 187128 615134 187448 615218
rect 187128 614898 187170 615134
rect 187406 614898 187448 615134
rect 187128 614866 187448 614898
rect 197368 615454 197688 615486
rect 197368 615218 197410 615454
rect 197646 615218 197688 615454
rect 197368 615134 197688 615218
rect 197368 614898 197410 615134
rect 197646 614898 197688 615134
rect 197368 614866 197688 614898
rect 207608 615454 207928 615486
rect 207608 615218 207650 615454
rect 207886 615218 207928 615454
rect 207608 615134 207928 615218
rect 207608 614898 207650 615134
rect 207886 614898 207928 615134
rect 207608 614866 207928 614898
rect 217848 615454 218168 615486
rect 217848 615218 217890 615454
rect 218126 615218 218168 615454
rect 217848 615134 218168 615218
rect 217848 614898 217890 615134
rect 218126 614898 218168 615134
rect 217848 614866 218168 614898
rect 228088 615454 228408 615486
rect 228088 615218 228130 615454
rect 228366 615218 228408 615454
rect 228088 615134 228408 615218
rect 228088 614898 228130 615134
rect 228366 614898 228408 615134
rect 228088 614866 228408 614898
rect 238328 615454 238648 615486
rect 238328 615218 238370 615454
rect 238606 615218 238648 615454
rect 238328 615134 238648 615218
rect 238328 614898 238370 615134
rect 238606 614898 238648 615134
rect 238328 614866 238648 614898
rect 248568 615454 248888 615486
rect 248568 615218 248610 615454
rect 248846 615218 248888 615454
rect 248568 615134 248888 615218
rect 248568 614898 248610 615134
rect 248846 614898 248888 615134
rect 248568 614866 248888 614898
rect 258808 615454 259128 615486
rect 258808 615218 258850 615454
rect 259086 615218 259128 615454
rect 258808 615134 259128 615218
rect 258808 614898 258850 615134
rect 259086 614898 259128 615134
rect 258808 614866 259128 614898
rect 269048 615454 269368 615486
rect 269048 615218 269090 615454
rect 269326 615218 269368 615454
rect 269048 615134 269368 615218
rect 269048 614898 269090 615134
rect 269326 614898 269368 615134
rect 269048 614866 269368 614898
rect 279288 615454 279608 615486
rect 279288 615218 279330 615454
rect 279566 615218 279608 615454
rect 279288 615134 279608 615218
rect 279288 614898 279330 615134
rect 279566 614898 279608 615134
rect 279288 614866 279608 614898
rect 289528 615454 289848 615486
rect 289528 615218 289570 615454
rect 289806 615218 289848 615454
rect 289528 615134 289848 615218
rect 289528 614898 289570 615134
rect 289806 614898 289848 615134
rect 289528 614866 289848 614898
rect 299768 615454 300088 615486
rect 299768 615218 299810 615454
rect 300046 615218 300088 615454
rect 299768 615134 300088 615218
rect 299768 614898 299810 615134
rect 300046 614898 300088 615134
rect 299768 614866 300088 614898
rect 310008 615454 310328 615486
rect 310008 615218 310050 615454
rect 310286 615218 310328 615454
rect 310008 615134 310328 615218
rect 310008 614898 310050 615134
rect 310286 614898 310328 615134
rect 310008 614866 310328 614898
rect 320248 615454 320568 615486
rect 320248 615218 320290 615454
rect 320526 615218 320568 615454
rect 320248 615134 320568 615218
rect 320248 614898 320290 615134
rect 320526 614898 320568 615134
rect 320248 614866 320568 614898
rect 330488 615454 330808 615486
rect 330488 615218 330530 615454
rect 330766 615218 330808 615454
rect 330488 615134 330808 615218
rect 330488 614898 330530 615134
rect 330766 614898 330808 615134
rect 330488 614866 330808 614898
rect 340728 615454 341048 615486
rect 340728 615218 340770 615454
rect 341006 615218 341048 615454
rect 340728 615134 341048 615218
rect 340728 614898 340770 615134
rect 341006 614898 341048 615134
rect 340728 614866 341048 614898
rect 350968 615454 351288 615486
rect 350968 615218 351010 615454
rect 351246 615218 351288 615454
rect 350968 615134 351288 615218
rect 350968 614898 351010 615134
rect 351246 614898 351288 615134
rect 350968 614866 351288 614898
rect 361208 615454 361528 615486
rect 361208 615218 361250 615454
rect 361486 615218 361528 615454
rect 361208 615134 361528 615218
rect 361208 614898 361250 615134
rect 361486 614898 361528 615134
rect 361208 614866 361528 614898
rect 371448 615454 371768 615486
rect 371448 615218 371490 615454
rect 371726 615218 371768 615454
rect 371448 615134 371768 615218
rect 371448 614898 371490 615134
rect 371726 614898 371768 615134
rect 371448 614866 371768 614898
rect 381688 615454 382008 615486
rect 381688 615218 381730 615454
rect 381966 615218 382008 615454
rect 381688 615134 382008 615218
rect 381688 614898 381730 615134
rect 381966 614898 382008 615134
rect 381688 614866 382008 614898
rect 391928 615454 392248 615486
rect 391928 615218 391970 615454
rect 392206 615218 392248 615454
rect 391928 615134 392248 615218
rect 391928 614898 391970 615134
rect 392206 614898 392248 615134
rect 391928 614866 392248 614898
rect 402168 615454 402488 615486
rect 402168 615218 402210 615454
rect 402446 615218 402488 615454
rect 402168 615134 402488 615218
rect 402168 614898 402210 615134
rect 402446 614898 402488 615134
rect 402168 614866 402488 614898
rect 412408 615454 412728 615486
rect 412408 615218 412450 615454
rect 412686 615218 412728 615454
rect 412408 615134 412728 615218
rect 412408 614898 412450 615134
rect 412686 614898 412728 615134
rect 412408 614866 412728 614898
rect 422648 615454 422968 615486
rect 422648 615218 422690 615454
rect 422926 615218 422968 615454
rect 422648 615134 422968 615218
rect 422648 614898 422690 615134
rect 422926 614898 422968 615134
rect 422648 614866 422968 614898
rect 432888 615454 433208 615486
rect 432888 615218 432930 615454
rect 433166 615218 433208 615454
rect 432888 615134 433208 615218
rect 432888 614898 432930 615134
rect 433166 614898 433208 615134
rect 432888 614866 433208 614898
rect 443128 615454 443448 615486
rect 443128 615218 443170 615454
rect 443406 615218 443448 615454
rect 443128 615134 443448 615218
rect 443128 614898 443170 615134
rect 443406 614898 443448 615134
rect 443128 614866 443448 614898
rect 453368 615454 453688 615486
rect 453368 615218 453410 615454
rect 453646 615218 453688 615454
rect 453368 615134 453688 615218
rect 453368 614898 453410 615134
rect 453646 614898 453688 615134
rect 453368 614866 453688 614898
rect 463608 615454 463928 615486
rect 463608 615218 463650 615454
rect 463886 615218 463928 615454
rect 463608 615134 463928 615218
rect 463608 614898 463650 615134
rect 463886 614898 463928 615134
rect 463608 614866 463928 614898
rect 473848 615454 474168 615486
rect 473848 615218 473890 615454
rect 474126 615218 474168 615454
rect 473848 615134 474168 615218
rect 473848 614898 473890 615134
rect 474126 614898 474168 615134
rect 473848 614866 474168 614898
rect 484088 615454 484408 615486
rect 484088 615218 484130 615454
rect 484366 615218 484408 615454
rect 484088 615134 484408 615218
rect 484088 614898 484130 615134
rect 484366 614898 484408 615134
rect 484088 614866 484408 614898
rect 494328 615454 494648 615486
rect 494328 615218 494370 615454
rect 494606 615218 494648 615454
rect 494328 615134 494648 615218
rect 494328 614898 494370 615134
rect 494606 614898 494648 615134
rect 494328 614866 494648 614898
rect 504568 615454 504888 615486
rect 504568 615218 504610 615454
rect 504846 615218 504888 615454
rect 504568 615134 504888 615218
rect 504568 614898 504610 615134
rect 504846 614898 504888 615134
rect 504568 614866 504888 614898
rect 514808 615454 515128 615486
rect 514808 615218 514850 615454
rect 515086 615218 515128 615454
rect 514808 615134 515128 615218
rect 514808 614898 514850 615134
rect 515086 614898 515128 615134
rect 514808 614866 515128 614898
rect 525048 615454 525368 615486
rect 525048 615218 525090 615454
rect 525326 615218 525368 615454
rect 525048 615134 525368 615218
rect 525048 614898 525090 615134
rect 525326 614898 525368 615134
rect 525048 614866 525368 614898
rect 535288 615454 535608 615486
rect 535288 615218 535330 615454
rect 535566 615218 535608 615454
rect 535288 615134 535608 615218
rect 535288 614898 535330 615134
rect 535566 614898 535608 615134
rect 535288 614866 535608 614898
rect 28408 597454 28728 597486
rect 28408 597218 28450 597454
rect 28686 597218 28728 597454
rect 28408 597134 28728 597218
rect 28408 596898 28450 597134
rect 28686 596898 28728 597134
rect 28408 596866 28728 596898
rect 38648 597454 38968 597486
rect 38648 597218 38690 597454
rect 38926 597218 38968 597454
rect 38648 597134 38968 597218
rect 38648 596898 38690 597134
rect 38926 596898 38968 597134
rect 38648 596866 38968 596898
rect 48888 597454 49208 597486
rect 48888 597218 48930 597454
rect 49166 597218 49208 597454
rect 48888 597134 49208 597218
rect 48888 596898 48930 597134
rect 49166 596898 49208 597134
rect 48888 596866 49208 596898
rect 59128 597454 59448 597486
rect 59128 597218 59170 597454
rect 59406 597218 59448 597454
rect 59128 597134 59448 597218
rect 59128 596898 59170 597134
rect 59406 596898 59448 597134
rect 59128 596866 59448 596898
rect 69368 597454 69688 597486
rect 69368 597218 69410 597454
rect 69646 597218 69688 597454
rect 69368 597134 69688 597218
rect 69368 596898 69410 597134
rect 69646 596898 69688 597134
rect 69368 596866 69688 596898
rect 79608 597454 79928 597486
rect 79608 597218 79650 597454
rect 79886 597218 79928 597454
rect 79608 597134 79928 597218
rect 79608 596898 79650 597134
rect 79886 596898 79928 597134
rect 79608 596866 79928 596898
rect 89848 597454 90168 597486
rect 89848 597218 89890 597454
rect 90126 597218 90168 597454
rect 89848 597134 90168 597218
rect 89848 596898 89890 597134
rect 90126 596898 90168 597134
rect 89848 596866 90168 596898
rect 100088 597454 100408 597486
rect 100088 597218 100130 597454
rect 100366 597218 100408 597454
rect 100088 597134 100408 597218
rect 100088 596898 100130 597134
rect 100366 596898 100408 597134
rect 100088 596866 100408 596898
rect 110328 597454 110648 597486
rect 110328 597218 110370 597454
rect 110606 597218 110648 597454
rect 110328 597134 110648 597218
rect 110328 596898 110370 597134
rect 110606 596898 110648 597134
rect 110328 596866 110648 596898
rect 120568 597454 120888 597486
rect 120568 597218 120610 597454
rect 120846 597218 120888 597454
rect 120568 597134 120888 597218
rect 120568 596898 120610 597134
rect 120846 596898 120888 597134
rect 120568 596866 120888 596898
rect 130808 597454 131128 597486
rect 130808 597218 130850 597454
rect 131086 597218 131128 597454
rect 130808 597134 131128 597218
rect 130808 596898 130850 597134
rect 131086 596898 131128 597134
rect 130808 596866 131128 596898
rect 141048 597454 141368 597486
rect 141048 597218 141090 597454
rect 141326 597218 141368 597454
rect 141048 597134 141368 597218
rect 141048 596898 141090 597134
rect 141326 596898 141368 597134
rect 141048 596866 141368 596898
rect 151288 597454 151608 597486
rect 151288 597218 151330 597454
rect 151566 597218 151608 597454
rect 151288 597134 151608 597218
rect 151288 596898 151330 597134
rect 151566 596898 151608 597134
rect 151288 596866 151608 596898
rect 161528 597454 161848 597486
rect 161528 597218 161570 597454
rect 161806 597218 161848 597454
rect 161528 597134 161848 597218
rect 161528 596898 161570 597134
rect 161806 596898 161848 597134
rect 161528 596866 161848 596898
rect 171768 597454 172088 597486
rect 171768 597218 171810 597454
rect 172046 597218 172088 597454
rect 171768 597134 172088 597218
rect 171768 596898 171810 597134
rect 172046 596898 172088 597134
rect 171768 596866 172088 596898
rect 182008 597454 182328 597486
rect 182008 597218 182050 597454
rect 182286 597218 182328 597454
rect 182008 597134 182328 597218
rect 182008 596898 182050 597134
rect 182286 596898 182328 597134
rect 182008 596866 182328 596898
rect 192248 597454 192568 597486
rect 192248 597218 192290 597454
rect 192526 597218 192568 597454
rect 192248 597134 192568 597218
rect 192248 596898 192290 597134
rect 192526 596898 192568 597134
rect 192248 596866 192568 596898
rect 202488 597454 202808 597486
rect 202488 597218 202530 597454
rect 202766 597218 202808 597454
rect 202488 597134 202808 597218
rect 202488 596898 202530 597134
rect 202766 596898 202808 597134
rect 202488 596866 202808 596898
rect 212728 597454 213048 597486
rect 212728 597218 212770 597454
rect 213006 597218 213048 597454
rect 212728 597134 213048 597218
rect 212728 596898 212770 597134
rect 213006 596898 213048 597134
rect 212728 596866 213048 596898
rect 222968 597454 223288 597486
rect 222968 597218 223010 597454
rect 223246 597218 223288 597454
rect 222968 597134 223288 597218
rect 222968 596898 223010 597134
rect 223246 596898 223288 597134
rect 222968 596866 223288 596898
rect 233208 597454 233528 597486
rect 233208 597218 233250 597454
rect 233486 597218 233528 597454
rect 233208 597134 233528 597218
rect 233208 596898 233250 597134
rect 233486 596898 233528 597134
rect 233208 596866 233528 596898
rect 243448 597454 243768 597486
rect 243448 597218 243490 597454
rect 243726 597218 243768 597454
rect 243448 597134 243768 597218
rect 243448 596898 243490 597134
rect 243726 596898 243768 597134
rect 243448 596866 243768 596898
rect 253688 597454 254008 597486
rect 253688 597218 253730 597454
rect 253966 597218 254008 597454
rect 253688 597134 254008 597218
rect 253688 596898 253730 597134
rect 253966 596898 254008 597134
rect 253688 596866 254008 596898
rect 263928 597454 264248 597486
rect 263928 597218 263970 597454
rect 264206 597218 264248 597454
rect 263928 597134 264248 597218
rect 263928 596898 263970 597134
rect 264206 596898 264248 597134
rect 263928 596866 264248 596898
rect 274168 597454 274488 597486
rect 274168 597218 274210 597454
rect 274446 597218 274488 597454
rect 274168 597134 274488 597218
rect 274168 596898 274210 597134
rect 274446 596898 274488 597134
rect 274168 596866 274488 596898
rect 284408 597454 284728 597486
rect 284408 597218 284450 597454
rect 284686 597218 284728 597454
rect 284408 597134 284728 597218
rect 284408 596898 284450 597134
rect 284686 596898 284728 597134
rect 284408 596866 284728 596898
rect 294648 597454 294968 597486
rect 294648 597218 294690 597454
rect 294926 597218 294968 597454
rect 294648 597134 294968 597218
rect 294648 596898 294690 597134
rect 294926 596898 294968 597134
rect 294648 596866 294968 596898
rect 304888 597454 305208 597486
rect 304888 597218 304930 597454
rect 305166 597218 305208 597454
rect 304888 597134 305208 597218
rect 304888 596898 304930 597134
rect 305166 596898 305208 597134
rect 304888 596866 305208 596898
rect 315128 597454 315448 597486
rect 315128 597218 315170 597454
rect 315406 597218 315448 597454
rect 315128 597134 315448 597218
rect 315128 596898 315170 597134
rect 315406 596898 315448 597134
rect 315128 596866 315448 596898
rect 325368 597454 325688 597486
rect 325368 597218 325410 597454
rect 325646 597218 325688 597454
rect 325368 597134 325688 597218
rect 325368 596898 325410 597134
rect 325646 596898 325688 597134
rect 325368 596866 325688 596898
rect 335608 597454 335928 597486
rect 335608 597218 335650 597454
rect 335886 597218 335928 597454
rect 335608 597134 335928 597218
rect 335608 596898 335650 597134
rect 335886 596898 335928 597134
rect 335608 596866 335928 596898
rect 345848 597454 346168 597486
rect 345848 597218 345890 597454
rect 346126 597218 346168 597454
rect 345848 597134 346168 597218
rect 345848 596898 345890 597134
rect 346126 596898 346168 597134
rect 345848 596866 346168 596898
rect 356088 597454 356408 597486
rect 356088 597218 356130 597454
rect 356366 597218 356408 597454
rect 356088 597134 356408 597218
rect 356088 596898 356130 597134
rect 356366 596898 356408 597134
rect 356088 596866 356408 596898
rect 366328 597454 366648 597486
rect 366328 597218 366370 597454
rect 366606 597218 366648 597454
rect 366328 597134 366648 597218
rect 366328 596898 366370 597134
rect 366606 596898 366648 597134
rect 366328 596866 366648 596898
rect 376568 597454 376888 597486
rect 376568 597218 376610 597454
rect 376846 597218 376888 597454
rect 376568 597134 376888 597218
rect 376568 596898 376610 597134
rect 376846 596898 376888 597134
rect 376568 596866 376888 596898
rect 386808 597454 387128 597486
rect 386808 597218 386850 597454
rect 387086 597218 387128 597454
rect 386808 597134 387128 597218
rect 386808 596898 386850 597134
rect 387086 596898 387128 597134
rect 386808 596866 387128 596898
rect 397048 597454 397368 597486
rect 397048 597218 397090 597454
rect 397326 597218 397368 597454
rect 397048 597134 397368 597218
rect 397048 596898 397090 597134
rect 397326 596898 397368 597134
rect 397048 596866 397368 596898
rect 407288 597454 407608 597486
rect 407288 597218 407330 597454
rect 407566 597218 407608 597454
rect 407288 597134 407608 597218
rect 407288 596898 407330 597134
rect 407566 596898 407608 597134
rect 407288 596866 407608 596898
rect 417528 597454 417848 597486
rect 417528 597218 417570 597454
rect 417806 597218 417848 597454
rect 417528 597134 417848 597218
rect 417528 596898 417570 597134
rect 417806 596898 417848 597134
rect 417528 596866 417848 596898
rect 427768 597454 428088 597486
rect 427768 597218 427810 597454
rect 428046 597218 428088 597454
rect 427768 597134 428088 597218
rect 427768 596898 427810 597134
rect 428046 596898 428088 597134
rect 427768 596866 428088 596898
rect 438008 597454 438328 597486
rect 438008 597218 438050 597454
rect 438286 597218 438328 597454
rect 438008 597134 438328 597218
rect 438008 596898 438050 597134
rect 438286 596898 438328 597134
rect 438008 596866 438328 596898
rect 448248 597454 448568 597486
rect 448248 597218 448290 597454
rect 448526 597218 448568 597454
rect 448248 597134 448568 597218
rect 448248 596898 448290 597134
rect 448526 596898 448568 597134
rect 448248 596866 448568 596898
rect 458488 597454 458808 597486
rect 458488 597218 458530 597454
rect 458766 597218 458808 597454
rect 458488 597134 458808 597218
rect 458488 596898 458530 597134
rect 458766 596898 458808 597134
rect 458488 596866 458808 596898
rect 468728 597454 469048 597486
rect 468728 597218 468770 597454
rect 469006 597218 469048 597454
rect 468728 597134 469048 597218
rect 468728 596898 468770 597134
rect 469006 596898 469048 597134
rect 468728 596866 469048 596898
rect 478968 597454 479288 597486
rect 478968 597218 479010 597454
rect 479246 597218 479288 597454
rect 478968 597134 479288 597218
rect 478968 596898 479010 597134
rect 479246 596898 479288 597134
rect 478968 596866 479288 596898
rect 489208 597454 489528 597486
rect 489208 597218 489250 597454
rect 489486 597218 489528 597454
rect 489208 597134 489528 597218
rect 489208 596898 489250 597134
rect 489486 596898 489528 597134
rect 489208 596866 489528 596898
rect 499448 597454 499768 597486
rect 499448 597218 499490 597454
rect 499726 597218 499768 597454
rect 499448 597134 499768 597218
rect 499448 596898 499490 597134
rect 499726 596898 499768 597134
rect 499448 596866 499768 596898
rect 509688 597454 510008 597486
rect 509688 597218 509730 597454
rect 509966 597218 510008 597454
rect 509688 597134 510008 597218
rect 509688 596898 509730 597134
rect 509966 596898 510008 597134
rect 509688 596866 510008 596898
rect 519928 597454 520248 597486
rect 519928 597218 519970 597454
rect 520206 597218 520248 597454
rect 519928 597134 520248 597218
rect 519928 596898 519970 597134
rect 520206 596898 520248 597134
rect 519928 596866 520248 596898
rect 530168 597454 530488 597486
rect 530168 597218 530210 597454
rect 530446 597218 530488 597454
rect 530168 597134 530488 597218
rect 530168 596898 530210 597134
rect 530446 596898 530488 597134
rect 530168 596866 530488 596898
rect 15754 582938 15786 583174
rect 16022 582938 16106 583174
rect 16342 582938 16374 583174
rect 15754 582854 16374 582938
rect 15754 582618 15786 582854
rect 16022 582618 16106 582854
rect 16342 582618 16374 582854
rect 15754 547174 16374 582618
rect 541714 586894 542334 622338
rect 541714 586658 541746 586894
rect 541982 586658 542066 586894
rect 542302 586658 542334 586894
rect 541714 586574 542334 586658
rect 541714 586338 541746 586574
rect 541982 586338 542066 586574
rect 542302 586338 542334 586574
rect 23288 579454 23608 579486
rect 23288 579218 23330 579454
rect 23566 579218 23608 579454
rect 23288 579134 23608 579218
rect 23288 578898 23330 579134
rect 23566 578898 23608 579134
rect 23288 578866 23608 578898
rect 33528 579454 33848 579486
rect 33528 579218 33570 579454
rect 33806 579218 33848 579454
rect 33528 579134 33848 579218
rect 33528 578898 33570 579134
rect 33806 578898 33848 579134
rect 33528 578866 33848 578898
rect 43768 579454 44088 579486
rect 43768 579218 43810 579454
rect 44046 579218 44088 579454
rect 43768 579134 44088 579218
rect 43768 578898 43810 579134
rect 44046 578898 44088 579134
rect 43768 578866 44088 578898
rect 54008 579454 54328 579486
rect 54008 579218 54050 579454
rect 54286 579218 54328 579454
rect 54008 579134 54328 579218
rect 54008 578898 54050 579134
rect 54286 578898 54328 579134
rect 54008 578866 54328 578898
rect 64248 579454 64568 579486
rect 64248 579218 64290 579454
rect 64526 579218 64568 579454
rect 64248 579134 64568 579218
rect 64248 578898 64290 579134
rect 64526 578898 64568 579134
rect 64248 578866 64568 578898
rect 74488 579454 74808 579486
rect 74488 579218 74530 579454
rect 74766 579218 74808 579454
rect 74488 579134 74808 579218
rect 74488 578898 74530 579134
rect 74766 578898 74808 579134
rect 74488 578866 74808 578898
rect 84728 579454 85048 579486
rect 84728 579218 84770 579454
rect 85006 579218 85048 579454
rect 84728 579134 85048 579218
rect 84728 578898 84770 579134
rect 85006 578898 85048 579134
rect 84728 578866 85048 578898
rect 94968 579454 95288 579486
rect 94968 579218 95010 579454
rect 95246 579218 95288 579454
rect 94968 579134 95288 579218
rect 94968 578898 95010 579134
rect 95246 578898 95288 579134
rect 94968 578866 95288 578898
rect 105208 579454 105528 579486
rect 105208 579218 105250 579454
rect 105486 579218 105528 579454
rect 105208 579134 105528 579218
rect 105208 578898 105250 579134
rect 105486 578898 105528 579134
rect 105208 578866 105528 578898
rect 115448 579454 115768 579486
rect 115448 579218 115490 579454
rect 115726 579218 115768 579454
rect 115448 579134 115768 579218
rect 115448 578898 115490 579134
rect 115726 578898 115768 579134
rect 115448 578866 115768 578898
rect 125688 579454 126008 579486
rect 125688 579218 125730 579454
rect 125966 579218 126008 579454
rect 125688 579134 126008 579218
rect 125688 578898 125730 579134
rect 125966 578898 126008 579134
rect 125688 578866 126008 578898
rect 135928 579454 136248 579486
rect 135928 579218 135970 579454
rect 136206 579218 136248 579454
rect 135928 579134 136248 579218
rect 135928 578898 135970 579134
rect 136206 578898 136248 579134
rect 135928 578866 136248 578898
rect 146168 579454 146488 579486
rect 146168 579218 146210 579454
rect 146446 579218 146488 579454
rect 146168 579134 146488 579218
rect 146168 578898 146210 579134
rect 146446 578898 146488 579134
rect 146168 578866 146488 578898
rect 156408 579454 156728 579486
rect 156408 579218 156450 579454
rect 156686 579218 156728 579454
rect 156408 579134 156728 579218
rect 156408 578898 156450 579134
rect 156686 578898 156728 579134
rect 156408 578866 156728 578898
rect 166648 579454 166968 579486
rect 166648 579218 166690 579454
rect 166926 579218 166968 579454
rect 166648 579134 166968 579218
rect 166648 578898 166690 579134
rect 166926 578898 166968 579134
rect 166648 578866 166968 578898
rect 176888 579454 177208 579486
rect 176888 579218 176930 579454
rect 177166 579218 177208 579454
rect 176888 579134 177208 579218
rect 176888 578898 176930 579134
rect 177166 578898 177208 579134
rect 176888 578866 177208 578898
rect 187128 579454 187448 579486
rect 187128 579218 187170 579454
rect 187406 579218 187448 579454
rect 187128 579134 187448 579218
rect 187128 578898 187170 579134
rect 187406 578898 187448 579134
rect 187128 578866 187448 578898
rect 197368 579454 197688 579486
rect 197368 579218 197410 579454
rect 197646 579218 197688 579454
rect 197368 579134 197688 579218
rect 197368 578898 197410 579134
rect 197646 578898 197688 579134
rect 197368 578866 197688 578898
rect 207608 579454 207928 579486
rect 207608 579218 207650 579454
rect 207886 579218 207928 579454
rect 207608 579134 207928 579218
rect 207608 578898 207650 579134
rect 207886 578898 207928 579134
rect 207608 578866 207928 578898
rect 217848 579454 218168 579486
rect 217848 579218 217890 579454
rect 218126 579218 218168 579454
rect 217848 579134 218168 579218
rect 217848 578898 217890 579134
rect 218126 578898 218168 579134
rect 217848 578866 218168 578898
rect 228088 579454 228408 579486
rect 228088 579218 228130 579454
rect 228366 579218 228408 579454
rect 228088 579134 228408 579218
rect 228088 578898 228130 579134
rect 228366 578898 228408 579134
rect 228088 578866 228408 578898
rect 238328 579454 238648 579486
rect 238328 579218 238370 579454
rect 238606 579218 238648 579454
rect 238328 579134 238648 579218
rect 238328 578898 238370 579134
rect 238606 578898 238648 579134
rect 238328 578866 238648 578898
rect 248568 579454 248888 579486
rect 248568 579218 248610 579454
rect 248846 579218 248888 579454
rect 248568 579134 248888 579218
rect 248568 578898 248610 579134
rect 248846 578898 248888 579134
rect 248568 578866 248888 578898
rect 258808 579454 259128 579486
rect 258808 579218 258850 579454
rect 259086 579218 259128 579454
rect 258808 579134 259128 579218
rect 258808 578898 258850 579134
rect 259086 578898 259128 579134
rect 258808 578866 259128 578898
rect 269048 579454 269368 579486
rect 269048 579218 269090 579454
rect 269326 579218 269368 579454
rect 269048 579134 269368 579218
rect 269048 578898 269090 579134
rect 269326 578898 269368 579134
rect 269048 578866 269368 578898
rect 279288 579454 279608 579486
rect 279288 579218 279330 579454
rect 279566 579218 279608 579454
rect 279288 579134 279608 579218
rect 279288 578898 279330 579134
rect 279566 578898 279608 579134
rect 279288 578866 279608 578898
rect 289528 579454 289848 579486
rect 289528 579218 289570 579454
rect 289806 579218 289848 579454
rect 289528 579134 289848 579218
rect 289528 578898 289570 579134
rect 289806 578898 289848 579134
rect 289528 578866 289848 578898
rect 299768 579454 300088 579486
rect 299768 579218 299810 579454
rect 300046 579218 300088 579454
rect 299768 579134 300088 579218
rect 299768 578898 299810 579134
rect 300046 578898 300088 579134
rect 299768 578866 300088 578898
rect 310008 579454 310328 579486
rect 310008 579218 310050 579454
rect 310286 579218 310328 579454
rect 310008 579134 310328 579218
rect 310008 578898 310050 579134
rect 310286 578898 310328 579134
rect 310008 578866 310328 578898
rect 320248 579454 320568 579486
rect 320248 579218 320290 579454
rect 320526 579218 320568 579454
rect 320248 579134 320568 579218
rect 320248 578898 320290 579134
rect 320526 578898 320568 579134
rect 320248 578866 320568 578898
rect 330488 579454 330808 579486
rect 330488 579218 330530 579454
rect 330766 579218 330808 579454
rect 330488 579134 330808 579218
rect 330488 578898 330530 579134
rect 330766 578898 330808 579134
rect 330488 578866 330808 578898
rect 340728 579454 341048 579486
rect 340728 579218 340770 579454
rect 341006 579218 341048 579454
rect 340728 579134 341048 579218
rect 340728 578898 340770 579134
rect 341006 578898 341048 579134
rect 340728 578866 341048 578898
rect 350968 579454 351288 579486
rect 350968 579218 351010 579454
rect 351246 579218 351288 579454
rect 350968 579134 351288 579218
rect 350968 578898 351010 579134
rect 351246 578898 351288 579134
rect 350968 578866 351288 578898
rect 361208 579454 361528 579486
rect 361208 579218 361250 579454
rect 361486 579218 361528 579454
rect 361208 579134 361528 579218
rect 361208 578898 361250 579134
rect 361486 578898 361528 579134
rect 361208 578866 361528 578898
rect 371448 579454 371768 579486
rect 371448 579218 371490 579454
rect 371726 579218 371768 579454
rect 371448 579134 371768 579218
rect 371448 578898 371490 579134
rect 371726 578898 371768 579134
rect 371448 578866 371768 578898
rect 381688 579454 382008 579486
rect 381688 579218 381730 579454
rect 381966 579218 382008 579454
rect 381688 579134 382008 579218
rect 381688 578898 381730 579134
rect 381966 578898 382008 579134
rect 381688 578866 382008 578898
rect 391928 579454 392248 579486
rect 391928 579218 391970 579454
rect 392206 579218 392248 579454
rect 391928 579134 392248 579218
rect 391928 578898 391970 579134
rect 392206 578898 392248 579134
rect 391928 578866 392248 578898
rect 402168 579454 402488 579486
rect 402168 579218 402210 579454
rect 402446 579218 402488 579454
rect 402168 579134 402488 579218
rect 402168 578898 402210 579134
rect 402446 578898 402488 579134
rect 402168 578866 402488 578898
rect 412408 579454 412728 579486
rect 412408 579218 412450 579454
rect 412686 579218 412728 579454
rect 412408 579134 412728 579218
rect 412408 578898 412450 579134
rect 412686 578898 412728 579134
rect 412408 578866 412728 578898
rect 422648 579454 422968 579486
rect 422648 579218 422690 579454
rect 422926 579218 422968 579454
rect 422648 579134 422968 579218
rect 422648 578898 422690 579134
rect 422926 578898 422968 579134
rect 422648 578866 422968 578898
rect 432888 579454 433208 579486
rect 432888 579218 432930 579454
rect 433166 579218 433208 579454
rect 432888 579134 433208 579218
rect 432888 578898 432930 579134
rect 433166 578898 433208 579134
rect 432888 578866 433208 578898
rect 443128 579454 443448 579486
rect 443128 579218 443170 579454
rect 443406 579218 443448 579454
rect 443128 579134 443448 579218
rect 443128 578898 443170 579134
rect 443406 578898 443448 579134
rect 443128 578866 443448 578898
rect 453368 579454 453688 579486
rect 453368 579218 453410 579454
rect 453646 579218 453688 579454
rect 453368 579134 453688 579218
rect 453368 578898 453410 579134
rect 453646 578898 453688 579134
rect 453368 578866 453688 578898
rect 463608 579454 463928 579486
rect 463608 579218 463650 579454
rect 463886 579218 463928 579454
rect 463608 579134 463928 579218
rect 463608 578898 463650 579134
rect 463886 578898 463928 579134
rect 463608 578866 463928 578898
rect 473848 579454 474168 579486
rect 473848 579218 473890 579454
rect 474126 579218 474168 579454
rect 473848 579134 474168 579218
rect 473848 578898 473890 579134
rect 474126 578898 474168 579134
rect 473848 578866 474168 578898
rect 484088 579454 484408 579486
rect 484088 579218 484130 579454
rect 484366 579218 484408 579454
rect 484088 579134 484408 579218
rect 484088 578898 484130 579134
rect 484366 578898 484408 579134
rect 484088 578866 484408 578898
rect 494328 579454 494648 579486
rect 494328 579218 494370 579454
rect 494606 579218 494648 579454
rect 494328 579134 494648 579218
rect 494328 578898 494370 579134
rect 494606 578898 494648 579134
rect 494328 578866 494648 578898
rect 504568 579454 504888 579486
rect 504568 579218 504610 579454
rect 504846 579218 504888 579454
rect 504568 579134 504888 579218
rect 504568 578898 504610 579134
rect 504846 578898 504888 579134
rect 504568 578866 504888 578898
rect 514808 579454 515128 579486
rect 514808 579218 514850 579454
rect 515086 579218 515128 579454
rect 514808 579134 515128 579218
rect 514808 578898 514850 579134
rect 515086 578898 515128 579134
rect 514808 578866 515128 578898
rect 525048 579454 525368 579486
rect 525048 579218 525090 579454
rect 525326 579218 525368 579454
rect 525048 579134 525368 579218
rect 525048 578898 525090 579134
rect 525326 578898 525368 579134
rect 525048 578866 525368 578898
rect 535288 579454 535608 579486
rect 535288 579218 535330 579454
rect 535566 579218 535608 579454
rect 535288 579134 535608 579218
rect 535288 578898 535330 579134
rect 535566 578898 535608 579134
rect 535288 578866 535608 578898
rect 28408 561454 28728 561486
rect 28408 561218 28450 561454
rect 28686 561218 28728 561454
rect 28408 561134 28728 561218
rect 28408 560898 28450 561134
rect 28686 560898 28728 561134
rect 28408 560866 28728 560898
rect 38648 561454 38968 561486
rect 38648 561218 38690 561454
rect 38926 561218 38968 561454
rect 38648 561134 38968 561218
rect 38648 560898 38690 561134
rect 38926 560898 38968 561134
rect 38648 560866 38968 560898
rect 48888 561454 49208 561486
rect 48888 561218 48930 561454
rect 49166 561218 49208 561454
rect 48888 561134 49208 561218
rect 48888 560898 48930 561134
rect 49166 560898 49208 561134
rect 48888 560866 49208 560898
rect 59128 561454 59448 561486
rect 59128 561218 59170 561454
rect 59406 561218 59448 561454
rect 59128 561134 59448 561218
rect 59128 560898 59170 561134
rect 59406 560898 59448 561134
rect 59128 560866 59448 560898
rect 69368 561454 69688 561486
rect 69368 561218 69410 561454
rect 69646 561218 69688 561454
rect 69368 561134 69688 561218
rect 69368 560898 69410 561134
rect 69646 560898 69688 561134
rect 69368 560866 69688 560898
rect 79608 561454 79928 561486
rect 79608 561218 79650 561454
rect 79886 561218 79928 561454
rect 79608 561134 79928 561218
rect 79608 560898 79650 561134
rect 79886 560898 79928 561134
rect 79608 560866 79928 560898
rect 89848 561454 90168 561486
rect 89848 561218 89890 561454
rect 90126 561218 90168 561454
rect 89848 561134 90168 561218
rect 89848 560898 89890 561134
rect 90126 560898 90168 561134
rect 89848 560866 90168 560898
rect 100088 561454 100408 561486
rect 100088 561218 100130 561454
rect 100366 561218 100408 561454
rect 100088 561134 100408 561218
rect 100088 560898 100130 561134
rect 100366 560898 100408 561134
rect 100088 560866 100408 560898
rect 110328 561454 110648 561486
rect 110328 561218 110370 561454
rect 110606 561218 110648 561454
rect 110328 561134 110648 561218
rect 110328 560898 110370 561134
rect 110606 560898 110648 561134
rect 110328 560866 110648 560898
rect 120568 561454 120888 561486
rect 120568 561218 120610 561454
rect 120846 561218 120888 561454
rect 120568 561134 120888 561218
rect 120568 560898 120610 561134
rect 120846 560898 120888 561134
rect 120568 560866 120888 560898
rect 130808 561454 131128 561486
rect 130808 561218 130850 561454
rect 131086 561218 131128 561454
rect 130808 561134 131128 561218
rect 130808 560898 130850 561134
rect 131086 560898 131128 561134
rect 130808 560866 131128 560898
rect 141048 561454 141368 561486
rect 141048 561218 141090 561454
rect 141326 561218 141368 561454
rect 141048 561134 141368 561218
rect 141048 560898 141090 561134
rect 141326 560898 141368 561134
rect 141048 560866 141368 560898
rect 151288 561454 151608 561486
rect 151288 561218 151330 561454
rect 151566 561218 151608 561454
rect 151288 561134 151608 561218
rect 151288 560898 151330 561134
rect 151566 560898 151608 561134
rect 151288 560866 151608 560898
rect 161528 561454 161848 561486
rect 161528 561218 161570 561454
rect 161806 561218 161848 561454
rect 161528 561134 161848 561218
rect 161528 560898 161570 561134
rect 161806 560898 161848 561134
rect 161528 560866 161848 560898
rect 171768 561454 172088 561486
rect 171768 561218 171810 561454
rect 172046 561218 172088 561454
rect 171768 561134 172088 561218
rect 171768 560898 171810 561134
rect 172046 560898 172088 561134
rect 171768 560866 172088 560898
rect 182008 561454 182328 561486
rect 182008 561218 182050 561454
rect 182286 561218 182328 561454
rect 182008 561134 182328 561218
rect 182008 560898 182050 561134
rect 182286 560898 182328 561134
rect 182008 560866 182328 560898
rect 192248 561454 192568 561486
rect 192248 561218 192290 561454
rect 192526 561218 192568 561454
rect 192248 561134 192568 561218
rect 192248 560898 192290 561134
rect 192526 560898 192568 561134
rect 192248 560866 192568 560898
rect 202488 561454 202808 561486
rect 202488 561218 202530 561454
rect 202766 561218 202808 561454
rect 202488 561134 202808 561218
rect 202488 560898 202530 561134
rect 202766 560898 202808 561134
rect 202488 560866 202808 560898
rect 212728 561454 213048 561486
rect 212728 561218 212770 561454
rect 213006 561218 213048 561454
rect 212728 561134 213048 561218
rect 212728 560898 212770 561134
rect 213006 560898 213048 561134
rect 212728 560866 213048 560898
rect 222968 561454 223288 561486
rect 222968 561218 223010 561454
rect 223246 561218 223288 561454
rect 222968 561134 223288 561218
rect 222968 560898 223010 561134
rect 223246 560898 223288 561134
rect 222968 560866 223288 560898
rect 233208 561454 233528 561486
rect 233208 561218 233250 561454
rect 233486 561218 233528 561454
rect 233208 561134 233528 561218
rect 233208 560898 233250 561134
rect 233486 560898 233528 561134
rect 233208 560866 233528 560898
rect 243448 561454 243768 561486
rect 243448 561218 243490 561454
rect 243726 561218 243768 561454
rect 243448 561134 243768 561218
rect 243448 560898 243490 561134
rect 243726 560898 243768 561134
rect 243448 560866 243768 560898
rect 253688 561454 254008 561486
rect 253688 561218 253730 561454
rect 253966 561218 254008 561454
rect 253688 561134 254008 561218
rect 253688 560898 253730 561134
rect 253966 560898 254008 561134
rect 253688 560866 254008 560898
rect 263928 561454 264248 561486
rect 263928 561218 263970 561454
rect 264206 561218 264248 561454
rect 263928 561134 264248 561218
rect 263928 560898 263970 561134
rect 264206 560898 264248 561134
rect 263928 560866 264248 560898
rect 274168 561454 274488 561486
rect 274168 561218 274210 561454
rect 274446 561218 274488 561454
rect 274168 561134 274488 561218
rect 274168 560898 274210 561134
rect 274446 560898 274488 561134
rect 274168 560866 274488 560898
rect 284408 561454 284728 561486
rect 284408 561218 284450 561454
rect 284686 561218 284728 561454
rect 284408 561134 284728 561218
rect 284408 560898 284450 561134
rect 284686 560898 284728 561134
rect 284408 560866 284728 560898
rect 294648 561454 294968 561486
rect 294648 561218 294690 561454
rect 294926 561218 294968 561454
rect 294648 561134 294968 561218
rect 294648 560898 294690 561134
rect 294926 560898 294968 561134
rect 294648 560866 294968 560898
rect 304888 561454 305208 561486
rect 304888 561218 304930 561454
rect 305166 561218 305208 561454
rect 304888 561134 305208 561218
rect 304888 560898 304930 561134
rect 305166 560898 305208 561134
rect 304888 560866 305208 560898
rect 315128 561454 315448 561486
rect 315128 561218 315170 561454
rect 315406 561218 315448 561454
rect 315128 561134 315448 561218
rect 315128 560898 315170 561134
rect 315406 560898 315448 561134
rect 315128 560866 315448 560898
rect 325368 561454 325688 561486
rect 325368 561218 325410 561454
rect 325646 561218 325688 561454
rect 325368 561134 325688 561218
rect 325368 560898 325410 561134
rect 325646 560898 325688 561134
rect 325368 560866 325688 560898
rect 335608 561454 335928 561486
rect 335608 561218 335650 561454
rect 335886 561218 335928 561454
rect 335608 561134 335928 561218
rect 335608 560898 335650 561134
rect 335886 560898 335928 561134
rect 335608 560866 335928 560898
rect 345848 561454 346168 561486
rect 345848 561218 345890 561454
rect 346126 561218 346168 561454
rect 345848 561134 346168 561218
rect 345848 560898 345890 561134
rect 346126 560898 346168 561134
rect 345848 560866 346168 560898
rect 356088 561454 356408 561486
rect 356088 561218 356130 561454
rect 356366 561218 356408 561454
rect 356088 561134 356408 561218
rect 356088 560898 356130 561134
rect 356366 560898 356408 561134
rect 356088 560866 356408 560898
rect 366328 561454 366648 561486
rect 366328 561218 366370 561454
rect 366606 561218 366648 561454
rect 366328 561134 366648 561218
rect 366328 560898 366370 561134
rect 366606 560898 366648 561134
rect 366328 560866 366648 560898
rect 376568 561454 376888 561486
rect 376568 561218 376610 561454
rect 376846 561218 376888 561454
rect 376568 561134 376888 561218
rect 376568 560898 376610 561134
rect 376846 560898 376888 561134
rect 376568 560866 376888 560898
rect 386808 561454 387128 561486
rect 386808 561218 386850 561454
rect 387086 561218 387128 561454
rect 386808 561134 387128 561218
rect 386808 560898 386850 561134
rect 387086 560898 387128 561134
rect 386808 560866 387128 560898
rect 397048 561454 397368 561486
rect 397048 561218 397090 561454
rect 397326 561218 397368 561454
rect 397048 561134 397368 561218
rect 397048 560898 397090 561134
rect 397326 560898 397368 561134
rect 397048 560866 397368 560898
rect 407288 561454 407608 561486
rect 407288 561218 407330 561454
rect 407566 561218 407608 561454
rect 407288 561134 407608 561218
rect 407288 560898 407330 561134
rect 407566 560898 407608 561134
rect 407288 560866 407608 560898
rect 417528 561454 417848 561486
rect 417528 561218 417570 561454
rect 417806 561218 417848 561454
rect 417528 561134 417848 561218
rect 417528 560898 417570 561134
rect 417806 560898 417848 561134
rect 417528 560866 417848 560898
rect 427768 561454 428088 561486
rect 427768 561218 427810 561454
rect 428046 561218 428088 561454
rect 427768 561134 428088 561218
rect 427768 560898 427810 561134
rect 428046 560898 428088 561134
rect 427768 560866 428088 560898
rect 438008 561454 438328 561486
rect 438008 561218 438050 561454
rect 438286 561218 438328 561454
rect 438008 561134 438328 561218
rect 438008 560898 438050 561134
rect 438286 560898 438328 561134
rect 438008 560866 438328 560898
rect 448248 561454 448568 561486
rect 448248 561218 448290 561454
rect 448526 561218 448568 561454
rect 448248 561134 448568 561218
rect 448248 560898 448290 561134
rect 448526 560898 448568 561134
rect 448248 560866 448568 560898
rect 458488 561454 458808 561486
rect 458488 561218 458530 561454
rect 458766 561218 458808 561454
rect 458488 561134 458808 561218
rect 458488 560898 458530 561134
rect 458766 560898 458808 561134
rect 458488 560866 458808 560898
rect 468728 561454 469048 561486
rect 468728 561218 468770 561454
rect 469006 561218 469048 561454
rect 468728 561134 469048 561218
rect 468728 560898 468770 561134
rect 469006 560898 469048 561134
rect 468728 560866 469048 560898
rect 478968 561454 479288 561486
rect 478968 561218 479010 561454
rect 479246 561218 479288 561454
rect 478968 561134 479288 561218
rect 478968 560898 479010 561134
rect 479246 560898 479288 561134
rect 478968 560866 479288 560898
rect 489208 561454 489528 561486
rect 489208 561218 489250 561454
rect 489486 561218 489528 561454
rect 489208 561134 489528 561218
rect 489208 560898 489250 561134
rect 489486 560898 489528 561134
rect 489208 560866 489528 560898
rect 499448 561454 499768 561486
rect 499448 561218 499490 561454
rect 499726 561218 499768 561454
rect 499448 561134 499768 561218
rect 499448 560898 499490 561134
rect 499726 560898 499768 561134
rect 499448 560866 499768 560898
rect 509688 561454 510008 561486
rect 509688 561218 509730 561454
rect 509966 561218 510008 561454
rect 509688 561134 510008 561218
rect 509688 560898 509730 561134
rect 509966 560898 510008 561134
rect 509688 560866 510008 560898
rect 519928 561454 520248 561486
rect 519928 561218 519970 561454
rect 520206 561218 520248 561454
rect 519928 561134 520248 561218
rect 519928 560898 519970 561134
rect 520206 560898 520248 561134
rect 519928 560866 520248 560898
rect 530168 561454 530488 561486
rect 530168 561218 530210 561454
rect 530446 561218 530488 561454
rect 530168 561134 530488 561218
rect 530168 560898 530210 561134
rect 530446 560898 530488 561134
rect 530168 560866 530488 560898
rect 15754 546938 15786 547174
rect 16022 546938 16106 547174
rect 16342 546938 16374 547174
rect 15754 546854 16374 546938
rect 15754 546618 15786 546854
rect 16022 546618 16106 546854
rect 16342 546618 16374 546854
rect 15754 511174 16374 546618
rect 541714 550894 542334 586338
rect 541714 550658 541746 550894
rect 541982 550658 542066 550894
rect 542302 550658 542334 550894
rect 541714 550574 542334 550658
rect 541714 550338 541746 550574
rect 541982 550338 542066 550574
rect 542302 550338 542334 550574
rect 23288 543454 23608 543486
rect 23288 543218 23330 543454
rect 23566 543218 23608 543454
rect 23288 543134 23608 543218
rect 23288 542898 23330 543134
rect 23566 542898 23608 543134
rect 23288 542866 23608 542898
rect 33528 543454 33848 543486
rect 33528 543218 33570 543454
rect 33806 543218 33848 543454
rect 33528 543134 33848 543218
rect 33528 542898 33570 543134
rect 33806 542898 33848 543134
rect 33528 542866 33848 542898
rect 43768 543454 44088 543486
rect 43768 543218 43810 543454
rect 44046 543218 44088 543454
rect 43768 543134 44088 543218
rect 43768 542898 43810 543134
rect 44046 542898 44088 543134
rect 43768 542866 44088 542898
rect 54008 543454 54328 543486
rect 54008 543218 54050 543454
rect 54286 543218 54328 543454
rect 54008 543134 54328 543218
rect 54008 542898 54050 543134
rect 54286 542898 54328 543134
rect 54008 542866 54328 542898
rect 64248 543454 64568 543486
rect 64248 543218 64290 543454
rect 64526 543218 64568 543454
rect 64248 543134 64568 543218
rect 64248 542898 64290 543134
rect 64526 542898 64568 543134
rect 64248 542866 64568 542898
rect 74488 543454 74808 543486
rect 74488 543218 74530 543454
rect 74766 543218 74808 543454
rect 74488 543134 74808 543218
rect 74488 542898 74530 543134
rect 74766 542898 74808 543134
rect 74488 542866 74808 542898
rect 84728 543454 85048 543486
rect 84728 543218 84770 543454
rect 85006 543218 85048 543454
rect 84728 543134 85048 543218
rect 84728 542898 84770 543134
rect 85006 542898 85048 543134
rect 84728 542866 85048 542898
rect 94968 543454 95288 543486
rect 94968 543218 95010 543454
rect 95246 543218 95288 543454
rect 94968 543134 95288 543218
rect 94968 542898 95010 543134
rect 95246 542898 95288 543134
rect 94968 542866 95288 542898
rect 105208 543454 105528 543486
rect 105208 543218 105250 543454
rect 105486 543218 105528 543454
rect 105208 543134 105528 543218
rect 105208 542898 105250 543134
rect 105486 542898 105528 543134
rect 105208 542866 105528 542898
rect 115448 543454 115768 543486
rect 115448 543218 115490 543454
rect 115726 543218 115768 543454
rect 115448 543134 115768 543218
rect 115448 542898 115490 543134
rect 115726 542898 115768 543134
rect 115448 542866 115768 542898
rect 125688 543454 126008 543486
rect 125688 543218 125730 543454
rect 125966 543218 126008 543454
rect 125688 543134 126008 543218
rect 125688 542898 125730 543134
rect 125966 542898 126008 543134
rect 125688 542866 126008 542898
rect 135928 543454 136248 543486
rect 135928 543218 135970 543454
rect 136206 543218 136248 543454
rect 135928 543134 136248 543218
rect 135928 542898 135970 543134
rect 136206 542898 136248 543134
rect 135928 542866 136248 542898
rect 146168 543454 146488 543486
rect 146168 543218 146210 543454
rect 146446 543218 146488 543454
rect 146168 543134 146488 543218
rect 146168 542898 146210 543134
rect 146446 542898 146488 543134
rect 146168 542866 146488 542898
rect 156408 543454 156728 543486
rect 156408 543218 156450 543454
rect 156686 543218 156728 543454
rect 156408 543134 156728 543218
rect 156408 542898 156450 543134
rect 156686 542898 156728 543134
rect 156408 542866 156728 542898
rect 166648 543454 166968 543486
rect 166648 543218 166690 543454
rect 166926 543218 166968 543454
rect 166648 543134 166968 543218
rect 166648 542898 166690 543134
rect 166926 542898 166968 543134
rect 166648 542866 166968 542898
rect 176888 543454 177208 543486
rect 176888 543218 176930 543454
rect 177166 543218 177208 543454
rect 176888 543134 177208 543218
rect 176888 542898 176930 543134
rect 177166 542898 177208 543134
rect 176888 542866 177208 542898
rect 187128 543454 187448 543486
rect 187128 543218 187170 543454
rect 187406 543218 187448 543454
rect 187128 543134 187448 543218
rect 187128 542898 187170 543134
rect 187406 542898 187448 543134
rect 187128 542866 187448 542898
rect 197368 543454 197688 543486
rect 197368 543218 197410 543454
rect 197646 543218 197688 543454
rect 197368 543134 197688 543218
rect 197368 542898 197410 543134
rect 197646 542898 197688 543134
rect 197368 542866 197688 542898
rect 207608 543454 207928 543486
rect 207608 543218 207650 543454
rect 207886 543218 207928 543454
rect 207608 543134 207928 543218
rect 207608 542898 207650 543134
rect 207886 542898 207928 543134
rect 207608 542866 207928 542898
rect 217848 543454 218168 543486
rect 217848 543218 217890 543454
rect 218126 543218 218168 543454
rect 217848 543134 218168 543218
rect 217848 542898 217890 543134
rect 218126 542898 218168 543134
rect 217848 542866 218168 542898
rect 228088 543454 228408 543486
rect 228088 543218 228130 543454
rect 228366 543218 228408 543454
rect 228088 543134 228408 543218
rect 228088 542898 228130 543134
rect 228366 542898 228408 543134
rect 228088 542866 228408 542898
rect 238328 543454 238648 543486
rect 238328 543218 238370 543454
rect 238606 543218 238648 543454
rect 238328 543134 238648 543218
rect 238328 542898 238370 543134
rect 238606 542898 238648 543134
rect 238328 542866 238648 542898
rect 248568 543454 248888 543486
rect 248568 543218 248610 543454
rect 248846 543218 248888 543454
rect 248568 543134 248888 543218
rect 248568 542898 248610 543134
rect 248846 542898 248888 543134
rect 248568 542866 248888 542898
rect 258808 543454 259128 543486
rect 258808 543218 258850 543454
rect 259086 543218 259128 543454
rect 258808 543134 259128 543218
rect 258808 542898 258850 543134
rect 259086 542898 259128 543134
rect 258808 542866 259128 542898
rect 269048 543454 269368 543486
rect 269048 543218 269090 543454
rect 269326 543218 269368 543454
rect 269048 543134 269368 543218
rect 269048 542898 269090 543134
rect 269326 542898 269368 543134
rect 269048 542866 269368 542898
rect 279288 543454 279608 543486
rect 279288 543218 279330 543454
rect 279566 543218 279608 543454
rect 279288 543134 279608 543218
rect 279288 542898 279330 543134
rect 279566 542898 279608 543134
rect 279288 542866 279608 542898
rect 289528 543454 289848 543486
rect 289528 543218 289570 543454
rect 289806 543218 289848 543454
rect 289528 543134 289848 543218
rect 289528 542898 289570 543134
rect 289806 542898 289848 543134
rect 289528 542866 289848 542898
rect 299768 543454 300088 543486
rect 299768 543218 299810 543454
rect 300046 543218 300088 543454
rect 299768 543134 300088 543218
rect 299768 542898 299810 543134
rect 300046 542898 300088 543134
rect 299768 542866 300088 542898
rect 310008 543454 310328 543486
rect 310008 543218 310050 543454
rect 310286 543218 310328 543454
rect 310008 543134 310328 543218
rect 310008 542898 310050 543134
rect 310286 542898 310328 543134
rect 310008 542866 310328 542898
rect 320248 543454 320568 543486
rect 320248 543218 320290 543454
rect 320526 543218 320568 543454
rect 320248 543134 320568 543218
rect 320248 542898 320290 543134
rect 320526 542898 320568 543134
rect 320248 542866 320568 542898
rect 330488 543454 330808 543486
rect 330488 543218 330530 543454
rect 330766 543218 330808 543454
rect 330488 543134 330808 543218
rect 330488 542898 330530 543134
rect 330766 542898 330808 543134
rect 330488 542866 330808 542898
rect 340728 543454 341048 543486
rect 340728 543218 340770 543454
rect 341006 543218 341048 543454
rect 340728 543134 341048 543218
rect 340728 542898 340770 543134
rect 341006 542898 341048 543134
rect 340728 542866 341048 542898
rect 350968 543454 351288 543486
rect 350968 543218 351010 543454
rect 351246 543218 351288 543454
rect 350968 543134 351288 543218
rect 350968 542898 351010 543134
rect 351246 542898 351288 543134
rect 350968 542866 351288 542898
rect 361208 543454 361528 543486
rect 361208 543218 361250 543454
rect 361486 543218 361528 543454
rect 361208 543134 361528 543218
rect 361208 542898 361250 543134
rect 361486 542898 361528 543134
rect 361208 542866 361528 542898
rect 371448 543454 371768 543486
rect 371448 543218 371490 543454
rect 371726 543218 371768 543454
rect 371448 543134 371768 543218
rect 371448 542898 371490 543134
rect 371726 542898 371768 543134
rect 371448 542866 371768 542898
rect 381688 543454 382008 543486
rect 381688 543218 381730 543454
rect 381966 543218 382008 543454
rect 381688 543134 382008 543218
rect 381688 542898 381730 543134
rect 381966 542898 382008 543134
rect 381688 542866 382008 542898
rect 391928 543454 392248 543486
rect 391928 543218 391970 543454
rect 392206 543218 392248 543454
rect 391928 543134 392248 543218
rect 391928 542898 391970 543134
rect 392206 542898 392248 543134
rect 391928 542866 392248 542898
rect 402168 543454 402488 543486
rect 402168 543218 402210 543454
rect 402446 543218 402488 543454
rect 402168 543134 402488 543218
rect 402168 542898 402210 543134
rect 402446 542898 402488 543134
rect 402168 542866 402488 542898
rect 412408 543454 412728 543486
rect 412408 543218 412450 543454
rect 412686 543218 412728 543454
rect 412408 543134 412728 543218
rect 412408 542898 412450 543134
rect 412686 542898 412728 543134
rect 412408 542866 412728 542898
rect 422648 543454 422968 543486
rect 422648 543218 422690 543454
rect 422926 543218 422968 543454
rect 422648 543134 422968 543218
rect 422648 542898 422690 543134
rect 422926 542898 422968 543134
rect 422648 542866 422968 542898
rect 432888 543454 433208 543486
rect 432888 543218 432930 543454
rect 433166 543218 433208 543454
rect 432888 543134 433208 543218
rect 432888 542898 432930 543134
rect 433166 542898 433208 543134
rect 432888 542866 433208 542898
rect 443128 543454 443448 543486
rect 443128 543218 443170 543454
rect 443406 543218 443448 543454
rect 443128 543134 443448 543218
rect 443128 542898 443170 543134
rect 443406 542898 443448 543134
rect 443128 542866 443448 542898
rect 453368 543454 453688 543486
rect 453368 543218 453410 543454
rect 453646 543218 453688 543454
rect 453368 543134 453688 543218
rect 453368 542898 453410 543134
rect 453646 542898 453688 543134
rect 453368 542866 453688 542898
rect 463608 543454 463928 543486
rect 463608 543218 463650 543454
rect 463886 543218 463928 543454
rect 463608 543134 463928 543218
rect 463608 542898 463650 543134
rect 463886 542898 463928 543134
rect 463608 542866 463928 542898
rect 473848 543454 474168 543486
rect 473848 543218 473890 543454
rect 474126 543218 474168 543454
rect 473848 543134 474168 543218
rect 473848 542898 473890 543134
rect 474126 542898 474168 543134
rect 473848 542866 474168 542898
rect 484088 543454 484408 543486
rect 484088 543218 484130 543454
rect 484366 543218 484408 543454
rect 484088 543134 484408 543218
rect 484088 542898 484130 543134
rect 484366 542898 484408 543134
rect 484088 542866 484408 542898
rect 494328 543454 494648 543486
rect 494328 543218 494370 543454
rect 494606 543218 494648 543454
rect 494328 543134 494648 543218
rect 494328 542898 494370 543134
rect 494606 542898 494648 543134
rect 494328 542866 494648 542898
rect 504568 543454 504888 543486
rect 504568 543218 504610 543454
rect 504846 543218 504888 543454
rect 504568 543134 504888 543218
rect 504568 542898 504610 543134
rect 504846 542898 504888 543134
rect 504568 542866 504888 542898
rect 514808 543454 515128 543486
rect 514808 543218 514850 543454
rect 515086 543218 515128 543454
rect 514808 543134 515128 543218
rect 514808 542898 514850 543134
rect 515086 542898 515128 543134
rect 514808 542866 515128 542898
rect 525048 543454 525368 543486
rect 525048 543218 525090 543454
rect 525326 543218 525368 543454
rect 525048 543134 525368 543218
rect 525048 542898 525090 543134
rect 525326 542898 525368 543134
rect 525048 542866 525368 542898
rect 535288 543454 535608 543486
rect 535288 543218 535330 543454
rect 535566 543218 535608 543454
rect 535288 543134 535608 543218
rect 535288 542898 535330 543134
rect 535566 542898 535608 543134
rect 535288 542866 535608 542898
rect 28408 525454 28728 525486
rect 28408 525218 28450 525454
rect 28686 525218 28728 525454
rect 28408 525134 28728 525218
rect 28408 524898 28450 525134
rect 28686 524898 28728 525134
rect 28408 524866 28728 524898
rect 38648 525454 38968 525486
rect 38648 525218 38690 525454
rect 38926 525218 38968 525454
rect 38648 525134 38968 525218
rect 38648 524898 38690 525134
rect 38926 524898 38968 525134
rect 38648 524866 38968 524898
rect 48888 525454 49208 525486
rect 48888 525218 48930 525454
rect 49166 525218 49208 525454
rect 48888 525134 49208 525218
rect 48888 524898 48930 525134
rect 49166 524898 49208 525134
rect 48888 524866 49208 524898
rect 59128 525454 59448 525486
rect 59128 525218 59170 525454
rect 59406 525218 59448 525454
rect 59128 525134 59448 525218
rect 59128 524898 59170 525134
rect 59406 524898 59448 525134
rect 59128 524866 59448 524898
rect 69368 525454 69688 525486
rect 69368 525218 69410 525454
rect 69646 525218 69688 525454
rect 69368 525134 69688 525218
rect 69368 524898 69410 525134
rect 69646 524898 69688 525134
rect 69368 524866 69688 524898
rect 79608 525454 79928 525486
rect 79608 525218 79650 525454
rect 79886 525218 79928 525454
rect 79608 525134 79928 525218
rect 79608 524898 79650 525134
rect 79886 524898 79928 525134
rect 79608 524866 79928 524898
rect 89848 525454 90168 525486
rect 89848 525218 89890 525454
rect 90126 525218 90168 525454
rect 89848 525134 90168 525218
rect 89848 524898 89890 525134
rect 90126 524898 90168 525134
rect 89848 524866 90168 524898
rect 100088 525454 100408 525486
rect 100088 525218 100130 525454
rect 100366 525218 100408 525454
rect 100088 525134 100408 525218
rect 100088 524898 100130 525134
rect 100366 524898 100408 525134
rect 100088 524866 100408 524898
rect 110328 525454 110648 525486
rect 110328 525218 110370 525454
rect 110606 525218 110648 525454
rect 110328 525134 110648 525218
rect 110328 524898 110370 525134
rect 110606 524898 110648 525134
rect 110328 524866 110648 524898
rect 120568 525454 120888 525486
rect 120568 525218 120610 525454
rect 120846 525218 120888 525454
rect 120568 525134 120888 525218
rect 120568 524898 120610 525134
rect 120846 524898 120888 525134
rect 120568 524866 120888 524898
rect 130808 525454 131128 525486
rect 130808 525218 130850 525454
rect 131086 525218 131128 525454
rect 130808 525134 131128 525218
rect 130808 524898 130850 525134
rect 131086 524898 131128 525134
rect 130808 524866 131128 524898
rect 141048 525454 141368 525486
rect 141048 525218 141090 525454
rect 141326 525218 141368 525454
rect 141048 525134 141368 525218
rect 141048 524898 141090 525134
rect 141326 524898 141368 525134
rect 141048 524866 141368 524898
rect 151288 525454 151608 525486
rect 151288 525218 151330 525454
rect 151566 525218 151608 525454
rect 151288 525134 151608 525218
rect 151288 524898 151330 525134
rect 151566 524898 151608 525134
rect 151288 524866 151608 524898
rect 161528 525454 161848 525486
rect 161528 525218 161570 525454
rect 161806 525218 161848 525454
rect 161528 525134 161848 525218
rect 161528 524898 161570 525134
rect 161806 524898 161848 525134
rect 161528 524866 161848 524898
rect 171768 525454 172088 525486
rect 171768 525218 171810 525454
rect 172046 525218 172088 525454
rect 171768 525134 172088 525218
rect 171768 524898 171810 525134
rect 172046 524898 172088 525134
rect 171768 524866 172088 524898
rect 182008 525454 182328 525486
rect 182008 525218 182050 525454
rect 182286 525218 182328 525454
rect 182008 525134 182328 525218
rect 182008 524898 182050 525134
rect 182286 524898 182328 525134
rect 182008 524866 182328 524898
rect 192248 525454 192568 525486
rect 192248 525218 192290 525454
rect 192526 525218 192568 525454
rect 192248 525134 192568 525218
rect 192248 524898 192290 525134
rect 192526 524898 192568 525134
rect 192248 524866 192568 524898
rect 202488 525454 202808 525486
rect 202488 525218 202530 525454
rect 202766 525218 202808 525454
rect 202488 525134 202808 525218
rect 202488 524898 202530 525134
rect 202766 524898 202808 525134
rect 202488 524866 202808 524898
rect 212728 525454 213048 525486
rect 212728 525218 212770 525454
rect 213006 525218 213048 525454
rect 212728 525134 213048 525218
rect 212728 524898 212770 525134
rect 213006 524898 213048 525134
rect 212728 524866 213048 524898
rect 222968 525454 223288 525486
rect 222968 525218 223010 525454
rect 223246 525218 223288 525454
rect 222968 525134 223288 525218
rect 222968 524898 223010 525134
rect 223246 524898 223288 525134
rect 222968 524866 223288 524898
rect 233208 525454 233528 525486
rect 233208 525218 233250 525454
rect 233486 525218 233528 525454
rect 233208 525134 233528 525218
rect 233208 524898 233250 525134
rect 233486 524898 233528 525134
rect 233208 524866 233528 524898
rect 243448 525454 243768 525486
rect 243448 525218 243490 525454
rect 243726 525218 243768 525454
rect 243448 525134 243768 525218
rect 243448 524898 243490 525134
rect 243726 524898 243768 525134
rect 243448 524866 243768 524898
rect 253688 525454 254008 525486
rect 253688 525218 253730 525454
rect 253966 525218 254008 525454
rect 253688 525134 254008 525218
rect 253688 524898 253730 525134
rect 253966 524898 254008 525134
rect 253688 524866 254008 524898
rect 263928 525454 264248 525486
rect 263928 525218 263970 525454
rect 264206 525218 264248 525454
rect 263928 525134 264248 525218
rect 263928 524898 263970 525134
rect 264206 524898 264248 525134
rect 263928 524866 264248 524898
rect 274168 525454 274488 525486
rect 274168 525218 274210 525454
rect 274446 525218 274488 525454
rect 274168 525134 274488 525218
rect 274168 524898 274210 525134
rect 274446 524898 274488 525134
rect 274168 524866 274488 524898
rect 284408 525454 284728 525486
rect 284408 525218 284450 525454
rect 284686 525218 284728 525454
rect 284408 525134 284728 525218
rect 284408 524898 284450 525134
rect 284686 524898 284728 525134
rect 284408 524866 284728 524898
rect 294648 525454 294968 525486
rect 294648 525218 294690 525454
rect 294926 525218 294968 525454
rect 294648 525134 294968 525218
rect 294648 524898 294690 525134
rect 294926 524898 294968 525134
rect 294648 524866 294968 524898
rect 304888 525454 305208 525486
rect 304888 525218 304930 525454
rect 305166 525218 305208 525454
rect 304888 525134 305208 525218
rect 304888 524898 304930 525134
rect 305166 524898 305208 525134
rect 304888 524866 305208 524898
rect 315128 525454 315448 525486
rect 315128 525218 315170 525454
rect 315406 525218 315448 525454
rect 315128 525134 315448 525218
rect 315128 524898 315170 525134
rect 315406 524898 315448 525134
rect 315128 524866 315448 524898
rect 325368 525454 325688 525486
rect 325368 525218 325410 525454
rect 325646 525218 325688 525454
rect 325368 525134 325688 525218
rect 325368 524898 325410 525134
rect 325646 524898 325688 525134
rect 325368 524866 325688 524898
rect 335608 525454 335928 525486
rect 335608 525218 335650 525454
rect 335886 525218 335928 525454
rect 335608 525134 335928 525218
rect 335608 524898 335650 525134
rect 335886 524898 335928 525134
rect 335608 524866 335928 524898
rect 345848 525454 346168 525486
rect 345848 525218 345890 525454
rect 346126 525218 346168 525454
rect 345848 525134 346168 525218
rect 345848 524898 345890 525134
rect 346126 524898 346168 525134
rect 345848 524866 346168 524898
rect 356088 525454 356408 525486
rect 356088 525218 356130 525454
rect 356366 525218 356408 525454
rect 356088 525134 356408 525218
rect 356088 524898 356130 525134
rect 356366 524898 356408 525134
rect 356088 524866 356408 524898
rect 366328 525454 366648 525486
rect 366328 525218 366370 525454
rect 366606 525218 366648 525454
rect 366328 525134 366648 525218
rect 366328 524898 366370 525134
rect 366606 524898 366648 525134
rect 366328 524866 366648 524898
rect 376568 525454 376888 525486
rect 376568 525218 376610 525454
rect 376846 525218 376888 525454
rect 376568 525134 376888 525218
rect 376568 524898 376610 525134
rect 376846 524898 376888 525134
rect 376568 524866 376888 524898
rect 386808 525454 387128 525486
rect 386808 525218 386850 525454
rect 387086 525218 387128 525454
rect 386808 525134 387128 525218
rect 386808 524898 386850 525134
rect 387086 524898 387128 525134
rect 386808 524866 387128 524898
rect 397048 525454 397368 525486
rect 397048 525218 397090 525454
rect 397326 525218 397368 525454
rect 397048 525134 397368 525218
rect 397048 524898 397090 525134
rect 397326 524898 397368 525134
rect 397048 524866 397368 524898
rect 407288 525454 407608 525486
rect 407288 525218 407330 525454
rect 407566 525218 407608 525454
rect 407288 525134 407608 525218
rect 407288 524898 407330 525134
rect 407566 524898 407608 525134
rect 407288 524866 407608 524898
rect 417528 525454 417848 525486
rect 417528 525218 417570 525454
rect 417806 525218 417848 525454
rect 417528 525134 417848 525218
rect 417528 524898 417570 525134
rect 417806 524898 417848 525134
rect 417528 524866 417848 524898
rect 427768 525454 428088 525486
rect 427768 525218 427810 525454
rect 428046 525218 428088 525454
rect 427768 525134 428088 525218
rect 427768 524898 427810 525134
rect 428046 524898 428088 525134
rect 427768 524866 428088 524898
rect 438008 525454 438328 525486
rect 438008 525218 438050 525454
rect 438286 525218 438328 525454
rect 438008 525134 438328 525218
rect 438008 524898 438050 525134
rect 438286 524898 438328 525134
rect 438008 524866 438328 524898
rect 448248 525454 448568 525486
rect 448248 525218 448290 525454
rect 448526 525218 448568 525454
rect 448248 525134 448568 525218
rect 448248 524898 448290 525134
rect 448526 524898 448568 525134
rect 448248 524866 448568 524898
rect 458488 525454 458808 525486
rect 458488 525218 458530 525454
rect 458766 525218 458808 525454
rect 458488 525134 458808 525218
rect 458488 524898 458530 525134
rect 458766 524898 458808 525134
rect 458488 524866 458808 524898
rect 468728 525454 469048 525486
rect 468728 525218 468770 525454
rect 469006 525218 469048 525454
rect 468728 525134 469048 525218
rect 468728 524898 468770 525134
rect 469006 524898 469048 525134
rect 468728 524866 469048 524898
rect 478968 525454 479288 525486
rect 478968 525218 479010 525454
rect 479246 525218 479288 525454
rect 478968 525134 479288 525218
rect 478968 524898 479010 525134
rect 479246 524898 479288 525134
rect 478968 524866 479288 524898
rect 489208 525454 489528 525486
rect 489208 525218 489250 525454
rect 489486 525218 489528 525454
rect 489208 525134 489528 525218
rect 489208 524898 489250 525134
rect 489486 524898 489528 525134
rect 489208 524866 489528 524898
rect 499448 525454 499768 525486
rect 499448 525218 499490 525454
rect 499726 525218 499768 525454
rect 499448 525134 499768 525218
rect 499448 524898 499490 525134
rect 499726 524898 499768 525134
rect 499448 524866 499768 524898
rect 509688 525454 510008 525486
rect 509688 525218 509730 525454
rect 509966 525218 510008 525454
rect 509688 525134 510008 525218
rect 509688 524898 509730 525134
rect 509966 524898 510008 525134
rect 509688 524866 510008 524898
rect 519928 525454 520248 525486
rect 519928 525218 519970 525454
rect 520206 525218 520248 525454
rect 519928 525134 520248 525218
rect 519928 524898 519970 525134
rect 520206 524898 520248 525134
rect 519928 524866 520248 524898
rect 530168 525454 530488 525486
rect 530168 525218 530210 525454
rect 530446 525218 530488 525454
rect 530168 525134 530488 525218
rect 530168 524898 530210 525134
rect 530446 524898 530488 525134
rect 530168 524866 530488 524898
rect 15754 510938 15786 511174
rect 16022 510938 16106 511174
rect 16342 510938 16374 511174
rect 15754 510854 16374 510938
rect 15754 510618 15786 510854
rect 16022 510618 16106 510854
rect 16342 510618 16374 510854
rect 15754 475174 16374 510618
rect 541714 514894 542334 550338
rect 541714 514658 541746 514894
rect 541982 514658 542066 514894
rect 542302 514658 542334 514894
rect 541714 514574 542334 514658
rect 541714 514338 541746 514574
rect 541982 514338 542066 514574
rect 542302 514338 542334 514574
rect 23288 507454 23608 507486
rect 23288 507218 23330 507454
rect 23566 507218 23608 507454
rect 23288 507134 23608 507218
rect 23288 506898 23330 507134
rect 23566 506898 23608 507134
rect 23288 506866 23608 506898
rect 33528 507454 33848 507486
rect 33528 507218 33570 507454
rect 33806 507218 33848 507454
rect 33528 507134 33848 507218
rect 33528 506898 33570 507134
rect 33806 506898 33848 507134
rect 33528 506866 33848 506898
rect 43768 507454 44088 507486
rect 43768 507218 43810 507454
rect 44046 507218 44088 507454
rect 43768 507134 44088 507218
rect 43768 506898 43810 507134
rect 44046 506898 44088 507134
rect 43768 506866 44088 506898
rect 54008 507454 54328 507486
rect 54008 507218 54050 507454
rect 54286 507218 54328 507454
rect 54008 507134 54328 507218
rect 54008 506898 54050 507134
rect 54286 506898 54328 507134
rect 54008 506866 54328 506898
rect 64248 507454 64568 507486
rect 64248 507218 64290 507454
rect 64526 507218 64568 507454
rect 64248 507134 64568 507218
rect 64248 506898 64290 507134
rect 64526 506898 64568 507134
rect 64248 506866 64568 506898
rect 74488 507454 74808 507486
rect 74488 507218 74530 507454
rect 74766 507218 74808 507454
rect 74488 507134 74808 507218
rect 74488 506898 74530 507134
rect 74766 506898 74808 507134
rect 74488 506866 74808 506898
rect 84728 507454 85048 507486
rect 84728 507218 84770 507454
rect 85006 507218 85048 507454
rect 84728 507134 85048 507218
rect 84728 506898 84770 507134
rect 85006 506898 85048 507134
rect 84728 506866 85048 506898
rect 94968 507454 95288 507486
rect 94968 507218 95010 507454
rect 95246 507218 95288 507454
rect 94968 507134 95288 507218
rect 94968 506898 95010 507134
rect 95246 506898 95288 507134
rect 94968 506866 95288 506898
rect 105208 507454 105528 507486
rect 105208 507218 105250 507454
rect 105486 507218 105528 507454
rect 105208 507134 105528 507218
rect 105208 506898 105250 507134
rect 105486 506898 105528 507134
rect 105208 506866 105528 506898
rect 115448 507454 115768 507486
rect 115448 507218 115490 507454
rect 115726 507218 115768 507454
rect 115448 507134 115768 507218
rect 115448 506898 115490 507134
rect 115726 506898 115768 507134
rect 115448 506866 115768 506898
rect 125688 507454 126008 507486
rect 125688 507218 125730 507454
rect 125966 507218 126008 507454
rect 125688 507134 126008 507218
rect 125688 506898 125730 507134
rect 125966 506898 126008 507134
rect 125688 506866 126008 506898
rect 135928 507454 136248 507486
rect 135928 507218 135970 507454
rect 136206 507218 136248 507454
rect 135928 507134 136248 507218
rect 135928 506898 135970 507134
rect 136206 506898 136248 507134
rect 135928 506866 136248 506898
rect 146168 507454 146488 507486
rect 146168 507218 146210 507454
rect 146446 507218 146488 507454
rect 146168 507134 146488 507218
rect 146168 506898 146210 507134
rect 146446 506898 146488 507134
rect 146168 506866 146488 506898
rect 156408 507454 156728 507486
rect 156408 507218 156450 507454
rect 156686 507218 156728 507454
rect 156408 507134 156728 507218
rect 156408 506898 156450 507134
rect 156686 506898 156728 507134
rect 156408 506866 156728 506898
rect 166648 507454 166968 507486
rect 166648 507218 166690 507454
rect 166926 507218 166968 507454
rect 166648 507134 166968 507218
rect 166648 506898 166690 507134
rect 166926 506898 166968 507134
rect 166648 506866 166968 506898
rect 176888 507454 177208 507486
rect 176888 507218 176930 507454
rect 177166 507218 177208 507454
rect 176888 507134 177208 507218
rect 176888 506898 176930 507134
rect 177166 506898 177208 507134
rect 176888 506866 177208 506898
rect 187128 507454 187448 507486
rect 187128 507218 187170 507454
rect 187406 507218 187448 507454
rect 187128 507134 187448 507218
rect 187128 506898 187170 507134
rect 187406 506898 187448 507134
rect 187128 506866 187448 506898
rect 197368 507454 197688 507486
rect 197368 507218 197410 507454
rect 197646 507218 197688 507454
rect 197368 507134 197688 507218
rect 197368 506898 197410 507134
rect 197646 506898 197688 507134
rect 197368 506866 197688 506898
rect 207608 507454 207928 507486
rect 207608 507218 207650 507454
rect 207886 507218 207928 507454
rect 207608 507134 207928 507218
rect 207608 506898 207650 507134
rect 207886 506898 207928 507134
rect 207608 506866 207928 506898
rect 217848 507454 218168 507486
rect 217848 507218 217890 507454
rect 218126 507218 218168 507454
rect 217848 507134 218168 507218
rect 217848 506898 217890 507134
rect 218126 506898 218168 507134
rect 217848 506866 218168 506898
rect 228088 507454 228408 507486
rect 228088 507218 228130 507454
rect 228366 507218 228408 507454
rect 228088 507134 228408 507218
rect 228088 506898 228130 507134
rect 228366 506898 228408 507134
rect 228088 506866 228408 506898
rect 238328 507454 238648 507486
rect 238328 507218 238370 507454
rect 238606 507218 238648 507454
rect 238328 507134 238648 507218
rect 238328 506898 238370 507134
rect 238606 506898 238648 507134
rect 238328 506866 238648 506898
rect 248568 507454 248888 507486
rect 248568 507218 248610 507454
rect 248846 507218 248888 507454
rect 248568 507134 248888 507218
rect 248568 506898 248610 507134
rect 248846 506898 248888 507134
rect 248568 506866 248888 506898
rect 258808 507454 259128 507486
rect 258808 507218 258850 507454
rect 259086 507218 259128 507454
rect 258808 507134 259128 507218
rect 258808 506898 258850 507134
rect 259086 506898 259128 507134
rect 258808 506866 259128 506898
rect 269048 507454 269368 507486
rect 269048 507218 269090 507454
rect 269326 507218 269368 507454
rect 269048 507134 269368 507218
rect 269048 506898 269090 507134
rect 269326 506898 269368 507134
rect 269048 506866 269368 506898
rect 279288 507454 279608 507486
rect 279288 507218 279330 507454
rect 279566 507218 279608 507454
rect 279288 507134 279608 507218
rect 279288 506898 279330 507134
rect 279566 506898 279608 507134
rect 279288 506866 279608 506898
rect 289528 507454 289848 507486
rect 289528 507218 289570 507454
rect 289806 507218 289848 507454
rect 289528 507134 289848 507218
rect 289528 506898 289570 507134
rect 289806 506898 289848 507134
rect 289528 506866 289848 506898
rect 299768 507454 300088 507486
rect 299768 507218 299810 507454
rect 300046 507218 300088 507454
rect 299768 507134 300088 507218
rect 299768 506898 299810 507134
rect 300046 506898 300088 507134
rect 299768 506866 300088 506898
rect 310008 507454 310328 507486
rect 310008 507218 310050 507454
rect 310286 507218 310328 507454
rect 310008 507134 310328 507218
rect 310008 506898 310050 507134
rect 310286 506898 310328 507134
rect 310008 506866 310328 506898
rect 320248 507454 320568 507486
rect 320248 507218 320290 507454
rect 320526 507218 320568 507454
rect 320248 507134 320568 507218
rect 320248 506898 320290 507134
rect 320526 506898 320568 507134
rect 320248 506866 320568 506898
rect 330488 507454 330808 507486
rect 330488 507218 330530 507454
rect 330766 507218 330808 507454
rect 330488 507134 330808 507218
rect 330488 506898 330530 507134
rect 330766 506898 330808 507134
rect 330488 506866 330808 506898
rect 340728 507454 341048 507486
rect 340728 507218 340770 507454
rect 341006 507218 341048 507454
rect 340728 507134 341048 507218
rect 340728 506898 340770 507134
rect 341006 506898 341048 507134
rect 340728 506866 341048 506898
rect 350968 507454 351288 507486
rect 350968 507218 351010 507454
rect 351246 507218 351288 507454
rect 350968 507134 351288 507218
rect 350968 506898 351010 507134
rect 351246 506898 351288 507134
rect 350968 506866 351288 506898
rect 361208 507454 361528 507486
rect 361208 507218 361250 507454
rect 361486 507218 361528 507454
rect 361208 507134 361528 507218
rect 361208 506898 361250 507134
rect 361486 506898 361528 507134
rect 361208 506866 361528 506898
rect 371448 507454 371768 507486
rect 371448 507218 371490 507454
rect 371726 507218 371768 507454
rect 371448 507134 371768 507218
rect 371448 506898 371490 507134
rect 371726 506898 371768 507134
rect 371448 506866 371768 506898
rect 381688 507454 382008 507486
rect 381688 507218 381730 507454
rect 381966 507218 382008 507454
rect 381688 507134 382008 507218
rect 381688 506898 381730 507134
rect 381966 506898 382008 507134
rect 381688 506866 382008 506898
rect 391928 507454 392248 507486
rect 391928 507218 391970 507454
rect 392206 507218 392248 507454
rect 391928 507134 392248 507218
rect 391928 506898 391970 507134
rect 392206 506898 392248 507134
rect 391928 506866 392248 506898
rect 402168 507454 402488 507486
rect 402168 507218 402210 507454
rect 402446 507218 402488 507454
rect 402168 507134 402488 507218
rect 402168 506898 402210 507134
rect 402446 506898 402488 507134
rect 402168 506866 402488 506898
rect 412408 507454 412728 507486
rect 412408 507218 412450 507454
rect 412686 507218 412728 507454
rect 412408 507134 412728 507218
rect 412408 506898 412450 507134
rect 412686 506898 412728 507134
rect 412408 506866 412728 506898
rect 422648 507454 422968 507486
rect 422648 507218 422690 507454
rect 422926 507218 422968 507454
rect 422648 507134 422968 507218
rect 422648 506898 422690 507134
rect 422926 506898 422968 507134
rect 422648 506866 422968 506898
rect 432888 507454 433208 507486
rect 432888 507218 432930 507454
rect 433166 507218 433208 507454
rect 432888 507134 433208 507218
rect 432888 506898 432930 507134
rect 433166 506898 433208 507134
rect 432888 506866 433208 506898
rect 443128 507454 443448 507486
rect 443128 507218 443170 507454
rect 443406 507218 443448 507454
rect 443128 507134 443448 507218
rect 443128 506898 443170 507134
rect 443406 506898 443448 507134
rect 443128 506866 443448 506898
rect 453368 507454 453688 507486
rect 453368 507218 453410 507454
rect 453646 507218 453688 507454
rect 453368 507134 453688 507218
rect 453368 506898 453410 507134
rect 453646 506898 453688 507134
rect 453368 506866 453688 506898
rect 463608 507454 463928 507486
rect 463608 507218 463650 507454
rect 463886 507218 463928 507454
rect 463608 507134 463928 507218
rect 463608 506898 463650 507134
rect 463886 506898 463928 507134
rect 463608 506866 463928 506898
rect 473848 507454 474168 507486
rect 473848 507218 473890 507454
rect 474126 507218 474168 507454
rect 473848 507134 474168 507218
rect 473848 506898 473890 507134
rect 474126 506898 474168 507134
rect 473848 506866 474168 506898
rect 484088 507454 484408 507486
rect 484088 507218 484130 507454
rect 484366 507218 484408 507454
rect 484088 507134 484408 507218
rect 484088 506898 484130 507134
rect 484366 506898 484408 507134
rect 484088 506866 484408 506898
rect 494328 507454 494648 507486
rect 494328 507218 494370 507454
rect 494606 507218 494648 507454
rect 494328 507134 494648 507218
rect 494328 506898 494370 507134
rect 494606 506898 494648 507134
rect 494328 506866 494648 506898
rect 504568 507454 504888 507486
rect 504568 507218 504610 507454
rect 504846 507218 504888 507454
rect 504568 507134 504888 507218
rect 504568 506898 504610 507134
rect 504846 506898 504888 507134
rect 504568 506866 504888 506898
rect 514808 507454 515128 507486
rect 514808 507218 514850 507454
rect 515086 507218 515128 507454
rect 514808 507134 515128 507218
rect 514808 506898 514850 507134
rect 515086 506898 515128 507134
rect 514808 506866 515128 506898
rect 525048 507454 525368 507486
rect 525048 507218 525090 507454
rect 525326 507218 525368 507454
rect 525048 507134 525368 507218
rect 525048 506898 525090 507134
rect 525326 506898 525368 507134
rect 525048 506866 525368 506898
rect 535288 507454 535608 507486
rect 535288 507218 535330 507454
rect 535566 507218 535608 507454
rect 535288 507134 535608 507218
rect 535288 506898 535330 507134
rect 535566 506898 535608 507134
rect 535288 506866 535608 506898
rect 28408 489454 28728 489486
rect 28408 489218 28450 489454
rect 28686 489218 28728 489454
rect 28408 489134 28728 489218
rect 28408 488898 28450 489134
rect 28686 488898 28728 489134
rect 28408 488866 28728 488898
rect 38648 489454 38968 489486
rect 38648 489218 38690 489454
rect 38926 489218 38968 489454
rect 38648 489134 38968 489218
rect 38648 488898 38690 489134
rect 38926 488898 38968 489134
rect 38648 488866 38968 488898
rect 48888 489454 49208 489486
rect 48888 489218 48930 489454
rect 49166 489218 49208 489454
rect 48888 489134 49208 489218
rect 48888 488898 48930 489134
rect 49166 488898 49208 489134
rect 48888 488866 49208 488898
rect 59128 489454 59448 489486
rect 59128 489218 59170 489454
rect 59406 489218 59448 489454
rect 59128 489134 59448 489218
rect 59128 488898 59170 489134
rect 59406 488898 59448 489134
rect 59128 488866 59448 488898
rect 69368 489454 69688 489486
rect 69368 489218 69410 489454
rect 69646 489218 69688 489454
rect 69368 489134 69688 489218
rect 69368 488898 69410 489134
rect 69646 488898 69688 489134
rect 69368 488866 69688 488898
rect 79608 489454 79928 489486
rect 79608 489218 79650 489454
rect 79886 489218 79928 489454
rect 79608 489134 79928 489218
rect 79608 488898 79650 489134
rect 79886 488898 79928 489134
rect 79608 488866 79928 488898
rect 89848 489454 90168 489486
rect 89848 489218 89890 489454
rect 90126 489218 90168 489454
rect 89848 489134 90168 489218
rect 89848 488898 89890 489134
rect 90126 488898 90168 489134
rect 89848 488866 90168 488898
rect 100088 489454 100408 489486
rect 100088 489218 100130 489454
rect 100366 489218 100408 489454
rect 100088 489134 100408 489218
rect 100088 488898 100130 489134
rect 100366 488898 100408 489134
rect 100088 488866 100408 488898
rect 110328 489454 110648 489486
rect 110328 489218 110370 489454
rect 110606 489218 110648 489454
rect 110328 489134 110648 489218
rect 110328 488898 110370 489134
rect 110606 488898 110648 489134
rect 110328 488866 110648 488898
rect 120568 489454 120888 489486
rect 120568 489218 120610 489454
rect 120846 489218 120888 489454
rect 120568 489134 120888 489218
rect 120568 488898 120610 489134
rect 120846 488898 120888 489134
rect 120568 488866 120888 488898
rect 130808 489454 131128 489486
rect 130808 489218 130850 489454
rect 131086 489218 131128 489454
rect 130808 489134 131128 489218
rect 130808 488898 130850 489134
rect 131086 488898 131128 489134
rect 130808 488866 131128 488898
rect 141048 489454 141368 489486
rect 141048 489218 141090 489454
rect 141326 489218 141368 489454
rect 141048 489134 141368 489218
rect 141048 488898 141090 489134
rect 141326 488898 141368 489134
rect 141048 488866 141368 488898
rect 151288 489454 151608 489486
rect 151288 489218 151330 489454
rect 151566 489218 151608 489454
rect 151288 489134 151608 489218
rect 151288 488898 151330 489134
rect 151566 488898 151608 489134
rect 151288 488866 151608 488898
rect 161528 489454 161848 489486
rect 161528 489218 161570 489454
rect 161806 489218 161848 489454
rect 161528 489134 161848 489218
rect 161528 488898 161570 489134
rect 161806 488898 161848 489134
rect 161528 488866 161848 488898
rect 171768 489454 172088 489486
rect 171768 489218 171810 489454
rect 172046 489218 172088 489454
rect 171768 489134 172088 489218
rect 171768 488898 171810 489134
rect 172046 488898 172088 489134
rect 171768 488866 172088 488898
rect 182008 489454 182328 489486
rect 182008 489218 182050 489454
rect 182286 489218 182328 489454
rect 182008 489134 182328 489218
rect 182008 488898 182050 489134
rect 182286 488898 182328 489134
rect 182008 488866 182328 488898
rect 192248 489454 192568 489486
rect 192248 489218 192290 489454
rect 192526 489218 192568 489454
rect 192248 489134 192568 489218
rect 192248 488898 192290 489134
rect 192526 488898 192568 489134
rect 192248 488866 192568 488898
rect 202488 489454 202808 489486
rect 202488 489218 202530 489454
rect 202766 489218 202808 489454
rect 202488 489134 202808 489218
rect 202488 488898 202530 489134
rect 202766 488898 202808 489134
rect 202488 488866 202808 488898
rect 212728 489454 213048 489486
rect 212728 489218 212770 489454
rect 213006 489218 213048 489454
rect 212728 489134 213048 489218
rect 212728 488898 212770 489134
rect 213006 488898 213048 489134
rect 212728 488866 213048 488898
rect 222968 489454 223288 489486
rect 222968 489218 223010 489454
rect 223246 489218 223288 489454
rect 222968 489134 223288 489218
rect 222968 488898 223010 489134
rect 223246 488898 223288 489134
rect 222968 488866 223288 488898
rect 233208 489454 233528 489486
rect 233208 489218 233250 489454
rect 233486 489218 233528 489454
rect 233208 489134 233528 489218
rect 233208 488898 233250 489134
rect 233486 488898 233528 489134
rect 233208 488866 233528 488898
rect 243448 489454 243768 489486
rect 243448 489218 243490 489454
rect 243726 489218 243768 489454
rect 243448 489134 243768 489218
rect 243448 488898 243490 489134
rect 243726 488898 243768 489134
rect 243448 488866 243768 488898
rect 253688 489454 254008 489486
rect 253688 489218 253730 489454
rect 253966 489218 254008 489454
rect 253688 489134 254008 489218
rect 253688 488898 253730 489134
rect 253966 488898 254008 489134
rect 253688 488866 254008 488898
rect 263928 489454 264248 489486
rect 263928 489218 263970 489454
rect 264206 489218 264248 489454
rect 263928 489134 264248 489218
rect 263928 488898 263970 489134
rect 264206 488898 264248 489134
rect 263928 488866 264248 488898
rect 274168 489454 274488 489486
rect 274168 489218 274210 489454
rect 274446 489218 274488 489454
rect 274168 489134 274488 489218
rect 274168 488898 274210 489134
rect 274446 488898 274488 489134
rect 274168 488866 274488 488898
rect 284408 489454 284728 489486
rect 284408 489218 284450 489454
rect 284686 489218 284728 489454
rect 284408 489134 284728 489218
rect 284408 488898 284450 489134
rect 284686 488898 284728 489134
rect 284408 488866 284728 488898
rect 294648 489454 294968 489486
rect 294648 489218 294690 489454
rect 294926 489218 294968 489454
rect 294648 489134 294968 489218
rect 294648 488898 294690 489134
rect 294926 488898 294968 489134
rect 294648 488866 294968 488898
rect 304888 489454 305208 489486
rect 304888 489218 304930 489454
rect 305166 489218 305208 489454
rect 304888 489134 305208 489218
rect 304888 488898 304930 489134
rect 305166 488898 305208 489134
rect 304888 488866 305208 488898
rect 315128 489454 315448 489486
rect 315128 489218 315170 489454
rect 315406 489218 315448 489454
rect 315128 489134 315448 489218
rect 315128 488898 315170 489134
rect 315406 488898 315448 489134
rect 315128 488866 315448 488898
rect 325368 489454 325688 489486
rect 325368 489218 325410 489454
rect 325646 489218 325688 489454
rect 325368 489134 325688 489218
rect 325368 488898 325410 489134
rect 325646 488898 325688 489134
rect 325368 488866 325688 488898
rect 335608 489454 335928 489486
rect 335608 489218 335650 489454
rect 335886 489218 335928 489454
rect 335608 489134 335928 489218
rect 335608 488898 335650 489134
rect 335886 488898 335928 489134
rect 335608 488866 335928 488898
rect 345848 489454 346168 489486
rect 345848 489218 345890 489454
rect 346126 489218 346168 489454
rect 345848 489134 346168 489218
rect 345848 488898 345890 489134
rect 346126 488898 346168 489134
rect 345848 488866 346168 488898
rect 356088 489454 356408 489486
rect 356088 489218 356130 489454
rect 356366 489218 356408 489454
rect 356088 489134 356408 489218
rect 356088 488898 356130 489134
rect 356366 488898 356408 489134
rect 356088 488866 356408 488898
rect 366328 489454 366648 489486
rect 366328 489218 366370 489454
rect 366606 489218 366648 489454
rect 366328 489134 366648 489218
rect 366328 488898 366370 489134
rect 366606 488898 366648 489134
rect 366328 488866 366648 488898
rect 376568 489454 376888 489486
rect 376568 489218 376610 489454
rect 376846 489218 376888 489454
rect 376568 489134 376888 489218
rect 376568 488898 376610 489134
rect 376846 488898 376888 489134
rect 376568 488866 376888 488898
rect 386808 489454 387128 489486
rect 386808 489218 386850 489454
rect 387086 489218 387128 489454
rect 386808 489134 387128 489218
rect 386808 488898 386850 489134
rect 387086 488898 387128 489134
rect 386808 488866 387128 488898
rect 397048 489454 397368 489486
rect 397048 489218 397090 489454
rect 397326 489218 397368 489454
rect 397048 489134 397368 489218
rect 397048 488898 397090 489134
rect 397326 488898 397368 489134
rect 397048 488866 397368 488898
rect 407288 489454 407608 489486
rect 407288 489218 407330 489454
rect 407566 489218 407608 489454
rect 407288 489134 407608 489218
rect 407288 488898 407330 489134
rect 407566 488898 407608 489134
rect 407288 488866 407608 488898
rect 417528 489454 417848 489486
rect 417528 489218 417570 489454
rect 417806 489218 417848 489454
rect 417528 489134 417848 489218
rect 417528 488898 417570 489134
rect 417806 488898 417848 489134
rect 417528 488866 417848 488898
rect 427768 489454 428088 489486
rect 427768 489218 427810 489454
rect 428046 489218 428088 489454
rect 427768 489134 428088 489218
rect 427768 488898 427810 489134
rect 428046 488898 428088 489134
rect 427768 488866 428088 488898
rect 438008 489454 438328 489486
rect 438008 489218 438050 489454
rect 438286 489218 438328 489454
rect 438008 489134 438328 489218
rect 438008 488898 438050 489134
rect 438286 488898 438328 489134
rect 438008 488866 438328 488898
rect 448248 489454 448568 489486
rect 448248 489218 448290 489454
rect 448526 489218 448568 489454
rect 448248 489134 448568 489218
rect 448248 488898 448290 489134
rect 448526 488898 448568 489134
rect 448248 488866 448568 488898
rect 458488 489454 458808 489486
rect 458488 489218 458530 489454
rect 458766 489218 458808 489454
rect 458488 489134 458808 489218
rect 458488 488898 458530 489134
rect 458766 488898 458808 489134
rect 458488 488866 458808 488898
rect 468728 489454 469048 489486
rect 468728 489218 468770 489454
rect 469006 489218 469048 489454
rect 468728 489134 469048 489218
rect 468728 488898 468770 489134
rect 469006 488898 469048 489134
rect 468728 488866 469048 488898
rect 478968 489454 479288 489486
rect 478968 489218 479010 489454
rect 479246 489218 479288 489454
rect 478968 489134 479288 489218
rect 478968 488898 479010 489134
rect 479246 488898 479288 489134
rect 478968 488866 479288 488898
rect 489208 489454 489528 489486
rect 489208 489218 489250 489454
rect 489486 489218 489528 489454
rect 489208 489134 489528 489218
rect 489208 488898 489250 489134
rect 489486 488898 489528 489134
rect 489208 488866 489528 488898
rect 499448 489454 499768 489486
rect 499448 489218 499490 489454
rect 499726 489218 499768 489454
rect 499448 489134 499768 489218
rect 499448 488898 499490 489134
rect 499726 488898 499768 489134
rect 499448 488866 499768 488898
rect 509688 489454 510008 489486
rect 509688 489218 509730 489454
rect 509966 489218 510008 489454
rect 509688 489134 510008 489218
rect 509688 488898 509730 489134
rect 509966 488898 510008 489134
rect 509688 488866 510008 488898
rect 519928 489454 520248 489486
rect 519928 489218 519970 489454
rect 520206 489218 520248 489454
rect 519928 489134 520248 489218
rect 519928 488898 519970 489134
rect 520206 488898 520248 489134
rect 519928 488866 520248 488898
rect 530168 489454 530488 489486
rect 530168 489218 530210 489454
rect 530446 489218 530488 489454
rect 530168 489134 530488 489218
rect 530168 488898 530210 489134
rect 530446 488898 530488 489134
rect 530168 488866 530488 488898
rect 15754 474938 15786 475174
rect 16022 474938 16106 475174
rect 16342 474938 16374 475174
rect 15754 474854 16374 474938
rect 15754 474618 15786 474854
rect 16022 474618 16106 474854
rect 16342 474618 16374 474854
rect 15754 439174 16374 474618
rect 541714 478894 542334 514338
rect 541714 478658 541746 478894
rect 541982 478658 542066 478894
rect 542302 478658 542334 478894
rect 541714 478574 542334 478658
rect 541714 478338 541746 478574
rect 541982 478338 542066 478574
rect 542302 478338 542334 478574
rect 23288 471454 23608 471486
rect 23288 471218 23330 471454
rect 23566 471218 23608 471454
rect 23288 471134 23608 471218
rect 23288 470898 23330 471134
rect 23566 470898 23608 471134
rect 23288 470866 23608 470898
rect 33528 471454 33848 471486
rect 33528 471218 33570 471454
rect 33806 471218 33848 471454
rect 33528 471134 33848 471218
rect 33528 470898 33570 471134
rect 33806 470898 33848 471134
rect 33528 470866 33848 470898
rect 43768 471454 44088 471486
rect 43768 471218 43810 471454
rect 44046 471218 44088 471454
rect 43768 471134 44088 471218
rect 43768 470898 43810 471134
rect 44046 470898 44088 471134
rect 43768 470866 44088 470898
rect 54008 471454 54328 471486
rect 54008 471218 54050 471454
rect 54286 471218 54328 471454
rect 54008 471134 54328 471218
rect 54008 470898 54050 471134
rect 54286 470898 54328 471134
rect 54008 470866 54328 470898
rect 64248 471454 64568 471486
rect 64248 471218 64290 471454
rect 64526 471218 64568 471454
rect 64248 471134 64568 471218
rect 64248 470898 64290 471134
rect 64526 470898 64568 471134
rect 64248 470866 64568 470898
rect 74488 471454 74808 471486
rect 74488 471218 74530 471454
rect 74766 471218 74808 471454
rect 74488 471134 74808 471218
rect 74488 470898 74530 471134
rect 74766 470898 74808 471134
rect 74488 470866 74808 470898
rect 84728 471454 85048 471486
rect 84728 471218 84770 471454
rect 85006 471218 85048 471454
rect 84728 471134 85048 471218
rect 84728 470898 84770 471134
rect 85006 470898 85048 471134
rect 84728 470866 85048 470898
rect 94968 471454 95288 471486
rect 94968 471218 95010 471454
rect 95246 471218 95288 471454
rect 94968 471134 95288 471218
rect 94968 470898 95010 471134
rect 95246 470898 95288 471134
rect 94968 470866 95288 470898
rect 105208 471454 105528 471486
rect 105208 471218 105250 471454
rect 105486 471218 105528 471454
rect 105208 471134 105528 471218
rect 105208 470898 105250 471134
rect 105486 470898 105528 471134
rect 105208 470866 105528 470898
rect 115448 471454 115768 471486
rect 115448 471218 115490 471454
rect 115726 471218 115768 471454
rect 115448 471134 115768 471218
rect 115448 470898 115490 471134
rect 115726 470898 115768 471134
rect 115448 470866 115768 470898
rect 125688 471454 126008 471486
rect 125688 471218 125730 471454
rect 125966 471218 126008 471454
rect 125688 471134 126008 471218
rect 125688 470898 125730 471134
rect 125966 470898 126008 471134
rect 125688 470866 126008 470898
rect 135928 471454 136248 471486
rect 135928 471218 135970 471454
rect 136206 471218 136248 471454
rect 135928 471134 136248 471218
rect 135928 470898 135970 471134
rect 136206 470898 136248 471134
rect 135928 470866 136248 470898
rect 146168 471454 146488 471486
rect 146168 471218 146210 471454
rect 146446 471218 146488 471454
rect 146168 471134 146488 471218
rect 146168 470898 146210 471134
rect 146446 470898 146488 471134
rect 146168 470866 146488 470898
rect 156408 471454 156728 471486
rect 156408 471218 156450 471454
rect 156686 471218 156728 471454
rect 156408 471134 156728 471218
rect 156408 470898 156450 471134
rect 156686 470898 156728 471134
rect 156408 470866 156728 470898
rect 166648 471454 166968 471486
rect 166648 471218 166690 471454
rect 166926 471218 166968 471454
rect 166648 471134 166968 471218
rect 166648 470898 166690 471134
rect 166926 470898 166968 471134
rect 166648 470866 166968 470898
rect 176888 471454 177208 471486
rect 176888 471218 176930 471454
rect 177166 471218 177208 471454
rect 176888 471134 177208 471218
rect 176888 470898 176930 471134
rect 177166 470898 177208 471134
rect 176888 470866 177208 470898
rect 187128 471454 187448 471486
rect 187128 471218 187170 471454
rect 187406 471218 187448 471454
rect 187128 471134 187448 471218
rect 187128 470898 187170 471134
rect 187406 470898 187448 471134
rect 187128 470866 187448 470898
rect 197368 471454 197688 471486
rect 197368 471218 197410 471454
rect 197646 471218 197688 471454
rect 197368 471134 197688 471218
rect 197368 470898 197410 471134
rect 197646 470898 197688 471134
rect 197368 470866 197688 470898
rect 207608 471454 207928 471486
rect 207608 471218 207650 471454
rect 207886 471218 207928 471454
rect 207608 471134 207928 471218
rect 207608 470898 207650 471134
rect 207886 470898 207928 471134
rect 207608 470866 207928 470898
rect 217848 471454 218168 471486
rect 217848 471218 217890 471454
rect 218126 471218 218168 471454
rect 217848 471134 218168 471218
rect 217848 470898 217890 471134
rect 218126 470898 218168 471134
rect 217848 470866 218168 470898
rect 228088 471454 228408 471486
rect 228088 471218 228130 471454
rect 228366 471218 228408 471454
rect 228088 471134 228408 471218
rect 228088 470898 228130 471134
rect 228366 470898 228408 471134
rect 228088 470866 228408 470898
rect 238328 471454 238648 471486
rect 238328 471218 238370 471454
rect 238606 471218 238648 471454
rect 238328 471134 238648 471218
rect 238328 470898 238370 471134
rect 238606 470898 238648 471134
rect 238328 470866 238648 470898
rect 248568 471454 248888 471486
rect 248568 471218 248610 471454
rect 248846 471218 248888 471454
rect 248568 471134 248888 471218
rect 248568 470898 248610 471134
rect 248846 470898 248888 471134
rect 248568 470866 248888 470898
rect 258808 471454 259128 471486
rect 258808 471218 258850 471454
rect 259086 471218 259128 471454
rect 258808 471134 259128 471218
rect 258808 470898 258850 471134
rect 259086 470898 259128 471134
rect 258808 470866 259128 470898
rect 269048 471454 269368 471486
rect 269048 471218 269090 471454
rect 269326 471218 269368 471454
rect 269048 471134 269368 471218
rect 269048 470898 269090 471134
rect 269326 470898 269368 471134
rect 269048 470866 269368 470898
rect 279288 471454 279608 471486
rect 279288 471218 279330 471454
rect 279566 471218 279608 471454
rect 279288 471134 279608 471218
rect 279288 470898 279330 471134
rect 279566 470898 279608 471134
rect 279288 470866 279608 470898
rect 289528 471454 289848 471486
rect 289528 471218 289570 471454
rect 289806 471218 289848 471454
rect 289528 471134 289848 471218
rect 289528 470898 289570 471134
rect 289806 470898 289848 471134
rect 289528 470866 289848 470898
rect 299768 471454 300088 471486
rect 299768 471218 299810 471454
rect 300046 471218 300088 471454
rect 299768 471134 300088 471218
rect 299768 470898 299810 471134
rect 300046 470898 300088 471134
rect 299768 470866 300088 470898
rect 310008 471454 310328 471486
rect 310008 471218 310050 471454
rect 310286 471218 310328 471454
rect 310008 471134 310328 471218
rect 310008 470898 310050 471134
rect 310286 470898 310328 471134
rect 310008 470866 310328 470898
rect 320248 471454 320568 471486
rect 320248 471218 320290 471454
rect 320526 471218 320568 471454
rect 320248 471134 320568 471218
rect 320248 470898 320290 471134
rect 320526 470898 320568 471134
rect 320248 470866 320568 470898
rect 330488 471454 330808 471486
rect 330488 471218 330530 471454
rect 330766 471218 330808 471454
rect 330488 471134 330808 471218
rect 330488 470898 330530 471134
rect 330766 470898 330808 471134
rect 330488 470866 330808 470898
rect 340728 471454 341048 471486
rect 340728 471218 340770 471454
rect 341006 471218 341048 471454
rect 340728 471134 341048 471218
rect 340728 470898 340770 471134
rect 341006 470898 341048 471134
rect 340728 470866 341048 470898
rect 350968 471454 351288 471486
rect 350968 471218 351010 471454
rect 351246 471218 351288 471454
rect 350968 471134 351288 471218
rect 350968 470898 351010 471134
rect 351246 470898 351288 471134
rect 350968 470866 351288 470898
rect 361208 471454 361528 471486
rect 361208 471218 361250 471454
rect 361486 471218 361528 471454
rect 361208 471134 361528 471218
rect 361208 470898 361250 471134
rect 361486 470898 361528 471134
rect 361208 470866 361528 470898
rect 371448 471454 371768 471486
rect 371448 471218 371490 471454
rect 371726 471218 371768 471454
rect 371448 471134 371768 471218
rect 371448 470898 371490 471134
rect 371726 470898 371768 471134
rect 371448 470866 371768 470898
rect 381688 471454 382008 471486
rect 381688 471218 381730 471454
rect 381966 471218 382008 471454
rect 381688 471134 382008 471218
rect 381688 470898 381730 471134
rect 381966 470898 382008 471134
rect 381688 470866 382008 470898
rect 391928 471454 392248 471486
rect 391928 471218 391970 471454
rect 392206 471218 392248 471454
rect 391928 471134 392248 471218
rect 391928 470898 391970 471134
rect 392206 470898 392248 471134
rect 391928 470866 392248 470898
rect 402168 471454 402488 471486
rect 402168 471218 402210 471454
rect 402446 471218 402488 471454
rect 402168 471134 402488 471218
rect 402168 470898 402210 471134
rect 402446 470898 402488 471134
rect 402168 470866 402488 470898
rect 412408 471454 412728 471486
rect 412408 471218 412450 471454
rect 412686 471218 412728 471454
rect 412408 471134 412728 471218
rect 412408 470898 412450 471134
rect 412686 470898 412728 471134
rect 412408 470866 412728 470898
rect 422648 471454 422968 471486
rect 422648 471218 422690 471454
rect 422926 471218 422968 471454
rect 422648 471134 422968 471218
rect 422648 470898 422690 471134
rect 422926 470898 422968 471134
rect 422648 470866 422968 470898
rect 432888 471454 433208 471486
rect 432888 471218 432930 471454
rect 433166 471218 433208 471454
rect 432888 471134 433208 471218
rect 432888 470898 432930 471134
rect 433166 470898 433208 471134
rect 432888 470866 433208 470898
rect 443128 471454 443448 471486
rect 443128 471218 443170 471454
rect 443406 471218 443448 471454
rect 443128 471134 443448 471218
rect 443128 470898 443170 471134
rect 443406 470898 443448 471134
rect 443128 470866 443448 470898
rect 453368 471454 453688 471486
rect 453368 471218 453410 471454
rect 453646 471218 453688 471454
rect 453368 471134 453688 471218
rect 453368 470898 453410 471134
rect 453646 470898 453688 471134
rect 453368 470866 453688 470898
rect 463608 471454 463928 471486
rect 463608 471218 463650 471454
rect 463886 471218 463928 471454
rect 463608 471134 463928 471218
rect 463608 470898 463650 471134
rect 463886 470898 463928 471134
rect 463608 470866 463928 470898
rect 473848 471454 474168 471486
rect 473848 471218 473890 471454
rect 474126 471218 474168 471454
rect 473848 471134 474168 471218
rect 473848 470898 473890 471134
rect 474126 470898 474168 471134
rect 473848 470866 474168 470898
rect 484088 471454 484408 471486
rect 484088 471218 484130 471454
rect 484366 471218 484408 471454
rect 484088 471134 484408 471218
rect 484088 470898 484130 471134
rect 484366 470898 484408 471134
rect 484088 470866 484408 470898
rect 494328 471454 494648 471486
rect 494328 471218 494370 471454
rect 494606 471218 494648 471454
rect 494328 471134 494648 471218
rect 494328 470898 494370 471134
rect 494606 470898 494648 471134
rect 494328 470866 494648 470898
rect 504568 471454 504888 471486
rect 504568 471218 504610 471454
rect 504846 471218 504888 471454
rect 504568 471134 504888 471218
rect 504568 470898 504610 471134
rect 504846 470898 504888 471134
rect 504568 470866 504888 470898
rect 514808 471454 515128 471486
rect 514808 471218 514850 471454
rect 515086 471218 515128 471454
rect 514808 471134 515128 471218
rect 514808 470898 514850 471134
rect 515086 470898 515128 471134
rect 514808 470866 515128 470898
rect 525048 471454 525368 471486
rect 525048 471218 525090 471454
rect 525326 471218 525368 471454
rect 525048 471134 525368 471218
rect 525048 470898 525090 471134
rect 525326 470898 525368 471134
rect 525048 470866 525368 470898
rect 535288 471454 535608 471486
rect 535288 471218 535330 471454
rect 535566 471218 535608 471454
rect 535288 471134 535608 471218
rect 535288 470898 535330 471134
rect 535566 470898 535608 471134
rect 535288 470866 535608 470898
rect 28408 453454 28728 453486
rect 28408 453218 28450 453454
rect 28686 453218 28728 453454
rect 28408 453134 28728 453218
rect 28408 452898 28450 453134
rect 28686 452898 28728 453134
rect 28408 452866 28728 452898
rect 38648 453454 38968 453486
rect 38648 453218 38690 453454
rect 38926 453218 38968 453454
rect 38648 453134 38968 453218
rect 38648 452898 38690 453134
rect 38926 452898 38968 453134
rect 38648 452866 38968 452898
rect 48888 453454 49208 453486
rect 48888 453218 48930 453454
rect 49166 453218 49208 453454
rect 48888 453134 49208 453218
rect 48888 452898 48930 453134
rect 49166 452898 49208 453134
rect 48888 452866 49208 452898
rect 59128 453454 59448 453486
rect 59128 453218 59170 453454
rect 59406 453218 59448 453454
rect 59128 453134 59448 453218
rect 59128 452898 59170 453134
rect 59406 452898 59448 453134
rect 59128 452866 59448 452898
rect 69368 453454 69688 453486
rect 69368 453218 69410 453454
rect 69646 453218 69688 453454
rect 69368 453134 69688 453218
rect 69368 452898 69410 453134
rect 69646 452898 69688 453134
rect 69368 452866 69688 452898
rect 79608 453454 79928 453486
rect 79608 453218 79650 453454
rect 79886 453218 79928 453454
rect 79608 453134 79928 453218
rect 79608 452898 79650 453134
rect 79886 452898 79928 453134
rect 79608 452866 79928 452898
rect 89848 453454 90168 453486
rect 89848 453218 89890 453454
rect 90126 453218 90168 453454
rect 89848 453134 90168 453218
rect 89848 452898 89890 453134
rect 90126 452898 90168 453134
rect 89848 452866 90168 452898
rect 100088 453454 100408 453486
rect 100088 453218 100130 453454
rect 100366 453218 100408 453454
rect 100088 453134 100408 453218
rect 100088 452898 100130 453134
rect 100366 452898 100408 453134
rect 100088 452866 100408 452898
rect 110328 453454 110648 453486
rect 110328 453218 110370 453454
rect 110606 453218 110648 453454
rect 110328 453134 110648 453218
rect 110328 452898 110370 453134
rect 110606 452898 110648 453134
rect 110328 452866 110648 452898
rect 120568 453454 120888 453486
rect 120568 453218 120610 453454
rect 120846 453218 120888 453454
rect 120568 453134 120888 453218
rect 120568 452898 120610 453134
rect 120846 452898 120888 453134
rect 120568 452866 120888 452898
rect 130808 453454 131128 453486
rect 130808 453218 130850 453454
rect 131086 453218 131128 453454
rect 130808 453134 131128 453218
rect 130808 452898 130850 453134
rect 131086 452898 131128 453134
rect 130808 452866 131128 452898
rect 141048 453454 141368 453486
rect 141048 453218 141090 453454
rect 141326 453218 141368 453454
rect 141048 453134 141368 453218
rect 141048 452898 141090 453134
rect 141326 452898 141368 453134
rect 141048 452866 141368 452898
rect 151288 453454 151608 453486
rect 151288 453218 151330 453454
rect 151566 453218 151608 453454
rect 151288 453134 151608 453218
rect 151288 452898 151330 453134
rect 151566 452898 151608 453134
rect 151288 452866 151608 452898
rect 161528 453454 161848 453486
rect 161528 453218 161570 453454
rect 161806 453218 161848 453454
rect 161528 453134 161848 453218
rect 161528 452898 161570 453134
rect 161806 452898 161848 453134
rect 161528 452866 161848 452898
rect 171768 453454 172088 453486
rect 171768 453218 171810 453454
rect 172046 453218 172088 453454
rect 171768 453134 172088 453218
rect 171768 452898 171810 453134
rect 172046 452898 172088 453134
rect 171768 452866 172088 452898
rect 182008 453454 182328 453486
rect 182008 453218 182050 453454
rect 182286 453218 182328 453454
rect 182008 453134 182328 453218
rect 182008 452898 182050 453134
rect 182286 452898 182328 453134
rect 182008 452866 182328 452898
rect 192248 453454 192568 453486
rect 192248 453218 192290 453454
rect 192526 453218 192568 453454
rect 192248 453134 192568 453218
rect 192248 452898 192290 453134
rect 192526 452898 192568 453134
rect 192248 452866 192568 452898
rect 202488 453454 202808 453486
rect 202488 453218 202530 453454
rect 202766 453218 202808 453454
rect 202488 453134 202808 453218
rect 202488 452898 202530 453134
rect 202766 452898 202808 453134
rect 202488 452866 202808 452898
rect 212728 453454 213048 453486
rect 212728 453218 212770 453454
rect 213006 453218 213048 453454
rect 212728 453134 213048 453218
rect 212728 452898 212770 453134
rect 213006 452898 213048 453134
rect 212728 452866 213048 452898
rect 222968 453454 223288 453486
rect 222968 453218 223010 453454
rect 223246 453218 223288 453454
rect 222968 453134 223288 453218
rect 222968 452898 223010 453134
rect 223246 452898 223288 453134
rect 222968 452866 223288 452898
rect 233208 453454 233528 453486
rect 233208 453218 233250 453454
rect 233486 453218 233528 453454
rect 233208 453134 233528 453218
rect 233208 452898 233250 453134
rect 233486 452898 233528 453134
rect 233208 452866 233528 452898
rect 243448 453454 243768 453486
rect 243448 453218 243490 453454
rect 243726 453218 243768 453454
rect 243448 453134 243768 453218
rect 243448 452898 243490 453134
rect 243726 452898 243768 453134
rect 243448 452866 243768 452898
rect 253688 453454 254008 453486
rect 253688 453218 253730 453454
rect 253966 453218 254008 453454
rect 253688 453134 254008 453218
rect 253688 452898 253730 453134
rect 253966 452898 254008 453134
rect 253688 452866 254008 452898
rect 263928 453454 264248 453486
rect 263928 453218 263970 453454
rect 264206 453218 264248 453454
rect 263928 453134 264248 453218
rect 263928 452898 263970 453134
rect 264206 452898 264248 453134
rect 263928 452866 264248 452898
rect 274168 453454 274488 453486
rect 274168 453218 274210 453454
rect 274446 453218 274488 453454
rect 274168 453134 274488 453218
rect 274168 452898 274210 453134
rect 274446 452898 274488 453134
rect 274168 452866 274488 452898
rect 284408 453454 284728 453486
rect 284408 453218 284450 453454
rect 284686 453218 284728 453454
rect 284408 453134 284728 453218
rect 284408 452898 284450 453134
rect 284686 452898 284728 453134
rect 284408 452866 284728 452898
rect 294648 453454 294968 453486
rect 294648 453218 294690 453454
rect 294926 453218 294968 453454
rect 294648 453134 294968 453218
rect 294648 452898 294690 453134
rect 294926 452898 294968 453134
rect 294648 452866 294968 452898
rect 304888 453454 305208 453486
rect 304888 453218 304930 453454
rect 305166 453218 305208 453454
rect 304888 453134 305208 453218
rect 304888 452898 304930 453134
rect 305166 452898 305208 453134
rect 304888 452866 305208 452898
rect 315128 453454 315448 453486
rect 315128 453218 315170 453454
rect 315406 453218 315448 453454
rect 315128 453134 315448 453218
rect 315128 452898 315170 453134
rect 315406 452898 315448 453134
rect 315128 452866 315448 452898
rect 325368 453454 325688 453486
rect 325368 453218 325410 453454
rect 325646 453218 325688 453454
rect 325368 453134 325688 453218
rect 325368 452898 325410 453134
rect 325646 452898 325688 453134
rect 325368 452866 325688 452898
rect 335608 453454 335928 453486
rect 335608 453218 335650 453454
rect 335886 453218 335928 453454
rect 335608 453134 335928 453218
rect 335608 452898 335650 453134
rect 335886 452898 335928 453134
rect 335608 452866 335928 452898
rect 345848 453454 346168 453486
rect 345848 453218 345890 453454
rect 346126 453218 346168 453454
rect 345848 453134 346168 453218
rect 345848 452898 345890 453134
rect 346126 452898 346168 453134
rect 345848 452866 346168 452898
rect 356088 453454 356408 453486
rect 356088 453218 356130 453454
rect 356366 453218 356408 453454
rect 356088 453134 356408 453218
rect 356088 452898 356130 453134
rect 356366 452898 356408 453134
rect 356088 452866 356408 452898
rect 366328 453454 366648 453486
rect 366328 453218 366370 453454
rect 366606 453218 366648 453454
rect 366328 453134 366648 453218
rect 366328 452898 366370 453134
rect 366606 452898 366648 453134
rect 366328 452866 366648 452898
rect 376568 453454 376888 453486
rect 376568 453218 376610 453454
rect 376846 453218 376888 453454
rect 376568 453134 376888 453218
rect 376568 452898 376610 453134
rect 376846 452898 376888 453134
rect 376568 452866 376888 452898
rect 386808 453454 387128 453486
rect 386808 453218 386850 453454
rect 387086 453218 387128 453454
rect 386808 453134 387128 453218
rect 386808 452898 386850 453134
rect 387086 452898 387128 453134
rect 386808 452866 387128 452898
rect 397048 453454 397368 453486
rect 397048 453218 397090 453454
rect 397326 453218 397368 453454
rect 397048 453134 397368 453218
rect 397048 452898 397090 453134
rect 397326 452898 397368 453134
rect 397048 452866 397368 452898
rect 407288 453454 407608 453486
rect 407288 453218 407330 453454
rect 407566 453218 407608 453454
rect 407288 453134 407608 453218
rect 407288 452898 407330 453134
rect 407566 452898 407608 453134
rect 407288 452866 407608 452898
rect 417528 453454 417848 453486
rect 417528 453218 417570 453454
rect 417806 453218 417848 453454
rect 417528 453134 417848 453218
rect 417528 452898 417570 453134
rect 417806 452898 417848 453134
rect 417528 452866 417848 452898
rect 427768 453454 428088 453486
rect 427768 453218 427810 453454
rect 428046 453218 428088 453454
rect 427768 453134 428088 453218
rect 427768 452898 427810 453134
rect 428046 452898 428088 453134
rect 427768 452866 428088 452898
rect 438008 453454 438328 453486
rect 438008 453218 438050 453454
rect 438286 453218 438328 453454
rect 438008 453134 438328 453218
rect 438008 452898 438050 453134
rect 438286 452898 438328 453134
rect 438008 452866 438328 452898
rect 448248 453454 448568 453486
rect 448248 453218 448290 453454
rect 448526 453218 448568 453454
rect 448248 453134 448568 453218
rect 448248 452898 448290 453134
rect 448526 452898 448568 453134
rect 448248 452866 448568 452898
rect 458488 453454 458808 453486
rect 458488 453218 458530 453454
rect 458766 453218 458808 453454
rect 458488 453134 458808 453218
rect 458488 452898 458530 453134
rect 458766 452898 458808 453134
rect 458488 452866 458808 452898
rect 468728 453454 469048 453486
rect 468728 453218 468770 453454
rect 469006 453218 469048 453454
rect 468728 453134 469048 453218
rect 468728 452898 468770 453134
rect 469006 452898 469048 453134
rect 468728 452866 469048 452898
rect 478968 453454 479288 453486
rect 478968 453218 479010 453454
rect 479246 453218 479288 453454
rect 478968 453134 479288 453218
rect 478968 452898 479010 453134
rect 479246 452898 479288 453134
rect 478968 452866 479288 452898
rect 489208 453454 489528 453486
rect 489208 453218 489250 453454
rect 489486 453218 489528 453454
rect 489208 453134 489528 453218
rect 489208 452898 489250 453134
rect 489486 452898 489528 453134
rect 489208 452866 489528 452898
rect 499448 453454 499768 453486
rect 499448 453218 499490 453454
rect 499726 453218 499768 453454
rect 499448 453134 499768 453218
rect 499448 452898 499490 453134
rect 499726 452898 499768 453134
rect 499448 452866 499768 452898
rect 509688 453454 510008 453486
rect 509688 453218 509730 453454
rect 509966 453218 510008 453454
rect 509688 453134 510008 453218
rect 509688 452898 509730 453134
rect 509966 452898 510008 453134
rect 509688 452866 510008 452898
rect 519928 453454 520248 453486
rect 519928 453218 519970 453454
rect 520206 453218 520248 453454
rect 519928 453134 520248 453218
rect 519928 452898 519970 453134
rect 520206 452898 520248 453134
rect 519928 452866 520248 452898
rect 530168 453454 530488 453486
rect 530168 453218 530210 453454
rect 530446 453218 530488 453454
rect 530168 453134 530488 453218
rect 530168 452898 530210 453134
rect 530446 452898 530488 453134
rect 530168 452866 530488 452898
rect 15754 438938 15786 439174
rect 16022 438938 16106 439174
rect 16342 438938 16374 439174
rect 15754 438854 16374 438938
rect 15754 438618 15786 438854
rect 16022 438618 16106 438854
rect 16342 438618 16374 438854
rect 15754 403174 16374 438618
rect 541714 442894 542334 478338
rect 541714 442658 541746 442894
rect 541982 442658 542066 442894
rect 542302 442658 542334 442894
rect 541714 442574 542334 442658
rect 541714 442338 541746 442574
rect 541982 442338 542066 442574
rect 542302 442338 542334 442574
rect 23288 435454 23608 435486
rect 23288 435218 23330 435454
rect 23566 435218 23608 435454
rect 23288 435134 23608 435218
rect 23288 434898 23330 435134
rect 23566 434898 23608 435134
rect 23288 434866 23608 434898
rect 33528 435454 33848 435486
rect 33528 435218 33570 435454
rect 33806 435218 33848 435454
rect 33528 435134 33848 435218
rect 33528 434898 33570 435134
rect 33806 434898 33848 435134
rect 33528 434866 33848 434898
rect 43768 435454 44088 435486
rect 43768 435218 43810 435454
rect 44046 435218 44088 435454
rect 43768 435134 44088 435218
rect 43768 434898 43810 435134
rect 44046 434898 44088 435134
rect 43768 434866 44088 434898
rect 54008 435454 54328 435486
rect 54008 435218 54050 435454
rect 54286 435218 54328 435454
rect 54008 435134 54328 435218
rect 54008 434898 54050 435134
rect 54286 434898 54328 435134
rect 54008 434866 54328 434898
rect 64248 435454 64568 435486
rect 64248 435218 64290 435454
rect 64526 435218 64568 435454
rect 64248 435134 64568 435218
rect 64248 434898 64290 435134
rect 64526 434898 64568 435134
rect 64248 434866 64568 434898
rect 74488 435454 74808 435486
rect 74488 435218 74530 435454
rect 74766 435218 74808 435454
rect 74488 435134 74808 435218
rect 74488 434898 74530 435134
rect 74766 434898 74808 435134
rect 74488 434866 74808 434898
rect 84728 435454 85048 435486
rect 84728 435218 84770 435454
rect 85006 435218 85048 435454
rect 84728 435134 85048 435218
rect 84728 434898 84770 435134
rect 85006 434898 85048 435134
rect 84728 434866 85048 434898
rect 94968 435454 95288 435486
rect 94968 435218 95010 435454
rect 95246 435218 95288 435454
rect 94968 435134 95288 435218
rect 94968 434898 95010 435134
rect 95246 434898 95288 435134
rect 94968 434866 95288 434898
rect 105208 435454 105528 435486
rect 105208 435218 105250 435454
rect 105486 435218 105528 435454
rect 105208 435134 105528 435218
rect 105208 434898 105250 435134
rect 105486 434898 105528 435134
rect 105208 434866 105528 434898
rect 115448 435454 115768 435486
rect 115448 435218 115490 435454
rect 115726 435218 115768 435454
rect 115448 435134 115768 435218
rect 115448 434898 115490 435134
rect 115726 434898 115768 435134
rect 115448 434866 115768 434898
rect 125688 435454 126008 435486
rect 125688 435218 125730 435454
rect 125966 435218 126008 435454
rect 125688 435134 126008 435218
rect 125688 434898 125730 435134
rect 125966 434898 126008 435134
rect 125688 434866 126008 434898
rect 135928 435454 136248 435486
rect 135928 435218 135970 435454
rect 136206 435218 136248 435454
rect 135928 435134 136248 435218
rect 135928 434898 135970 435134
rect 136206 434898 136248 435134
rect 135928 434866 136248 434898
rect 146168 435454 146488 435486
rect 146168 435218 146210 435454
rect 146446 435218 146488 435454
rect 146168 435134 146488 435218
rect 146168 434898 146210 435134
rect 146446 434898 146488 435134
rect 146168 434866 146488 434898
rect 156408 435454 156728 435486
rect 156408 435218 156450 435454
rect 156686 435218 156728 435454
rect 156408 435134 156728 435218
rect 156408 434898 156450 435134
rect 156686 434898 156728 435134
rect 156408 434866 156728 434898
rect 166648 435454 166968 435486
rect 166648 435218 166690 435454
rect 166926 435218 166968 435454
rect 166648 435134 166968 435218
rect 166648 434898 166690 435134
rect 166926 434898 166968 435134
rect 166648 434866 166968 434898
rect 176888 435454 177208 435486
rect 176888 435218 176930 435454
rect 177166 435218 177208 435454
rect 176888 435134 177208 435218
rect 176888 434898 176930 435134
rect 177166 434898 177208 435134
rect 176888 434866 177208 434898
rect 187128 435454 187448 435486
rect 187128 435218 187170 435454
rect 187406 435218 187448 435454
rect 187128 435134 187448 435218
rect 187128 434898 187170 435134
rect 187406 434898 187448 435134
rect 187128 434866 187448 434898
rect 197368 435454 197688 435486
rect 197368 435218 197410 435454
rect 197646 435218 197688 435454
rect 197368 435134 197688 435218
rect 197368 434898 197410 435134
rect 197646 434898 197688 435134
rect 197368 434866 197688 434898
rect 207608 435454 207928 435486
rect 207608 435218 207650 435454
rect 207886 435218 207928 435454
rect 207608 435134 207928 435218
rect 207608 434898 207650 435134
rect 207886 434898 207928 435134
rect 207608 434866 207928 434898
rect 217848 435454 218168 435486
rect 217848 435218 217890 435454
rect 218126 435218 218168 435454
rect 217848 435134 218168 435218
rect 217848 434898 217890 435134
rect 218126 434898 218168 435134
rect 217848 434866 218168 434898
rect 228088 435454 228408 435486
rect 228088 435218 228130 435454
rect 228366 435218 228408 435454
rect 228088 435134 228408 435218
rect 228088 434898 228130 435134
rect 228366 434898 228408 435134
rect 228088 434866 228408 434898
rect 238328 435454 238648 435486
rect 238328 435218 238370 435454
rect 238606 435218 238648 435454
rect 238328 435134 238648 435218
rect 238328 434898 238370 435134
rect 238606 434898 238648 435134
rect 238328 434866 238648 434898
rect 248568 435454 248888 435486
rect 248568 435218 248610 435454
rect 248846 435218 248888 435454
rect 248568 435134 248888 435218
rect 248568 434898 248610 435134
rect 248846 434898 248888 435134
rect 248568 434866 248888 434898
rect 258808 435454 259128 435486
rect 258808 435218 258850 435454
rect 259086 435218 259128 435454
rect 258808 435134 259128 435218
rect 258808 434898 258850 435134
rect 259086 434898 259128 435134
rect 258808 434866 259128 434898
rect 269048 435454 269368 435486
rect 269048 435218 269090 435454
rect 269326 435218 269368 435454
rect 269048 435134 269368 435218
rect 269048 434898 269090 435134
rect 269326 434898 269368 435134
rect 269048 434866 269368 434898
rect 279288 435454 279608 435486
rect 279288 435218 279330 435454
rect 279566 435218 279608 435454
rect 279288 435134 279608 435218
rect 279288 434898 279330 435134
rect 279566 434898 279608 435134
rect 279288 434866 279608 434898
rect 289528 435454 289848 435486
rect 289528 435218 289570 435454
rect 289806 435218 289848 435454
rect 289528 435134 289848 435218
rect 289528 434898 289570 435134
rect 289806 434898 289848 435134
rect 289528 434866 289848 434898
rect 299768 435454 300088 435486
rect 299768 435218 299810 435454
rect 300046 435218 300088 435454
rect 299768 435134 300088 435218
rect 299768 434898 299810 435134
rect 300046 434898 300088 435134
rect 299768 434866 300088 434898
rect 310008 435454 310328 435486
rect 310008 435218 310050 435454
rect 310286 435218 310328 435454
rect 310008 435134 310328 435218
rect 310008 434898 310050 435134
rect 310286 434898 310328 435134
rect 310008 434866 310328 434898
rect 320248 435454 320568 435486
rect 320248 435218 320290 435454
rect 320526 435218 320568 435454
rect 320248 435134 320568 435218
rect 320248 434898 320290 435134
rect 320526 434898 320568 435134
rect 320248 434866 320568 434898
rect 330488 435454 330808 435486
rect 330488 435218 330530 435454
rect 330766 435218 330808 435454
rect 330488 435134 330808 435218
rect 330488 434898 330530 435134
rect 330766 434898 330808 435134
rect 330488 434866 330808 434898
rect 340728 435454 341048 435486
rect 340728 435218 340770 435454
rect 341006 435218 341048 435454
rect 340728 435134 341048 435218
rect 340728 434898 340770 435134
rect 341006 434898 341048 435134
rect 340728 434866 341048 434898
rect 350968 435454 351288 435486
rect 350968 435218 351010 435454
rect 351246 435218 351288 435454
rect 350968 435134 351288 435218
rect 350968 434898 351010 435134
rect 351246 434898 351288 435134
rect 350968 434866 351288 434898
rect 361208 435454 361528 435486
rect 361208 435218 361250 435454
rect 361486 435218 361528 435454
rect 361208 435134 361528 435218
rect 361208 434898 361250 435134
rect 361486 434898 361528 435134
rect 361208 434866 361528 434898
rect 371448 435454 371768 435486
rect 371448 435218 371490 435454
rect 371726 435218 371768 435454
rect 371448 435134 371768 435218
rect 371448 434898 371490 435134
rect 371726 434898 371768 435134
rect 371448 434866 371768 434898
rect 381688 435454 382008 435486
rect 381688 435218 381730 435454
rect 381966 435218 382008 435454
rect 381688 435134 382008 435218
rect 381688 434898 381730 435134
rect 381966 434898 382008 435134
rect 381688 434866 382008 434898
rect 391928 435454 392248 435486
rect 391928 435218 391970 435454
rect 392206 435218 392248 435454
rect 391928 435134 392248 435218
rect 391928 434898 391970 435134
rect 392206 434898 392248 435134
rect 391928 434866 392248 434898
rect 402168 435454 402488 435486
rect 402168 435218 402210 435454
rect 402446 435218 402488 435454
rect 402168 435134 402488 435218
rect 402168 434898 402210 435134
rect 402446 434898 402488 435134
rect 402168 434866 402488 434898
rect 412408 435454 412728 435486
rect 412408 435218 412450 435454
rect 412686 435218 412728 435454
rect 412408 435134 412728 435218
rect 412408 434898 412450 435134
rect 412686 434898 412728 435134
rect 412408 434866 412728 434898
rect 422648 435454 422968 435486
rect 422648 435218 422690 435454
rect 422926 435218 422968 435454
rect 422648 435134 422968 435218
rect 422648 434898 422690 435134
rect 422926 434898 422968 435134
rect 422648 434866 422968 434898
rect 432888 435454 433208 435486
rect 432888 435218 432930 435454
rect 433166 435218 433208 435454
rect 432888 435134 433208 435218
rect 432888 434898 432930 435134
rect 433166 434898 433208 435134
rect 432888 434866 433208 434898
rect 443128 435454 443448 435486
rect 443128 435218 443170 435454
rect 443406 435218 443448 435454
rect 443128 435134 443448 435218
rect 443128 434898 443170 435134
rect 443406 434898 443448 435134
rect 443128 434866 443448 434898
rect 453368 435454 453688 435486
rect 453368 435218 453410 435454
rect 453646 435218 453688 435454
rect 453368 435134 453688 435218
rect 453368 434898 453410 435134
rect 453646 434898 453688 435134
rect 453368 434866 453688 434898
rect 463608 435454 463928 435486
rect 463608 435218 463650 435454
rect 463886 435218 463928 435454
rect 463608 435134 463928 435218
rect 463608 434898 463650 435134
rect 463886 434898 463928 435134
rect 463608 434866 463928 434898
rect 473848 435454 474168 435486
rect 473848 435218 473890 435454
rect 474126 435218 474168 435454
rect 473848 435134 474168 435218
rect 473848 434898 473890 435134
rect 474126 434898 474168 435134
rect 473848 434866 474168 434898
rect 484088 435454 484408 435486
rect 484088 435218 484130 435454
rect 484366 435218 484408 435454
rect 484088 435134 484408 435218
rect 484088 434898 484130 435134
rect 484366 434898 484408 435134
rect 484088 434866 484408 434898
rect 494328 435454 494648 435486
rect 494328 435218 494370 435454
rect 494606 435218 494648 435454
rect 494328 435134 494648 435218
rect 494328 434898 494370 435134
rect 494606 434898 494648 435134
rect 494328 434866 494648 434898
rect 504568 435454 504888 435486
rect 504568 435218 504610 435454
rect 504846 435218 504888 435454
rect 504568 435134 504888 435218
rect 504568 434898 504610 435134
rect 504846 434898 504888 435134
rect 504568 434866 504888 434898
rect 514808 435454 515128 435486
rect 514808 435218 514850 435454
rect 515086 435218 515128 435454
rect 514808 435134 515128 435218
rect 514808 434898 514850 435134
rect 515086 434898 515128 435134
rect 514808 434866 515128 434898
rect 525048 435454 525368 435486
rect 525048 435218 525090 435454
rect 525326 435218 525368 435454
rect 525048 435134 525368 435218
rect 525048 434898 525090 435134
rect 525326 434898 525368 435134
rect 525048 434866 525368 434898
rect 535288 435454 535608 435486
rect 535288 435218 535330 435454
rect 535566 435218 535608 435454
rect 535288 435134 535608 435218
rect 535288 434898 535330 435134
rect 535566 434898 535608 435134
rect 535288 434866 535608 434898
rect 28408 417454 28728 417486
rect 28408 417218 28450 417454
rect 28686 417218 28728 417454
rect 28408 417134 28728 417218
rect 28408 416898 28450 417134
rect 28686 416898 28728 417134
rect 28408 416866 28728 416898
rect 38648 417454 38968 417486
rect 38648 417218 38690 417454
rect 38926 417218 38968 417454
rect 38648 417134 38968 417218
rect 38648 416898 38690 417134
rect 38926 416898 38968 417134
rect 38648 416866 38968 416898
rect 48888 417454 49208 417486
rect 48888 417218 48930 417454
rect 49166 417218 49208 417454
rect 48888 417134 49208 417218
rect 48888 416898 48930 417134
rect 49166 416898 49208 417134
rect 48888 416866 49208 416898
rect 59128 417454 59448 417486
rect 59128 417218 59170 417454
rect 59406 417218 59448 417454
rect 59128 417134 59448 417218
rect 59128 416898 59170 417134
rect 59406 416898 59448 417134
rect 59128 416866 59448 416898
rect 69368 417454 69688 417486
rect 69368 417218 69410 417454
rect 69646 417218 69688 417454
rect 69368 417134 69688 417218
rect 69368 416898 69410 417134
rect 69646 416898 69688 417134
rect 69368 416866 69688 416898
rect 79608 417454 79928 417486
rect 79608 417218 79650 417454
rect 79886 417218 79928 417454
rect 79608 417134 79928 417218
rect 79608 416898 79650 417134
rect 79886 416898 79928 417134
rect 79608 416866 79928 416898
rect 89848 417454 90168 417486
rect 89848 417218 89890 417454
rect 90126 417218 90168 417454
rect 89848 417134 90168 417218
rect 89848 416898 89890 417134
rect 90126 416898 90168 417134
rect 89848 416866 90168 416898
rect 100088 417454 100408 417486
rect 100088 417218 100130 417454
rect 100366 417218 100408 417454
rect 100088 417134 100408 417218
rect 100088 416898 100130 417134
rect 100366 416898 100408 417134
rect 100088 416866 100408 416898
rect 110328 417454 110648 417486
rect 110328 417218 110370 417454
rect 110606 417218 110648 417454
rect 110328 417134 110648 417218
rect 110328 416898 110370 417134
rect 110606 416898 110648 417134
rect 110328 416866 110648 416898
rect 120568 417454 120888 417486
rect 120568 417218 120610 417454
rect 120846 417218 120888 417454
rect 120568 417134 120888 417218
rect 120568 416898 120610 417134
rect 120846 416898 120888 417134
rect 120568 416866 120888 416898
rect 130808 417454 131128 417486
rect 130808 417218 130850 417454
rect 131086 417218 131128 417454
rect 130808 417134 131128 417218
rect 130808 416898 130850 417134
rect 131086 416898 131128 417134
rect 130808 416866 131128 416898
rect 141048 417454 141368 417486
rect 141048 417218 141090 417454
rect 141326 417218 141368 417454
rect 141048 417134 141368 417218
rect 141048 416898 141090 417134
rect 141326 416898 141368 417134
rect 141048 416866 141368 416898
rect 151288 417454 151608 417486
rect 151288 417218 151330 417454
rect 151566 417218 151608 417454
rect 151288 417134 151608 417218
rect 151288 416898 151330 417134
rect 151566 416898 151608 417134
rect 151288 416866 151608 416898
rect 161528 417454 161848 417486
rect 161528 417218 161570 417454
rect 161806 417218 161848 417454
rect 161528 417134 161848 417218
rect 161528 416898 161570 417134
rect 161806 416898 161848 417134
rect 161528 416866 161848 416898
rect 171768 417454 172088 417486
rect 171768 417218 171810 417454
rect 172046 417218 172088 417454
rect 171768 417134 172088 417218
rect 171768 416898 171810 417134
rect 172046 416898 172088 417134
rect 171768 416866 172088 416898
rect 182008 417454 182328 417486
rect 182008 417218 182050 417454
rect 182286 417218 182328 417454
rect 182008 417134 182328 417218
rect 182008 416898 182050 417134
rect 182286 416898 182328 417134
rect 182008 416866 182328 416898
rect 192248 417454 192568 417486
rect 192248 417218 192290 417454
rect 192526 417218 192568 417454
rect 192248 417134 192568 417218
rect 192248 416898 192290 417134
rect 192526 416898 192568 417134
rect 192248 416866 192568 416898
rect 202488 417454 202808 417486
rect 202488 417218 202530 417454
rect 202766 417218 202808 417454
rect 202488 417134 202808 417218
rect 202488 416898 202530 417134
rect 202766 416898 202808 417134
rect 202488 416866 202808 416898
rect 212728 417454 213048 417486
rect 212728 417218 212770 417454
rect 213006 417218 213048 417454
rect 212728 417134 213048 417218
rect 212728 416898 212770 417134
rect 213006 416898 213048 417134
rect 212728 416866 213048 416898
rect 222968 417454 223288 417486
rect 222968 417218 223010 417454
rect 223246 417218 223288 417454
rect 222968 417134 223288 417218
rect 222968 416898 223010 417134
rect 223246 416898 223288 417134
rect 222968 416866 223288 416898
rect 233208 417454 233528 417486
rect 233208 417218 233250 417454
rect 233486 417218 233528 417454
rect 233208 417134 233528 417218
rect 233208 416898 233250 417134
rect 233486 416898 233528 417134
rect 233208 416866 233528 416898
rect 243448 417454 243768 417486
rect 243448 417218 243490 417454
rect 243726 417218 243768 417454
rect 243448 417134 243768 417218
rect 243448 416898 243490 417134
rect 243726 416898 243768 417134
rect 243448 416866 243768 416898
rect 253688 417454 254008 417486
rect 253688 417218 253730 417454
rect 253966 417218 254008 417454
rect 253688 417134 254008 417218
rect 253688 416898 253730 417134
rect 253966 416898 254008 417134
rect 253688 416866 254008 416898
rect 263928 417454 264248 417486
rect 263928 417218 263970 417454
rect 264206 417218 264248 417454
rect 263928 417134 264248 417218
rect 263928 416898 263970 417134
rect 264206 416898 264248 417134
rect 263928 416866 264248 416898
rect 274168 417454 274488 417486
rect 274168 417218 274210 417454
rect 274446 417218 274488 417454
rect 274168 417134 274488 417218
rect 274168 416898 274210 417134
rect 274446 416898 274488 417134
rect 274168 416866 274488 416898
rect 284408 417454 284728 417486
rect 284408 417218 284450 417454
rect 284686 417218 284728 417454
rect 284408 417134 284728 417218
rect 284408 416898 284450 417134
rect 284686 416898 284728 417134
rect 284408 416866 284728 416898
rect 294648 417454 294968 417486
rect 294648 417218 294690 417454
rect 294926 417218 294968 417454
rect 294648 417134 294968 417218
rect 294648 416898 294690 417134
rect 294926 416898 294968 417134
rect 294648 416866 294968 416898
rect 304888 417454 305208 417486
rect 304888 417218 304930 417454
rect 305166 417218 305208 417454
rect 304888 417134 305208 417218
rect 304888 416898 304930 417134
rect 305166 416898 305208 417134
rect 304888 416866 305208 416898
rect 315128 417454 315448 417486
rect 315128 417218 315170 417454
rect 315406 417218 315448 417454
rect 315128 417134 315448 417218
rect 315128 416898 315170 417134
rect 315406 416898 315448 417134
rect 315128 416866 315448 416898
rect 325368 417454 325688 417486
rect 325368 417218 325410 417454
rect 325646 417218 325688 417454
rect 325368 417134 325688 417218
rect 325368 416898 325410 417134
rect 325646 416898 325688 417134
rect 325368 416866 325688 416898
rect 335608 417454 335928 417486
rect 335608 417218 335650 417454
rect 335886 417218 335928 417454
rect 335608 417134 335928 417218
rect 335608 416898 335650 417134
rect 335886 416898 335928 417134
rect 335608 416866 335928 416898
rect 345848 417454 346168 417486
rect 345848 417218 345890 417454
rect 346126 417218 346168 417454
rect 345848 417134 346168 417218
rect 345848 416898 345890 417134
rect 346126 416898 346168 417134
rect 345848 416866 346168 416898
rect 356088 417454 356408 417486
rect 356088 417218 356130 417454
rect 356366 417218 356408 417454
rect 356088 417134 356408 417218
rect 356088 416898 356130 417134
rect 356366 416898 356408 417134
rect 356088 416866 356408 416898
rect 366328 417454 366648 417486
rect 366328 417218 366370 417454
rect 366606 417218 366648 417454
rect 366328 417134 366648 417218
rect 366328 416898 366370 417134
rect 366606 416898 366648 417134
rect 366328 416866 366648 416898
rect 376568 417454 376888 417486
rect 376568 417218 376610 417454
rect 376846 417218 376888 417454
rect 376568 417134 376888 417218
rect 376568 416898 376610 417134
rect 376846 416898 376888 417134
rect 376568 416866 376888 416898
rect 386808 417454 387128 417486
rect 386808 417218 386850 417454
rect 387086 417218 387128 417454
rect 386808 417134 387128 417218
rect 386808 416898 386850 417134
rect 387086 416898 387128 417134
rect 386808 416866 387128 416898
rect 397048 417454 397368 417486
rect 397048 417218 397090 417454
rect 397326 417218 397368 417454
rect 397048 417134 397368 417218
rect 397048 416898 397090 417134
rect 397326 416898 397368 417134
rect 397048 416866 397368 416898
rect 407288 417454 407608 417486
rect 407288 417218 407330 417454
rect 407566 417218 407608 417454
rect 407288 417134 407608 417218
rect 407288 416898 407330 417134
rect 407566 416898 407608 417134
rect 407288 416866 407608 416898
rect 417528 417454 417848 417486
rect 417528 417218 417570 417454
rect 417806 417218 417848 417454
rect 417528 417134 417848 417218
rect 417528 416898 417570 417134
rect 417806 416898 417848 417134
rect 417528 416866 417848 416898
rect 427768 417454 428088 417486
rect 427768 417218 427810 417454
rect 428046 417218 428088 417454
rect 427768 417134 428088 417218
rect 427768 416898 427810 417134
rect 428046 416898 428088 417134
rect 427768 416866 428088 416898
rect 438008 417454 438328 417486
rect 438008 417218 438050 417454
rect 438286 417218 438328 417454
rect 438008 417134 438328 417218
rect 438008 416898 438050 417134
rect 438286 416898 438328 417134
rect 438008 416866 438328 416898
rect 448248 417454 448568 417486
rect 448248 417218 448290 417454
rect 448526 417218 448568 417454
rect 448248 417134 448568 417218
rect 448248 416898 448290 417134
rect 448526 416898 448568 417134
rect 448248 416866 448568 416898
rect 458488 417454 458808 417486
rect 458488 417218 458530 417454
rect 458766 417218 458808 417454
rect 458488 417134 458808 417218
rect 458488 416898 458530 417134
rect 458766 416898 458808 417134
rect 458488 416866 458808 416898
rect 468728 417454 469048 417486
rect 468728 417218 468770 417454
rect 469006 417218 469048 417454
rect 468728 417134 469048 417218
rect 468728 416898 468770 417134
rect 469006 416898 469048 417134
rect 468728 416866 469048 416898
rect 478968 417454 479288 417486
rect 478968 417218 479010 417454
rect 479246 417218 479288 417454
rect 478968 417134 479288 417218
rect 478968 416898 479010 417134
rect 479246 416898 479288 417134
rect 478968 416866 479288 416898
rect 489208 417454 489528 417486
rect 489208 417218 489250 417454
rect 489486 417218 489528 417454
rect 489208 417134 489528 417218
rect 489208 416898 489250 417134
rect 489486 416898 489528 417134
rect 489208 416866 489528 416898
rect 499448 417454 499768 417486
rect 499448 417218 499490 417454
rect 499726 417218 499768 417454
rect 499448 417134 499768 417218
rect 499448 416898 499490 417134
rect 499726 416898 499768 417134
rect 499448 416866 499768 416898
rect 509688 417454 510008 417486
rect 509688 417218 509730 417454
rect 509966 417218 510008 417454
rect 509688 417134 510008 417218
rect 509688 416898 509730 417134
rect 509966 416898 510008 417134
rect 509688 416866 510008 416898
rect 519928 417454 520248 417486
rect 519928 417218 519970 417454
rect 520206 417218 520248 417454
rect 519928 417134 520248 417218
rect 519928 416898 519970 417134
rect 520206 416898 520248 417134
rect 519928 416866 520248 416898
rect 530168 417454 530488 417486
rect 530168 417218 530210 417454
rect 530446 417218 530488 417454
rect 530168 417134 530488 417218
rect 530168 416898 530210 417134
rect 530446 416898 530488 417134
rect 530168 416866 530488 416898
rect 15754 402938 15786 403174
rect 16022 402938 16106 403174
rect 16342 402938 16374 403174
rect 15754 402854 16374 402938
rect 15754 402618 15786 402854
rect 16022 402618 16106 402854
rect 16342 402618 16374 402854
rect 15754 367174 16374 402618
rect 541714 406894 542334 442338
rect 541714 406658 541746 406894
rect 541982 406658 542066 406894
rect 542302 406658 542334 406894
rect 541714 406574 542334 406658
rect 541714 406338 541746 406574
rect 541982 406338 542066 406574
rect 542302 406338 542334 406574
rect 23288 399454 23608 399486
rect 23288 399218 23330 399454
rect 23566 399218 23608 399454
rect 23288 399134 23608 399218
rect 23288 398898 23330 399134
rect 23566 398898 23608 399134
rect 23288 398866 23608 398898
rect 33528 399454 33848 399486
rect 33528 399218 33570 399454
rect 33806 399218 33848 399454
rect 33528 399134 33848 399218
rect 33528 398898 33570 399134
rect 33806 398898 33848 399134
rect 33528 398866 33848 398898
rect 43768 399454 44088 399486
rect 43768 399218 43810 399454
rect 44046 399218 44088 399454
rect 43768 399134 44088 399218
rect 43768 398898 43810 399134
rect 44046 398898 44088 399134
rect 43768 398866 44088 398898
rect 54008 399454 54328 399486
rect 54008 399218 54050 399454
rect 54286 399218 54328 399454
rect 54008 399134 54328 399218
rect 54008 398898 54050 399134
rect 54286 398898 54328 399134
rect 54008 398866 54328 398898
rect 64248 399454 64568 399486
rect 64248 399218 64290 399454
rect 64526 399218 64568 399454
rect 64248 399134 64568 399218
rect 64248 398898 64290 399134
rect 64526 398898 64568 399134
rect 64248 398866 64568 398898
rect 74488 399454 74808 399486
rect 74488 399218 74530 399454
rect 74766 399218 74808 399454
rect 74488 399134 74808 399218
rect 74488 398898 74530 399134
rect 74766 398898 74808 399134
rect 74488 398866 74808 398898
rect 84728 399454 85048 399486
rect 84728 399218 84770 399454
rect 85006 399218 85048 399454
rect 84728 399134 85048 399218
rect 84728 398898 84770 399134
rect 85006 398898 85048 399134
rect 84728 398866 85048 398898
rect 94968 399454 95288 399486
rect 94968 399218 95010 399454
rect 95246 399218 95288 399454
rect 94968 399134 95288 399218
rect 94968 398898 95010 399134
rect 95246 398898 95288 399134
rect 94968 398866 95288 398898
rect 105208 399454 105528 399486
rect 105208 399218 105250 399454
rect 105486 399218 105528 399454
rect 105208 399134 105528 399218
rect 105208 398898 105250 399134
rect 105486 398898 105528 399134
rect 105208 398866 105528 398898
rect 115448 399454 115768 399486
rect 115448 399218 115490 399454
rect 115726 399218 115768 399454
rect 115448 399134 115768 399218
rect 115448 398898 115490 399134
rect 115726 398898 115768 399134
rect 115448 398866 115768 398898
rect 125688 399454 126008 399486
rect 125688 399218 125730 399454
rect 125966 399218 126008 399454
rect 125688 399134 126008 399218
rect 125688 398898 125730 399134
rect 125966 398898 126008 399134
rect 125688 398866 126008 398898
rect 135928 399454 136248 399486
rect 135928 399218 135970 399454
rect 136206 399218 136248 399454
rect 135928 399134 136248 399218
rect 135928 398898 135970 399134
rect 136206 398898 136248 399134
rect 135928 398866 136248 398898
rect 146168 399454 146488 399486
rect 146168 399218 146210 399454
rect 146446 399218 146488 399454
rect 146168 399134 146488 399218
rect 146168 398898 146210 399134
rect 146446 398898 146488 399134
rect 146168 398866 146488 398898
rect 156408 399454 156728 399486
rect 156408 399218 156450 399454
rect 156686 399218 156728 399454
rect 156408 399134 156728 399218
rect 156408 398898 156450 399134
rect 156686 398898 156728 399134
rect 156408 398866 156728 398898
rect 166648 399454 166968 399486
rect 166648 399218 166690 399454
rect 166926 399218 166968 399454
rect 166648 399134 166968 399218
rect 166648 398898 166690 399134
rect 166926 398898 166968 399134
rect 166648 398866 166968 398898
rect 176888 399454 177208 399486
rect 176888 399218 176930 399454
rect 177166 399218 177208 399454
rect 176888 399134 177208 399218
rect 176888 398898 176930 399134
rect 177166 398898 177208 399134
rect 176888 398866 177208 398898
rect 187128 399454 187448 399486
rect 187128 399218 187170 399454
rect 187406 399218 187448 399454
rect 187128 399134 187448 399218
rect 187128 398898 187170 399134
rect 187406 398898 187448 399134
rect 187128 398866 187448 398898
rect 197368 399454 197688 399486
rect 197368 399218 197410 399454
rect 197646 399218 197688 399454
rect 197368 399134 197688 399218
rect 197368 398898 197410 399134
rect 197646 398898 197688 399134
rect 197368 398866 197688 398898
rect 207608 399454 207928 399486
rect 207608 399218 207650 399454
rect 207886 399218 207928 399454
rect 207608 399134 207928 399218
rect 207608 398898 207650 399134
rect 207886 398898 207928 399134
rect 207608 398866 207928 398898
rect 217848 399454 218168 399486
rect 217848 399218 217890 399454
rect 218126 399218 218168 399454
rect 217848 399134 218168 399218
rect 217848 398898 217890 399134
rect 218126 398898 218168 399134
rect 217848 398866 218168 398898
rect 228088 399454 228408 399486
rect 228088 399218 228130 399454
rect 228366 399218 228408 399454
rect 228088 399134 228408 399218
rect 228088 398898 228130 399134
rect 228366 398898 228408 399134
rect 228088 398866 228408 398898
rect 238328 399454 238648 399486
rect 238328 399218 238370 399454
rect 238606 399218 238648 399454
rect 238328 399134 238648 399218
rect 238328 398898 238370 399134
rect 238606 398898 238648 399134
rect 238328 398866 238648 398898
rect 248568 399454 248888 399486
rect 248568 399218 248610 399454
rect 248846 399218 248888 399454
rect 248568 399134 248888 399218
rect 248568 398898 248610 399134
rect 248846 398898 248888 399134
rect 248568 398866 248888 398898
rect 258808 399454 259128 399486
rect 258808 399218 258850 399454
rect 259086 399218 259128 399454
rect 258808 399134 259128 399218
rect 258808 398898 258850 399134
rect 259086 398898 259128 399134
rect 258808 398866 259128 398898
rect 269048 399454 269368 399486
rect 269048 399218 269090 399454
rect 269326 399218 269368 399454
rect 269048 399134 269368 399218
rect 269048 398898 269090 399134
rect 269326 398898 269368 399134
rect 269048 398866 269368 398898
rect 279288 399454 279608 399486
rect 279288 399218 279330 399454
rect 279566 399218 279608 399454
rect 279288 399134 279608 399218
rect 279288 398898 279330 399134
rect 279566 398898 279608 399134
rect 279288 398866 279608 398898
rect 289528 399454 289848 399486
rect 289528 399218 289570 399454
rect 289806 399218 289848 399454
rect 289528 399134 289848 399218
rect 289528 398898 289570 399134
rect 289806 398898 289848 399134
rect 289528 398866 289848 398898
rect 299768 399454 300088 399486
rect 299768 399218 299810 399454
rect 300046 399218 300088 399454
rect 299768 399134 300088 399218
rect 299768 398898 299810 399134
rect 300046 398898 300088 399134
rect 299768 398866 300088 398898
rect 310008 399454 310328 399486
rect 310008 399218 310050 399454
rect 310286 399218 310328 399454
rect 310008 399134 310328 399218
rect 310008 398898 310050 399134
rect 310286 398898 310328 399134
rect 310008 398866 310328 398898
rect 320248 399454 320568 399486
rect 320248 399218 320290 399454
rect 320526 399218 320568 399454
rect 320248 399134 320568 399218
rect 320248 398898 320290 399134
rect 320526 398898 320568 399134
rect 320248 398866 320568 398898
rect 330488 399454 330808 399486
rect 330488 399218 330530 399454
rect 330766 399218 330808 399454
rect 330488 399134 330808 399218
rect 330488 398898 330530 399134
rect 330766 398898 330808 399134
rect 330488 398866 330808 398898
rect 340728 399454 341048 399486
rect 340728 399218 340770 399454
rect 341006 399218 341048 399454
rect 340728 399134 341048 399218
rect 340728 398898 340770 399134
rect 341006 398898 341048 399134
rect 340728 398866 341048 398898
rect 350968 399454 351288 399486
rect 350968 399218 351010 399454
rect 351246 399218 351288 399454
rect 350968 399134 351288 399218
rect 350968 398898 351010 399134
rect 351246 398898 351288 399134
rect 350968 398866 351288 398898
rect 361208 399454 361528 399486
rect 361208 399218 361250 399454
rect 361486 399218 361528 399454
rect 361208 399134 361528 399218
rect 361208 398898 361250 399134
rect 361486 398898 361528 399134
rect 361208 398866 361528 398898
rect 371448 399454 371768 399486
rect 371448 399218 371490 399454
rect 371726 399218 371768 399454
rect 371448 399134 371768 399218
rect 371448 398898 371490 399134
rect 371726 398898 371768 399134
rect 371448 398866 371768 398898
rect 381688 399454 382008 399486
rect 381688 399218 381730 399454
rect 381966 399218 382008 399454
rect 381688 399134 382008 399218
rect 381688 398898 381730 399134
rect 381966 398898 382008 399134
rect 381688 398866 382008 398898
rect 391928 399454 392248 399486
rect 391928 399218 391970 399454
rect 392206 399218 392248 399454
rect 391928 399134 392248 399218
rect 391928 398898 391970 399134
rect 392206 398898 392248 399134
rect 391928 398866 392248 398898
rect 402168 399454 402488 399486
rect 402168 399218 402210 399454
rect 402446 399218 402488 399454
rect 402168 399134 402488 399218
rect 402168 398898 402210 399134
rect 402446 398898 402488 399134
rect 402168 398866 402488 398898
rect 412408 399454 412728 399486
rect 412408 399218 412450 399454
rect 412686 399218 412728 399454
rect 412408 399134 412728 399218
rect 412408 398898 412450 399134
rect 412686 398898 412728 399134
rect 412408 398866 412728 398898
rect 422648 399454 422968 399486
rect 422648 399218 422690 399454
rect 422926 399218 422968 399454
rect 422648 399134 422968 399218
rect 422648 398898 422690 399134
rect 422926 398898 422968 399134
rect 422648 398866 422968 398898
rect 432888 399454 433208 399486
rect 432888 399218 432930 399454
rect 433166 399218 433208 399454
rect 432888 399134 433208 399218
rect 432888 398898 432930 399134
rect 433166 398898 433208 399134
rect 432888 398866 433208 398898
rect 443128 399454 443448 399486
rect 443128 399218 443170 399454
rect 443406 399218 443448 399454
rect 443128 399134 443448 399218
rect 443128 398898 443170 399134
rect 443406 398898 443448 399134
rect 443128 398866 443448 398898
rect 453368 399454 453688 399486
rect 453368 399218 453410 399454
rect 453646 399218 453688 399454
rect 453368 399134 453688 399218
rect 453368 398898 453410 399134
rect 453646 398898 453688 399134
rect 453368 398866 453688 398898
rect 463608 399454 463928 399486
rect 463608 399218 463650 399454
rect 463886 399218 463928 399454
rect 463608 399134 463928 399218
rect 463608 398898 463650 399134
rect 463886 398898 463928 399134
rect 463608 398866 463928 398898
rect 473848 399454 474168 399486
rect 473848 399218 473890 399454
rect 474126 399218 474168 399454
rect 473848 399134 474168 399218
rect 473848 398898 473890 399134
rect 474126 398898 474168 399134
rect 473848 398866 474168 398898
rect 484088 399454 484408 399486
rect 484088 399218 484130 399454
rect 484366 399218 484408 399454
rect 484088 399134 484408 399218
rect 484088 398898 484130 399134
rect 484366 398898 484408 399134
rect 484088 398866 484408 398898
rect 494328 399454 494648 399486
rect 494328 399218 494370 399454
rect 494606 399218 494648 399454
rect 494328 399134 494648 399218
rect 494328 398898 494370 399134
rect 494606 398898 494648 399134
rect 494328 398866 494648 398898
rect 504568 399454 504888 399486
rect 504568 399218 504610 399454
rect 504846 399218 504888 399454
rect 504568 399134 504888 399218
rect 504568 398898 504610 399134
rect 504846 398898 504888 399134
rect 504568 398866 504888 398898
rect 514808 399454 515128 399486
rect 514808 399218 514850 399454
rect 515086 399218 515128 399454
rect 514808 399134 515128 399218
rect 514808 398898 514850 399134
rect 515086 398898 515128 399134
rect 514808 398866 515128 398898
rect 525048 399454 525368 399486
rect 525048 399218 525090 399454
rect 525326 399218 525368 399454
rect 525048 399134 525368 399218
rect 525048 398898 525090 399134
rect 525326 398898 525368 399134
rect 525048 398866 525368 398898
rect 535288 399454 535608 399486
rect 535288 399218 535330 399454
rect 535566 399218 535608 399454
rect 535288 399134 535608 399218
rect 535288 398898 535330 399134
rect 535566 398898 535608 399134
rect 535288 398866 535608 398898
rect 28408 381454 28728 381486
rect 28408 381218 28450 381454
rect 28686 381218 28728 381454
rect 28408 381134 28728 381218
rect 28408 380898 28450 381134
rect 28686 380898 28728 381134
rect 28408 380866 28728 380898
rect 38648 381454 38968 381486
rect 38648 381218 38690 381454
rect 38926 381218 38968 381454
rect 38648 381134 38968 381218
rect 38648 380898 38690 381134
rect 38926 380898 38968 381134
rect 38648 380866 38968 380898
rect 48888 381454 49208 381486
rect 48888 381218 48930 381454
rect 49166 381218 49208 381454
rect 48888 381134 49208 381218
rect 48888 380898 48930 381134
rect 49166 380898 49208 381134
rect 48888 380866 49208 380898
rect 59128 381454 59448 381486
rect 59128 381218 59170 381454
rect 59406 381218 59448 381454
rect 59128 381134 59448 381218
rect 59128 380898 59170 381134
rect 59406 380898 59448 381134
rect 59128 380866 59448 380898
rect 69368 381454 69688 381486
rect 69368 381218 69410 381454
rect 69646 381218 69688 381454
rect 69368 381134 69688 381218
rect 69368 380898 69410 381134
rect 69646 380898 69688 381134
rect 69368 380866 69688 380898
rect 79608 381454 79928 381486
rect 79608 381218 79650 381454
rect 79886 381218 79928 381454
rect 79608 381134 79928 381218
rect 79608 380898 79650 381134
rect 79886 380898 79928 381134
rect 79608 380866 79928 380898
rect 89848 381454 90168 381486
rect 89848 381218 89890 381454
rect 90126 381218 90168 381454
rect 89848 381134 90168 381218
rect 89848 380898 89890 381134
rect 90126 380898 90168 381134
rect 89848 380866 90168 380898
rect 100088 381454 100408 381486
rect 100088 381218 100130 381454
rect 100366 381218 100408 381454
rect 100088 381134 100408 381218
rect 100088 380898 100130 381134
rect 100366 380898 100408 381134
rect 100088 380866 100408 380898
rect 110328 381454 110648 381486
rect 110328 381218 110370 381454
rect 110606 381218 110648 381454
rect 110328 381134 110648 381218
rect 110328 380898 110370 381134
rect 110606 380898 110648 381134
rect 110328 380866 110648 380898
rect 120568 381454 120888 381486
rect 120568 381218 120610 381454
rect 120846 381218 120888 381454
rect 120568 381134 120888 381218
rect 120568 380898 120610 381134
rect 120846 380898 120888 381134
rect 120568 380866 120888 380898
rect 130808 381454 131128 381486
rect 130808 381218 130850 381454
rect 131086 381218 131128 381454
rect 130808 381134 131128 381218
rect 130808 380898 130850 381134
rect 131086 380898 131128 381134
rect 130808 380866 131128 380898
rect 141048 381454 141368 381486
rect 141048 381218 141090 381454
rect 141326 381218 141368 381454
rect 141048 381134 141368 381218
rect 141048 380898 141090 381134
rect 141326 380898 141368 381134
rect 141048 380866 141368 380898
rect 151288 381454 151608 381486
rect 151288 381218 151330 381454
rect 151566 381218 151608 381454
rect 151288 381134 151608 381218
rect 151288 380898 151330 381134
rect 151566 380898 151608 381134
rect 151288 380866 151608 380898
rect 161528 381454 161848 381486
rect 161528 381218 161570 381454
rect 161806 381218 161848 381454
rect 161528 381134 161848 381218
rect 161528 380898 161570 381134
rect 161806 380898 161848 381134
rect 161528 380866 161848 380898
rect 171768 381454 172088 381486
rect 171768 381218 171810 381454
rect 172046 381218 172088 381454
rect 171768 381134 172088 381218
rect 171768 380898 171810 381134
rect 172046 380898 172088 381134
rect 171768 380866 172088 380898
rect 182008 381454 182328 381486
rect 182008 381218 182050 381454
rect 182286 381218 182328 381454
rect 182008 381134 182328 381218
rect 182008 380898 182050 381134
rect 182286 380898 182328 381134
rect 182008 380866 182328 380898
rect 192248 381454 192568 381486
rect 192248 381218 192290 381454
rect 192526 381218 192568 381454
rect 192248 381134 192568 381218
rect 192248 380898 192290 381134
rect 192526 380898 192568 381134
rect 192248 380866 192568 380898
rect 202488 381454 202808 381486
rect 202488 381218 202530 381454
rect 202766 381218 202808 381454
rect 202488 381134 202808 381218
rect 202488 380898 202530 381134
rect 202766 380898 202808 381134
rect 202488 380866 202808 380898
rect 212728 381454 213048 381486
rect 212728 381218 212770 381454
rect 213006 381218 213048 381454
rect 212728 381134 213048 381218
rect 212728 380898 212770 381134
rect 213006 380898 213048 381134
rect 212728 380866 213048 380898
rect 222968 381454 223288 381486
rect 222968 381218 223010 381454
rect 223246 381218 223288 381454
rect 222968 381134 223288 381218
rect 222968 380898 223010 381134
rect 223246 380898 223288 381134
rect 222968 380866 223288 380898
rect 233208 381454 233528 381486
rect 233208 381218 233250 381454
rect 233486 381218 233528 381454
rect 233208 381134 233528 381218
rect 233208 380898 233250 381134
rect 233486 380898 233528 381134
rect 233208 380866 233528 380898
rect 243448 381454 243768 381486
rect 243448 381218 243490 381454
rect 243726 381218 243768 381454
rect 243448 381134 243768 381218
rect 243448 380898 243490 381134
rect 243726 380898 243768 381134
rect 243448 380866 243768 380898
rect 253688 381454 254008 381486
rect 253688 381218 253730 381454
rect 253966 381218 254008 381454
rect 253688 381134 254008 381218
rect 253688 380898 253730 381134
rect 253966 380898 254008 381134
rect 253688 380866 254008 380898
rect 263928 381454 264248 381486
rect 263928 381218 263970 381454
rect 264206 381218 264248 381454
rect 263928 381134 264248 381218
rect 263928 380898 263970 381134
rect 264206 380898 264248 381134
rect 263928 380866 264248 380898
rect 274168 381454 274488 381486
rect 274168 381218 274210 381454
rect 274446 381218 274488 381454
rect 274168 381134 274488 381218
rect 274168 380898 274210 381134
rect 274446 380898 274488 381134
rect 274168 380866 274488 380898
rect 284408 381454 284728 381486
rect 284408 381218 284450 381454
rect 284686 381218 284728 381454
rect 284408 381134 284728 381218
rect 284408 380898 284450 381134
rect 284686 380898 284728 381134
rect 284408 380866 284728 380898
rect 294648 381454 294968 381486
rect 294648 381218 294690 381454
rect 294926 381218 294968 381454
rect 294648 381134 294968 381218
rect 294648 380898 294690 381134
rect 294926 380898 294968 381134
rect 294648 380866 294968 380898
rect 304888 381454 305208 381486
rect 304888 381218 304930 381454
rect 305166 381218 305208 381454
rect 304888 381134 305208 381218
rect 304888 380898 304930 381134
rect 305166 380898 305208 381134
rect 304888 380866 305208 380898
rect 315128 381454 315448 381486
rect 315128 381218 315170 381454
rect 315406 381218 315448 381454
rect 315128 381134 315448 381218
rect 315128 380898 315170 381134
rect 315406 380898 315448 381134
rect 315128 380866 315448 380898
rect 325368 381454 325688 381486
rect 325368 381218 325410 381454
rect 325646 381218 325688 381454
rect 325368 381134 325688 381218
rect 325368 380898 325410 381134
rect 325646 380898 325688 381134
rect 325368 380866 325688 380898
rect 335608 381454 335928 381486
rect 335608 381218 335650 381454
rect 335886 381218 335928 381454
rect 335608 381134 335928 381218
rect 335608 380898 335650 381134
rect 335886 380898 335928 381134
rect 335608 380866 335928 380898
rect 345848 381454 346168 381486
rect 345848 381218 345890 381454
rect 346126 381218 346168 381454
rect 345848 381134 346168 381218
rect 345848 380898 345890 381134
rect 346126 380898 346168 381134
rect 345848 380866 346168 380898
rect 356088 381454 356408 381486
rect 356088 381218 356130 381454
rect 356366 381218 356408 381454
rect 356088 381134 356408 381218
rect 356088 380898 356130 381134
rect 356366 380898 356408 381134
rect 356088 380866 356408 380898
rect 366328 381454 366648 381486
rect 366328 381218 366370 381454
rect 366606 381218 366648 381454
rect 366328 381134 366648 381218
rect 366328 380898 366370 381134
rect 366606 380898 366648 381134
rect 366328 380866 366648 380898
rect 376568 381454 376888 381486
rect 376568 381218 376610 381454
rect 376846 381218 376888 381454
rect 376568 381134 376888 381218
rect 376568 380898 376610 381134
rect 376846 380898 376888 381134
rect 376568 380866 376888 380898
rect 386808 381454 387128 381486
rect 386808 381218 386850 381454
rect 387086 381218 387128 381454
rect 386808 381134 387128 381218
rect 386808 380898 386850 381134
rect 387086 380898 387128 381134
rect 386808 380866 387128 380898
rect 397048 381454 397368 381486
rect 397048 381218 397090 381454
rect 397326 381218 397368 381454
rect 397048 381134 397368 381218
rect 397048 380898 397090 381134
rect 397326 380898 397368 381134
rect 397048 380866 397368 380898
rect 407288 381454 407608 381486
rect 407288 381218 407330 381454
rect 407566 381218 407608 381454
rect 407288 381134 407608 381218
rect 407288 380898 407330 381134
rect 407566 380898 407608 381134
rect 407288 380866 407608 380898
rect 417528 381454 417848 381486
rect 417528 381218 417570 381454
rect 417806 381218 417848 381454
rect 417528 381134 417848 381218
rect 417528 380898 417570 381134
rect 417806 380898 417848 381134
rect 417528 380866 417848 380898
rect 427768 381454 428088 381486
rect 427768 381218 427810 381454
rect 428046 381218 428088 381454
rect 427768 381134 428088 381218
rect 427768 380898 427810 381134
rect 428046 380898 428088 381134
rect 427768 380866 428088 380898
rect 438008 381454 438328 381486
rect 438008 381218 438050 381454
rect 438286 381218 438328 381454
rect 438008 381134 438328 381218
rect 438008 380898 438050 381134
rect 438286 380898 438328 381134
rect 438008 380866 438328 380898
rect 448248 381454 448568 381486
rect 448248 381218 448290 381454
rect 448526 381218 448568 381454
rect 448248 381134 448568 381218
rect 448248 380898 448290 381134
rect 448526 380898 448568 381134
rect 448248 380866 448568 380898
rect 458488 381454 458808 381486
rect 458488 381218 458530 381454
rect 458766 381218 458808 381454
rect 458488 381134 458808 381218
rect 458488 380898 458530 381134
rect 458766 380898 458808 381134
rect 458488 380866 458808 380898
rect 468728 381454 469048 381486
rect 468728 381218 468770 381454
rect 469006 381218 469048 381454
rect 468728 381134 469048 381218
rect 468728 380898 468770 381134
rect 469006 380898 469048 381134
rect 468728 380866 469048 380898
rect 478968 381454 479288 381486
rect 478968 381218 479010 381454
rect 479246 381218 479288 381454
rect 478968 381134 479288 381218
rect 478968 380898 479010 381134
rect 479246 380898 479288 381134
rect 478968 380866 479288 380898
rect 489208 381454 489528 381486
rect 489208 381218 489250 381454
rect 489486 381218 489528 381454
rect 489208 381134 489528 381218
rect 489208 380898 489250 381134
rect 489486 380898 489528 381134
rect 489208 380866 489528 380898
rect 499448 381454 499768 381486
rect 499448 381218 499490 381454
rect 499726 381218 499768 381454
rect 499448 381134 499768 381218
rect 499448 380898 499490 381134
rect 499726 380898 499768 381134
rect 499448 380866 499768 380898
rect 509688 381454 510008 381486
rect 509688 381218 509730 381454
rect 509966 381218 510008 381454
rect 509688 381134 510008 381218
rect 509688 380898 509730 381134
rect 509966 380898 510008 381134
rect 509688 380866 510008 380898
rect 519928 381454 520248 381486
rect 519928 381218 519970 381454
rect 520206 381218 520248 381454
rect 519928 381134 520248 381218
rect 519928 380898 519970 381134
rect 520206 380898 520248 381134
rect 519928 380866 520248 380898
rect 530168 381454 530488 381486
rect 530168 381218 530210 381454
rect 530446 381218 530488 381454
rect 530168 381134 530488 381218
rect 530168 380898 530210 381134
rect 530446 380898 530488 381134
rect 530168 380866 530488 380898
rect 15754 366938 15786 367174
rect 16022 366938 16106 367174
rect 16342 366938 16374 367174
rect 15754 366854 16374 366938
rect 15754 366618 15786 366854
rect 16022 366618 16106 366854
rect 16342 366618 16374 366854
rect 15754 331174 16374 366618
rect 541714 370894 542334 406338
rect 541714 370658 541746 370894
rect 541982 370658 542066 370894
rect 542302 370658 542334 370894
rect 541714 370574 542334 370658
rect 541714 370338 541746 370574
rect 541982 370338 542066 370574
rect 542302 370338 542334 370574
rect 23288 363454 23608 363486
rect 23288 363218 23330 363454
rect 23566 363218 23608 363454
rect 23288 363134 23608 363218
rect 23288 362898 23330 363134
rect 23566 362898 23608 363134
rect 23288 362866 23608 362898
rect 33528 363454 33848 363486
rect 33528 363218 33570 363454
rect 33806 363218 33848 363454
rect 33528 363134 33848 363218
rect 33528 362898 33570 363134
rect 33806 362898 33848 363134
rect 33528 362866 33848 362898
rect 43768 363454 44088 363486
rect 43768 363218 43810 363454
rect 44046 363218 44088 363454
rect 43768 363134 44088 363218
rect 43768 362898 43810 363134
rect 44046 362898 44088 363134
rect 43768 362866 44088 362898
rect 54008 363454 54328 363486
rect 54008 363218 54050 363454
rect 54286 363218 54328 363454
rect 54008 363134 54328 363218
rect 54008 362898 54050 363134
rect 54286 362898 54328 363134
rect 54008 362866 54328 362898
rect 64248 363454 64568 363486
rect 64248 363218 64290 363454
rect 64526 363218 64568 363454
rect 64248 363134 64568 363218
rect 64248 362898 64290 363134
rect 64526 362898 64568 363134
rect 64248 362866 64568 362898
rect 74488 363454 74808 363486
rect 74488 363218 74530 363454
rect 74766 363218 74808 363454
rect 74488 363134 74808 363218
rect 74488 362898 74530 363134
rect 74766 362898 74808 363134
rect 74488 362866 74808 362898
rect 84728 363454 85048 363486
rect 84728 363218 84770 363454
rect 85006 363218 85048 363454
rect 84728 363134 85048 363218
rect 84728 362898 84770 363134
rect 85006 362898 85048 363134
rect 84728 362866 85048 362898
rect 94968 363454 95288 363486
rect 94968 363218 95010 363454
rect 95246 363218 95288 363454
rect 94968 363134 95288 363218
rect 94968 362898 95010 363134
rect 95246 362898 95288 363134
rect 94968 362866 95288 362898
rect 105208 363454 105528 363486
rect 105208 363218 105250 363454
rect 105486 363218 105528 363454
rect 105208 363134 105528 363218
rect 105208 362898 105250 363134
rect 105486 362898 105528 363134
rect 105208 362866 105528 362898
rect 115448 363454 115768 363486
rect 115448 363218 115490 363454
rect 115726 363218 115768 363454
rect 115448 363134 115768 363218
rect 115448 362898 115490 363134
rect 115726 362898 115768 363134
rect 115448 362866 115768 362898
rect 125688 363454 126008 363486
rect 125688 363218 125730 363454
rect 125966 363218 126008 363454
rect 125688 363134 126008 363218
rect 125688 362898 125730 363134
rect 125966 362898 126008 363134
rect 125688 362866 126008 362898
rect 135928 363454 136248 363486
rect 135928 363218 135970 363454
rect 136206 363218 136248 363454
rect 135928 363134 136248 363218
rect 135928 362898 135970 363134
rect 136206 362898 136248 363134
rect 135928 362866 136248 362898
rect 146168 363454 146488 363486
rect 146168 363218 146210 363454
rect 146446 363218 146488 363454
rect 146168 363134 146488 363218
rect 146168 362898 146210 363134
rect 146446 362898 146488 363134
rect 146168 362866 146488 362898
rect 156408 363454 156728 363486
rect 156408 363218 156450 363454
rect 156686 363218 156728 363454
rect 156408 363134 156728 363218
rect 156408 362898 156450 363134
rect 156686 362898 156728 363134
rect 156408 362866 156728 362898
rect 166648 363454 166968 363486
rect 166648 363218 166690 363454
rect 166926 363218 166968 363454
rect 166648 363134 166968 363218
rect 166648 362898 166690 363134
rect 166926 362898 166968 363134
rect 166648 362866 166968 362898
rect 176888 363454 177208 363486
rect 176888 363218 176930 363454
rect 177166 363218 177208 363454
rect 176888 363134 177208 363218
rect 176888 362898 176930 363134
rect 177166 362898 177208 363134
rect 176888 362866 177208 362898
rect 187128 363454 187448 363486
rect 187128 363218 187170 363454
rect 187406 363218 187448 363454
rect 187128 363134 187448 363218
rect 187128 362898 187170 363134
rect 187406 362898 187448 363134
rect 187128 362866 187448 362898
rect 197368 363454 197688 363486
rect 197368 363218 197410 363454
rect 197646 363218 197688 363454
rect 197368 363134 197688 363218
rect 197368 362898 197410 363134
rect 197646 362898 197688 363134
rect 197368 362866 197688 362898
rect 207608 363454 207928 363486
rect 207608 363218 207650 363454
rect 207886 363218 207928 363454
rect 207608 363134 207928 363218
rect 207608 362898 207650 363134
rect 207886 362898 207928 363134
rect 207608 362866 207928 362898
rect 217848 363454 218168 363486
rect 217848 363218 217890 363454
rect 218126 363218 218168 363454
rect 217848 363134 218168 363218
rect 217848 362898 217890 363134
rect 218126 362898 218168 363134
rect 217848 362866 218168 362898
rect 228088 363454 228408 363486
rect 228088 363218 228130 363454
rect 228366 363218 228408 363454
rect 228088 363134 228408 363218
rect 228088 362898 228130 363134
rect 228366 362898 228408 363134
rect 228088 362866 228408 362898
rect 238328 363454 238648 363486
rect 238328 363218 238370 363454
rect 238606 363218 238648 363454
rect 238328 363134 238648 363218
rect 238328 362898 238370 363134
rect 238606 362898 238648 363134
rect 238328 362866 238648 362898
rect 248568 363454 248888 363486
rect 248568 363218 248610 363454
rect 248846 363218 248888 363454
rect 248568 363134 248888 363218
rect 248568 362898 248610 363134
rect 248846 362898 248888 363134
rect 248568 362866 248888 362898
rect 258808 363454 259128 363486
rect 258808 363218 258850 363454
rect 259086 363218 259128 363454
rect 258808 363134 259128 363218
rect 258808 362898 258850 363134
rect 259086 362898 259128 363134
rect 258808 362866 259128 362898
rect 269048 363454 269368 363486
rect 269048 363218 269090 363454
rect 269326 363218 269368 363454
rect 269048 363134 269368 363218
rect 269048 362898 269090 363134
rect 269326 362898 269368 363134
rect 269048 362866 269368 362898
rect 279288 363454 279608 363486
rect 279288 363218 279330 363454
rect 279566 363218 279608 363454
rect 279288 363134 279608 363218
rect 279288 362898 279330 363134
rect 279566 362898 279608 363134
rect 279288 362866 279608 362898
rect 289528 363454 289848 363486
rect 289528 363218 289570 363454
rect 289806 363218 289848 363454
rect 289528 363134 289848 363218
rect 289528 362898 289570 363134
rect 289806 362898 289848 363134
rect 289528 362866 289848 362898
rect 299768 363454 300088 363486
rect 299768 363218 299810 363454
rect 300046 363218 300088 363454
rect 299768 363134 300088 363218
rect 299768 362898 299810 363134
rect 300046 362898 300088 363134
rect 299768 362866 300088 362898
rect 310008 363454 310328 363486
rect 310008 363218 310050 363454
rect 310286 363218 310328 363454
rect 310008 363134 310328 363218
rect 310008 362898 310050 363134
rect 310286 362898 310328 363134
rect 310008 362866 310328 362898
rect 320248 363454 320568 363486
rect 320248 363218 320290 363454
rect 320526 363218 320568 363454
rect 320248 363134 320568 363218
rect 320248 362898 320290 363134
rect 320526 362898 320568 363134
rect 320248 362866 320568 362898
rect 330488 363454 330808 363486
rect 330488 363218 330530 363454
rect 330766 363218 330808 363454
rect 330488 363134 330808 363218
rect 330488 362898 330530 363134
rect 330766 362898 330808 363134
rect 330488 362866 330808 362898
rect 340728 363454 341048 363486
rect 340728 363218 340770 363454
rect 341006 363218 341048 363454
rect 340728 363134 341048 363218
rect 340728 362898 340770 363134
rect 341006 362898 341048 363134
rect 340728 362866 341048 362898
rect 350968 363454 351288 363486
rect 350968 363218 351010 363454
rect 351246 363218 351288 363454
rect 350968 363134 351288 363218
rect 350968 362898 351010 363134
rect 351246 362898 351288 363134
rect 350968 362866 351288 362898
rect 361208 363454 361528 363486
rect 361208 363218 361250 363454
rect 361486 363218 361528 363454
rect 361208 363134 361528 363218
rect 361208 362898 361250 363134
rect 361486 362898 361528 363134
rect 361208 362866 361528 362898
rect 371448 363454 371768 363486
rect 371448 363218 371490 363454
rect 371726 363218 371768 363454
rect 371448 363134 371768 363218
rect 371448 362898 371490 363134
rect 371726 362898 371768 363134
rect 371448 362866 371768 362898
rect 381688 363454 382008 363486
rect 381688 363218 381730 363454
rect 381966 363218 382008 363454
rect 381688 363134 382008 363218
rect 381688 362898 381730 363134
rect 381966 362898 382008 363134
rect 381688 362866 382008 362898
rect 391928 363454 392248 363486
rect 391928 363218 391970 363454
rect 392206 363218 392248 363454
rect 391928 363134 392248 363218
rect 391928 362898 391970 363134
rect 392206 362898 392248 363134
rect 391928 362866 392248 362898
rect 402168 363454 402488 363486
rect 402168 363218 402210 363454
rect 402446 363218 402488 363454
rect 402168 363134 402488 363218
rect 402168 362898 402210 363134
rect 402446 362898 402488 363134
rect 402168 362866 402488 362898
rect 412408 363454 412728 363486
rect 412408 363218 412450 363454
rect 412686 363218 412728 363454
rect 412408 363134 412728 363218
rect 412408 362898 412450 363134
rect 412686 362898 412728 363134
rect 412408 362866 412728 362898
rect 422648 363454 422968 363486
rect 422648 363218 422690 363454
rect 422926 363218 422968 363454
rect 422648 363134 422968 363218
rect 422648 362898 422690 363134
rect 422926 362898 422968 363134
rect 422648 362866 422968 362898
rect 432888 363454 433208 363486
rect 432888 363218 432930 363454
rect 433166 363218 433208 363454
rect 432888 363134 433208 363218
rect 432888 362898 432930 363134
rect 433166 362898 433208 363134
rect 432888 362866 433208 362898
rect 443128 363454 443448 363486
rect 443128 363218 443170 363454
rect 443406 363218 443448 363454
rect 443128 363134 443448 363218
rect 443128 362898 443170 363134
rect 443406 362898 443448 363134
rect 443128 362866 443448 362898
rect 453368 363454 453688 363486
rect 453368 363218 453410 363454
rect 453646 363218 453688 363454
rect 453368 363134 453688 363218
rect 453368 362898 453410 363134
rect 453646 362898 453688 363134
rect 453368 362866 453688 362898
rect 463608 363454 463928 363486
rect 463608 363218 463650 363454
rect 463886 363218 463928 363454
rect 463608 363134 463928 363218
rect 463608 362898 463650 363134
rect 463886 362898 463928 363134
rect 463608 362866 463928 362898
rect 473848 363454 474168 363486
rect 473848 363218 473890 363454
rect 474126 363218 474168 363454
rect 473848 363134 474168 363218
rect 473848 362898 473890 363134
rect 474126 362898 474168 363134
rect 473848 362866 474168 362898
rect 484088 363454 484408 363486
rect 484088 363218 484130 363454
rect 484366 363218 484408 363454
rect 484088 363134 484408 363218
rect 484088 362898 484130 363134
rect 484366 362898 484408 363134
rect 484088 362866 484408 362898
rect 494328 363454 494648 363486
rect 494328 363218 494370 363454
rect 494606 363218 494648 363454
rect 494328 363134 494648 363218
rect 494328 362898 494370 363134
rect 494606 362898 494648 363134
rect 494328 362866 494648 362898
rect 504568 363454 504888 363486
rect 504568 363218 504610 363454
rect 504846 363218 504888 363454
rect 504568 363134 504888 363218
rect 504568 362898 504610 363134
rect 504846 362898 504888 363134
rect 504568 362866 504888 362898
rect 514808 363454 515128 363486
rect 514808 363218 514850 363454
rect 515086 363218 515128 363454
rect 514808 363134 515128 363218
rect 514808 362898 514850 363134
rect 515086 362898 515128 363134
rect 514808 362866 515128 362898
rect 525048 363454 525368 363486
rect 525048 363218 525090 363454
rect 525326 363218 525368 363454
rect 525048 363134 525368 363218
rect 525048 362898 525090 363134
rect 525326 362898 525368 363134
rect 525048 362866 525368 362898
rect 535288 363454 535608 363486
rect 535288 363218 535330 363454
rect 535566 363218 535608 363454
rect 535288 363134 535608 363218
rect 535288 362898 535330 363134
rect 535566 362898 535608 363134
rect 535288 362866 535608 362898
rect 28408 345454 28728 345486
rect 28408 345218 28450 345454
rect 28686 345218 28728 345454
rect 28408 345134 28728 345218
rect 28408 344898 28450 345134
rect 28686 344898 28728 345134
rect 28408 344866 28728 344898
rect 38648 345454 38968 345486
rect 38648 345218 38690 345454
rect 38926 345218 38968 345454
rect 38648 345134 38968 345218
rect 38648 344898 38690 345134
rect 38926 344898 38968 345134
rect 38648 344866 38968 344898
rect 48888 345454 49208 345486
rect 48888 345218 48930 345454
rect 49166 345218 49208 345454
rect 48888 345134 49208 345218
rect 48888 344898 48930 345134
rect 49166 344898 49208 345134
rect 48888 344866 49208 344898
rect 59128 345454 59448 345486
rect 59128 345218 59170 345454
rect 59406 345218 59448 345454
rect 59128 345134 59448 345218
rect 59128 344898 59170 345134
rect 59406 344898 59448 345134
rect 59128 344866 59448 344898
rect 69368 345454 69688 345486
rect 69368 345218 69410 345454
rect 69646 345218 69688 345454
rect 69368 345134 69688 345218
rect 69368 344898 69410 345134
rect 69646 344898 69688 345134
rect 69368 344866 69688 344898
rect 79608 345454 79928 345486
rect 79608 345218 79650 345454
rect 79886 345218 79928 345454
rect 79608 345134 79928 345218
rect 79608 344898 79650 345134
rect 79886 344898 79928 345134
rect 79608 344866 79928 344898
rect 89848 345454 90168 345486
rect 89848 345218 89890 345454
rect 90126 345218 90168 345454
rect 89848 345134 90168 345218
rect 89848 344898 89890 345134
rect 90126 344898 90168 345134
rect 89848 344866 90168 344898
rect 100088 345454 100408 345486
rect 100088 345218 100130 345454
rect 100366 345218 100408 345454
rect 100088 345134 100408 345218
rect 100088 344898 100130 345134
rect 100366 344898 100408 345134
rect 100088 344866 100408 344898
rect 110328 345454 110648 345486
rect 110328 345218 110370 345454
rect 110606 345218 110648 345454
rect 110328 345134 110648 345218
rect 110328 344898 110370 345134
rect 110606 344898 110648 345134
rect 110328 344866 110648 344898
rect 120568 345454 120888 345486
rect 120568 345218 120610 345454
rect 120846 345218 120888 345454
rect 120568 345134 120888 345218
rect 120568 344898 120610 345134
rect 120846 344898 120888 345134
rect 120568 344866 120888 344898
rect 130808 345454 131128 345486
rect 130808 345218 130850 345454
rect 131086 345218 131128 345454
rect 130808 345134 131128 345218
rect 130808 344898 130850 345134
rect 131086 344898 131128 345134
rect 130808 344866 131128 344898
rect 141048 345454 141368 345486
rect 141048 345218 141090 345454
rect 141326 345218 141368 345454
rect 141048 345134 141368 345218
rect 141048 344898 141090 345134
rect 141326 344898 141368 345134
rect 141048 344866 141368 344898
rect 151288 345454 151608 345486
rect 151288 345218 151330 345454
rect 151566 345218 151608 345454
rect 151288 345134 151608 345218
rect 151288 344898 151330 345134
rect 151566 344898 151608 345134
rect 151288 344866 151608 344898
rect 161528 345454 161848 345486
rect 161528 345218 161570 345454
rect 161806 345218 161848 345454
rect 161528 345134 161848 345218
rect 161528 344898 161570 345134
rect 161806 344898 161848 345134
rect 161528 344866 161848 344898
rect 171768 345454 172088 345486
rect 171768 345218 171810 345454
rect 172046 345218 172088 345454
rect 171768 345134 172088 345218
rect 171768 344898 171810 345134
rect 172046 344898 172088 345134
rect 171768 344866 172088 344898
rect 182008 345454 182328 345486
rect 182008 345218 182050 345454
rect 182286 345218 182328 345454
rect 182008 345134 182328 345218
rect 182008 344898 182050 345134
rect 182286 344898 182328 345134
rect 182008 344866 182328 344898
rect 192248 345454 192568 345486
rect 192248 345218 192290 345454
rect 192526 345218 192568 345454
rect 192248 345134 192568 345218
rect 192248 344898 192290 345134
rect 192526 344898 192568 345134
rect 192248 344866 192568 344898
rect 202488 345454 202808 345486
rect 202488 345218 202530 345454
rect 202766 345218 202808 345454
rect 202488 345134 202808 345218
rect 202488 344898 202530 345134
rect 202766 344898 202808 345134
rect 202488 344866 202808 344898
rect 212728 345454 213048 345486
rect 212728 345218 212770 345454
rect 213006 345218 213048 345454
rect 212728 345134 213048 345218
rect 212728 344898 212770 345134
rect 213006 344898 213048 345134
rect 212728 344866 213048 344898
rect 222968 345454 223288 345486
rect 222968 345218 223010 345454
rect 223246 345218 223288 345454
rect 222968 345134 223288 345218
rect 222968 344898 223010 345134
rect 223246 344898 223288 345134
rect 222968 344866 223288 344898
rect 233208 345454 233528 345486
rect 233208 345218 233250 345454
rect 233486 345218 233528 345454
rect 233208 345134 233528 345218
rect 233208 344898 233250 345134
rect 233486 344898 233528 345134
rect 233208 344866 233528 344898
rect 243448 345454 243768 345486
rect 243448 345218 243490 345454
rect 243726 345218 243768 345454
rect 243448 345134 243768 345218
rect 243448 344898 243490 345134
rect 243726 344898 243768 345134
rect 243448 344866 243768 344898
rect 253688 345454 254008 345486
rect 253688 345218 253730 345454
rect 253966 345218 254008 345454
rect 253688 345134 254008 345218
rect 253688 344898 253730 345134
rect 253966 344898 254008 345134
rect 253688 344866 254008 344898
rect 263928 345454 264248 345486
rect 263928 345218 263970 345454
rect 264206 345218 264248 345454
rect 263928 345134 264248 345218
rect 263928 344898 263970 345134
rect 264206 344898 264248 345134
rect 263928 344866 264248 344898
rect 274168 345454 274488 345486
rect 274168 345218 274210 345454
rect 274446 345218 274488 345454
rect 274168 345134 274488 345218
rect 274168 344898 274210 345134
rect 274446 344898 274488 345134
rect 274168 344866 274488 344898
rect 284408 345454 284728 345486
rect 284408 345218 284450 345454
rect 284686 345218 284728 345454
rect 284408 345134 284728 345218
rect 284408 344898 284450 345134
rect 284686 344898 284728 345134
rect 284408 344866 284728 344898
rect 294648 345454 294968 345486
rect 294648 345218 294690 345454
rect 294926 345218 294968 345454
rect 294648 345134 294968 345218
rect 294648 344898 294690 345134
rect 294926 344898 294968 345134
rect 294648 344866 294968 344898
rect 304888 345454 305208 345486
rect 304888 345218 304930 345454
rect 305166 345218 305208 345454
rect 304888 345134 305208 345218
rect 304888 344898 304930 345134
rect 305166 344898 305208 345134
rect 304888 344866 305208 344898
rect 315128 345454 315448 345486
rect 315128 345218 315170 345454
rect 315406 345218 315448 345454
rect 315128 345134 315448 345218
rect 315128 344898 315170 345134
rect 315406 344898 315448 345134
rect 315128 344866 315448 344898
rect 325368 345454 325688 345486
rect 325368 345218 325410 345454
rect 325646 345218 325688 345454
rect 325368 345134 325688 345218
rect 325368 344898 325410 345134
rect 325646 344898 325688 345134
rect 325368 344866 325688 344898
rect 335608 345454 335928 345486
rect 335608 345218 335650 345454
rect 335886 345218 335928 345454
rect 335608 345134 335928 345218
rect 335608 344898 335650 345134
rect 335886 344898 335928 345134
rect 335608 344866 335928 344898
rect 345848 345454 346168 345486
rect 345848 345218 345890 345454
rect 346126 345218 346168 345454
rect 345848 345134 346168 345218
rect 345848 344898 345890 345134
rect 346126 344898 346168 345134
rect 345848 344866 346168 344898
rect 356088 345454 356408 345486
rect 356088 345218 356130 345454
rect 356366 345218 356408 345454
rect 356088 345134 356408 345218
rect 356088 344898 356130 345134
rect 356366 344898 356408 345134
rect 356088 344866 356408 344898
rect 366328 345454 366648 345486
rect 366328 345218 366370 345454
rect 366606 345218 366648 345454
rect 366328 345134 366648 345218
rect 366328 344898 366370 345134
rect 366606 344898 366648 345134
rect 366328 344866 366648 344898
rect 376568 345454 376888 345486
rect 376568 345218 376610 345454
rect 376846 345218 376888 345454
rect 376568 345134 376888 345218
rect 376568 344898 376610 345134
rect 376846 344898 376888 345134
rect 376568 344866 376888 344898
rect 386808 345454 387128 345486
rect 386808 345218 386850 345454
rect 387086 345218 387128 345454
rect 386808 345134 387128 345218
rect 386808 344898 386850 345134
rect 387086 344898 387128 345134
rect 386808 344866 387128 344898
rect 397048 345454 397368 345486
rect 397048 345218 397090 345454
rect 397326 345218 397368 345454
rect 397048 345134 397368 345218
rect 397048 344898 397090 345134
rect 397326 344898 397368 345134
rect 397048 344866 397368 344898
rect 407288 345454 407608 345486
rect 407288 345218 407330 345454
rect 407566 345218 407608 345454
rect 407288 345134 407608 345218
rect 407288 344898 407330 345134
rect 407566 344898 407608 345134
rect 407288 344866 407608 344898
rect 417528 345454 417848 345486
rect 417528 345218 417570 345454
rect 417806 345218 417848 345454
rect 417528 345134 417848 345218
rect 417528 344898 417570 345134
rect 417806 344898 417848 345134
rect 417528 344866 417848 344898
rect 427768 345454 428088 345486
rect 427768 345218 427810 345454
rect 428046 345218 428088 345454
rect 427768 345134 428088 345218
rect 427768 344898 427810 345134
rect 428046 344898 428088 345134
rect 427768 344866 428088 344898
rect 438008 345454 438328 345486
rect 438008 345218 438050 345454
rect 438286 345218 438328 345454
rect 438008 345134 438328 345218
rect 438008 344898 438050 345134
rect 438286 344898 438328 345134
rect 438008 344866 438328 344898
rect 448248 345454 448568 345486
rect 448248 345218 448290 345454
rect 448526 345218 448568 345454
rect 448248 345134 448568 345218
rect 448248 344898 448290 345134
rect 448526 344898 448568 345134
rect 448248 344866 448568 344898
rect 458488 345454 458808 345486
rect 458488 345218 458530 345454
rect 458766 345218 458808 345454
rect 458488 345134 458808 345218
rect 458488 344898 458530 345134
rect 458766 344898 458808 345134
rect 458488 344866 458808 344898
rect 468728 345454 469048 345486
rect 468728 345218 468770 345454
rect 469006 345218 469048 345454
rect 468728 345134 469048 345218
rect 468728 344898 468770 345134
rect 469006 344898 469048 345134
rect 468728 344866 469048 344898
rect 478968 345454 479288 345486
rect 478968 345218 479010 345454
rect 479246 345218 479288 345454
rect 478968 345134 479288 345218
rect 478968 344898 479010 345134
rect 479246 344898 479288 345134
rect 478968 344866 479288 344898
rect 489208 345454 489528 345486
rect 489208 345218 489250 345454
rect 489486 345218 489528 345454
rect 489208 345134 489528 345218
rect 489208 344898 489250 345134
rect 489486 344898 489528 345134
rect 489208 344866 489528 344898
rect 499448 345454 499768 345486
rect 499448 345218 499490 345454
rect 499726 345218 499768 345454
rect 499448 345134 499768 345218
rect 499448 344898 499490 345134
rect 499726 344898 499768 345134
rect 499448 344866 499768 344898
rect 509688 345454 510008 345486
rect 509688 345218 509730 345454
rect 509966 345218 510008 345454
rect 509688 345134 510008 345218
rect 509688 344898 509730 345134
rect 509966 344898 510008 345134
rect 509688 344866 510008 344898
rect 519928 345454 520248 345486
rect 519928 345218 519970 345454
rect 520206 345218 520248 345454
rect 519928 345134 520248 345218
rect 519928 344898 519970 345134
rect 520206 344898 520248 345134
rect 519928 344866 520248 344898
rect 530168 345454 530488 345486
rect 530168 345218 530210 345454
rect 530446 345218 530488 345454
rect 530168 345134 530488 345218
rect 530168 344898 530210 345134
rect 530446 344898 530488 345134
rect 530168 344866 530488 344898
rect 15754 330938 15786 331174
rect 16022 330938 16106 331174
rect 16342 330938 16374 331174
rect 15754 330854 16374 330938
rect 15754 330618 15786 330854
rect 16022 330618 16106 330854
rect 16342 330618 16374 330854
rect 15754 295174 16374 330618
rect 541714 334894 542334 370338
rect 541714 334658 541746 334894
rect 541982 334658 542066 334894
rect 542302 334658 542334 334894
rect 541714 334574 542334 334658
rect 541714 334338 541746 334574
rect 541982 334338 542066 334574
rect 542302 334338 542334 334574
rect 23288 327454 23608 327486
rect 23288 327218 23330 327454
rect 23566 327218 23608 327454
rect 23288 327134 23608 327218
rect 23288 326898 23330 327134
rect 23566 326898 23608 327134
rect 23288 326866 23608 326898
rect 33528 327454 33848 327486
rect 33528 327218 33570 327454
rect 33806 327218 33848 327454
rect 33528 327134 33848 327218
rect 33528 326898 33570 327134
rect 33806 326898 33848 327134
rect 33528 326866 33848 326898
rect 43768 327454 44088 327486
rect 43768 327218 43810 327454
rect 44046 327218 44088 327454
rect 43768 327134 44088 327218
rect 43768 326898 43810 327134
rect 44046 326898 44088 327134
rect 43768 326866 44088 326898
rect 54008 327454 54328 327486
rect 54008 327218 54050 327454
rect 54286 327218 54328 327454
rect 54008 327134 54328 327218
rect 54008 326898 54050 327134
rect 54286 326898 54328 327134
rect 54008 326866 54328 326898
rect 64248 327454 64568 327486
rect 64248 327218 64290 327454
rect 64526 327218 64568 327454
rect 64248 327134 64568 327218
rect 64248 326898 64290 327134
rect 64526 326898 64568 327134
rect 64248 326866 64568 326898
rect 74488 327454 74808 327486
rect 74488 327218 74530 327454
rect 74766 327218 74808 327454
rect 74488 327134 74808 327218
rect 74488 326898 74530 327134
rect 74766 326898 74808 327134
rect 74488 326866 74808 326898
rect 84728 327454 85048 327486
rect 84728 327218 84770 327454
rect 85006 327218 85048 327454
rect 84728 327134 85048 327218
rect 84728 326898 84770 327134
rect 85006 326898 85048 327134
rect 84728 326866 85048 326898
rect 94968 327454 95288 327486
rect 94968 327218 95010 327454
rect 95246 327218 95288 327454
rect 94968 327134 95288 327218
rect 94968 326898 95010 327134
rect 95246 326898 95288 327134
rect 94968 326866 95288 326898
rect 105208 327454 105528 327486
rect 105208 327218 105250 327454
rect 105486 327218 105528 327454
rect 105208 327134 105528 327218
rect 105208 326898 105250 327134
rect 105486 326898 105528 327134
rect 105208 326866 105528 326898
rect 115448 327454 115768 327486
rect 115448 327218 115490 327454
rect 115726 327218 115768 327454
rect 115448 327134 115768 327218
rect 115448 326898 115490 327134
rect 115726 326898 115768 327134
rect 115448 326866 115768 326898
rect 125688 327454 126008 327486
rect 125688 327218 125730 327454
rect 125966 327218 126008 327454
rect 125688 327134 126008 327218
rect 125688 326898 125730 327134
rect 125966 326898 126008 327134
rect 125688 326866 126008 326898
rect 135928 327454 136248 327486
rect 135928 327218 135970 327454
rect 136206 327218 136248 327454
rect 135928 327134 136248 327218
rect 135928 326898 135970 327134
rect 136206 326898 136248 327134
rect 135928 326866 136248 326898
rect 146168 327454 146488 327486
rect 146168 327218 146210 327454
rect 146446 327218 146488 327454
rect 146168 327134 146488 327218
rect 146168 326898 146210 327134
rect 146446 326898 146488 327134
rect 146168 326866 146488 326898
rect 156408 327454 156728 327486
rect 156408 327218 156450 327454
rect 156686 327218 156728 327454
rect 156408 327134 156728 327218
rect 156408 326898 156450 327134
rect 156686 326898 156728 327134
rect 156408 326866 156728 326898
rect 166648 327454 166968 327486
rect 166648 327218 166690 327454
rect 166926 327218 166968 327454
rect 166648 327134 166968 327218
rect 166648 326898 166690 327134
rect 166926 326898 166968 327134
rect 166648 326866 166968 326898
rect 176888 327454 177208 327486
rect 176888 327218 176930 327454
rect 177166 327218 177208 327454
rect 176888 327134 177208 327218
rect 176888 326898 176930 327134
rect 177166 326898 177208 327134
rect 176888 326866 177208 326898
rect 187128 327454 187448 327486
rect 187128 327218 187170 327454
rect 187406 327218 187448 327454
rect 187128 327134 187448 327218
rect 187128 326898 187170 327134
rect 187406 326898 187448 327134
rect 187128 326866 187448 326898
rect 197368 327454 197688 327486
rect 197368 327218 197410 327454
rect 197646 327218 197688 327454
rect 197368 327134 197688 327218
rect 197368 326898 197410 327134
rect 197646 326898 197688 327134
rect 197368 326866 197688 326898
rect 207608 327454 207928 327486
rect 207608 327218 207650 327454
rect 207886 327218 207928 327454
rect 207608 327134 207928 327218
rect 207608 326898 207650 327134
rect 207886 326898 207928 327134
rect 207608 326866 207928 326898
rect 217848 327454 218168 327486
rect 217848 327218 217890 327454
rect 218126 327218 218168 327454
rect 217848 327134 218168 327218
rect 217848 326898 217890 327134
rect 218126 326898 218168 327134
rect 217848 326866 218168 326898
rect 228088 327454 228408 327486
rect 228088 327218 228130 327454
rect 228366 327218 228408 327454
rect 228088 327134 228408 327218
rect 228088 326898 228130 327134
rect 228366 326898 228408 327134
rect 228088 326866 228408 326898
rect 238328 327454 238648 327486
rect 238328 327218 238370 327454
rect 238606 327218 238648 327454
rect 238328 327134 238648 327218
rect 238328 326898 238370 327134
rect 238606 326898 238648 327134
rect 238328 326866 238648 326898
rect 248568 327454 248888 327486
rect 248568 327218 248610 327454
rect 248846 327218 248888 327454
rect 248568 327134 248888 327218
rect 248568 326898 248610 327134
rect 248846 326898 248888 327134
rect 248568 326866 248888 326898
rect 258808 327454 259128 327486
rect 258808 327218 258850 327454
rect 259086 327218 259128 327454
rect 258808 327134 259128 327218
rect 258808 326898 258850 327134
rect 259086 326898 259128 327134
rect 258808 326866 259128 326898
rect 269048 327454 269368 327486
rect 269048 327218 269090 327454
rect 269326 327218 269368 327454
rect 269048 327134 269368 327218
rect 269048 326898 269090 327134
rect 269326 326898 269368 327134
rect 269048 326866 269368 326898
rect 279288 327454 279608 327486
rect 279288 327218 279330 327454
rect 279566 327218 279608 327454
rect 279288 327134 279608 327218
rect 279288 326898 279330 327134
rect 279566 326898 279608 327134
rect 279288 326866 279608 326898
rect 289528 327454 289848 327486
rect 289528 327218 289570 327454
rect 289806 327218 289848 327454
rect 289528 327134 289848 327218
rect 289528 326898 289570 327134
rect 289806 326898 289848 327134
rect 289528 326866 289848 326898
rect 299768 327454 300088 327486
rect 299768 327218 299810 327454
rect 300046 327218 300088 327454
rect 299768 327134 300088 327218
rect 299768 326898 299810 327134
rect 300046 326898 300088 327134
rect 299768 326866 300088 326898
rect 310008 327454 310328 327486
rect 310008 327218 310050 327454
rect 310286 327218 310328 327454
rect 310008 327134 310328 327218
rect 310008 326898 310050 327134
rect 310286 326898 310328 327134
rect 310008 326866 310328 326898
rect 320248 327454 320568 327486
rect 320248 327218 320290 327454
rect 320526 327218 320568 327454
rect 320248 327134 320568 327218
rect 320248 326898 320290 327134
rect 320526 326898 320568 327134
rect 320248 326866 320568 326898
rect 330488 327454 330808 327486
rect 330488 327218 330530 327454
rect 330766 327218 330808 327454
rect 330488 327134 330808 327218
rect 330488 326898 330530 327134
rect 330766 326898 330808 327134
rect 330488 326866 330808 326898
rect 340728 327454 341048 327486
rect 340728 327218 340770 327454
rect 341006 327218 341048 327454
rect 340728 327134 341048 327218
rect 340728 326898 340770 327134
rect 341006 326898 341048 327134
rect 340728 326866 341048 326898
rect 350968 327454 351288 327486
rect 350968 327218 351010 327454
rect 351246 327218 351288 327454
rect 350968 327134 351288 327218
rect 350968 326898 351010 327134
rect 351246 326898 351288 327134
rect 350968 326866 351288 326898
rect 361208 327454 361528 327486
rect 361208 327218 361250 327454
rect 361486 327218 361528 327454
rect 361208 327134 361528 327218
rect 361208 326898 361250 327134
rect 361486 326898 361528 327134
rect 361208 326866 361528 326898
rect 371448 327454 371768 327486
rect 371448 327218 371490 327454
rect 371726 327218 371768 327454
rect 371448 327134 371768 327218
rect 371448 326898 371490 327134
rect 371726 326898 371768 327134
rect 371448 326866 371768 326898
rect 381688 327454 382008 327486
rect 381688 327218 381730 327454
rect 381966 327218 382008 327454
rect 381688 327134 382008 327218
rect 381688 326898 381730 327134
rect 381966 326898 382008 327134
rect 381688 326866 382008 326898
rect 391928 327454 392248 327486
rect 391928 327218 391970 327454
rect 392206 327218 392248 327454
rect 391928 327134 392248 327218
rect 391928 326898 391970 327134
rect 392206 326898 392248 327134
rect 391928 326866 392248 326898
rect 402168 327454 402488 327486
rect 402168 327218 402210 327454
rect 402446 327218 402488 327454
rect 402168 327134 402488 327218
rect 402168 326898 402210 327134
rect 402446 326898 402488 327134
rect 402168 326866 402488 326898
rect 412408 327454 412728 327486
rect 412408 327218 412450 327454
rect 412686 327218 412728 327454
rect 412408 327134 412728 327218
rect 412408 326898 412450 327134
rect 412686 326898 412728 327134
rect 412408 326866 412728 326898
rect 422648 327454 422968 327486
rect 422648 327218 422690 327454
rect 422926 327218 422968 327454
rect 422648 327134 422968 327218
rect 422648 326898 422690 327134
rect 422926 326898 422968 327134
rect 422648 326866 422968 326898
rect 432888 327454 433208 327486
rect 432888 327218 432930 327454
rect 433166 327218 433208 327454
rect 432888 327134 433208 327218
rect 432888 326898 432930 327134
rect 433166 326898 433208 327134
rect 432888 326866 433208 326898
rect 443128 327454 443448 327486
rect 443128 327218 443170 327454
rect 443406 327218 443448 327454
rect 443128 327134 443448 327218
rect 443128 326898 443170 327134
rect 443406 326898 443448 327134
rect 443128 326866 443448 326898
rect 453368 327454 453688 327486
rect 453368 327218 453410 327454
rect 453646 327218 453688 327454
rect 453368 327134 453688 327218
rect 453368 326898 453410 327134
rect 453646 326898 453688 327134
rect 453368 326866 453688 326898
rect 463608 327454 463928 327486
rect 463608 327218 463650 327454
rect 463886 327218 463928 327454
rect 463608 327134 463928 327218
rect 463608 326898 463650 327134
rect 463886 326898 463928 327134
rect 463608 326866 463928 326898
rect 473848 327454 474168 327486
rect 473848 327218 473890 327454
rect 474126 327218 474168 327454
rect 473848 327134 474168 327218
rect 473848 326898 473890 327134
rect 474126 326898 474168 327134
rect 473848 326866 474168 326898
rect 484088 327454 484408 327486
rect 484088 327218 484130 327454
rect 484366 327218 484408 327454
rect 484088 327134 484408 327218
rect 484088 326898 484130 327134
rect 484366 326898 484408 327134
rect 484088 326866 484408 326898
rect 494328 327454 494648 327486
rect 494328 327218 494370 327454
rect 494606 327218 494648 327454
rect 494328 327134 494648 327218
rect 494328 326898 494370 327134
rect 494606 326898 494648 327134
rect 494328 326866 494648 326898
rect 504568 327454 504888 327486
rect 504568 327218 504610 327454
rect 504846 327218 504888 327454
rect 504568 327134 504888 327218
rect 504568 326898 504610 327134
rect 504846 326898 504888 327134
rect 504568 326866 504888 326898
rect 514808 327454 515128 327486
rect 514808 327218 514850 327454
rect 515086 327218 515128 327454
rect 514808 327134 515128 327218
rect 514808 326898 514850 327134
rect 515086 326898 515128 327134
rect 514808 326866 515128 326898
rect 525048 327454 525368 327486
rect 525048 327218 525090 327454
rect 525326 327218 525368 327454
rect 525048 327134 525368 327218
rect 525048 326898 525090 327134
rect 525326 326898 525368 327134
rect 525048 326866 525368 326898
rect 535288 327454 535608 327486
rect 535288 327218 535330 327454
rect 535566 327218 535608 327454
rect 535288 327134 535608 327218
rect 535288 326898 535330 327134
rect 535566 326898 535608 327134
rect 535288 326866 535608 326898
rect 28408 309454 28728 309486
rect 28408 309218 28450 309454
rect 28686 309218 28728 309454
rect 28408 309134 28728 309218
rect 28408 308898 28450 309134
rect 28686 308898 28728 309134
rect 28408 308866 28728 308898
rect 38648 309454 38968 309486
rect 38648 309218 38690 309454
rect 38926 309218 38968 309454
rect 38648 309134 38968 309218
rect 38648 308898 38690 309134
rect 38926 308898 38968 309134
rect 38648 308866 38968 308898
rect 48888 309454 49208 309486
rect 48888 309218 48930 309454
rect 49166 309218 49208 309454
rect 48888 309134 49208 309218
rect 48888 308898 48930 309134
rect 49166 308898 49208 309134
rect 48888 308866 49208 308898
rect 59128 309454 59448 309486
rect 59128 309218 59170 309454
rect 59406 309218 59448 309454
rect 59128 309134 59448 309218
rect 59128 308898 59170 309134
rect 59406 308898 59448 309134
rect 59128 308866 59448 308898
rect 69368 309454 69688 309486
rect 69368 309218 69410 309454
rect 69646 309218 69688 309454
rect 69368 309134 69688 309218
rect 69368 308898 69410 309134
rect 69646 308898 69688 309134
rect 69368 308866 69688 308898
rect 79608 309454 79928 309486
rect 79608 309218 79650 309454
rect 79886 309218 79928 309454
rect 79608 309134 79928 309218
rect 79608 308898 79650 309134
rect 79886 308898 79928 309134
rect 79608 308866 79928 308898
rect 89848 309454 90168 309486
rect 89848 309218 89890 309454
rect 90126 309218 90168 309454
rect 89848 309134 90168 309218
rect 89848 308898 89890 309134
rect 90126 308898 90168 309134
rect 89848 308866 90168 308898
rect 100088 309454 100408 309486
rect 100088 309218 100130 309454
rect 100366 309218 100408 309454
rect 100088 309134 100408 309218
rect 100088 308898 100130 309134
rect 100366 308898 100408 309134
rect 100088 308866 100408 308898
rect 110328 309454 110648 309486
rect 110328 309218 110370 309454
rect 110606 309218 110648 309454
rect 110328 309134 110648 309218
rect 110328 308898 110370 309134
rect 110606 308898 110648 309134
rect 110328 308866 110648 308898
rect 120568 309454 120888 309486
rect 120568 309218 120610 309454
rect 120846 309218 120888 309454
rect 120568 309134 120888 309218
rect 120568 308898 120610 309134
rect 120846 308898 120888 309134
rect 120568 308866 120888 308898
rect 130808 309454 131128 309486
rect 130808 309218 130850 309454
rect 131086 309218 131128 309454
rect 130808 309134 131128 309218
rect 130808 308898 130850 309134
rect 131086 308898 131128 309134
rect 130808 308866 131128 308898
rect 141048 309454 141368 309486
rect 141048 309218 141090 309454
rect 141326 309218 141368 309454
rect 141048 309134 141368 309218
rect 141048 308898 141090 309134
rect 141326 308898 141368 309134
rect 141048 308866 141368 308898
rect 151288 309454 151608 309486
rect 151288 309218 151330 309454
rect 151566 309218 151608 309454
rect 151288 309134 151608 309218
rect 151288 308898 151330 309134
rect 151566 308898 151608 309134
rect 151288 308866 151608 308898
rect 161528 309454 161848 309486
rect 161528 309218 161570 309454
rect 161806 309218 161848 309454
rect 161528 309134 161848 309218
rect 161528 308898 161570 309134
rect 161806 308898 161848 309134
rect 161528 308866 161848 308898
rect 171768 309454 172088 309486
rect 171768 309218 171810 309454
rect 172046 309218 172088 309454
rect 171768 309134 172088 309218
rect 171768 308898 171810 309134
rect 172046 308898 172088 309134
rect 171768 308866 172088 308898
rect 182008 309454 182328 309486
rect 182008 309218 182050 309454
rect 182286 309218 182328 309454
rect 182008 309134 182328 309218
rect 182008 308898 182050 309134
rect 182286 308898 182328 309134
rect 182008 308866 182328 308898
rect 192248 309454 192568 309486
rect 192248 309218 192290 309454
rect 192526 309218 192568 309454
rect 192248 309134 192568 309218
rect 192248 308898 192290 309134
rect 192526 308898 192568 309134
rect 192248 308866 192568 308898
rect 202488 309454 202808 309486
rect 202488 309218 202530 309454
rect 202766 309218 202808 309454
rect 202488 309134 202808 309218
rect 202488 308898 202530 309134
rect 202766 308898 202808 309134
rect 202488 308866 202808 308898
rect 212728 309454 213048 309486
rect 212728 309218 212770 309454
rect 213006 309218 213048 309454
rect 212728 309134 213048 309218
rect 212728 308898 212770 309134
rect 213006 308898 213048 309134
rect 212728 308866 213048 308898
rect 222968 309454 223288 309486
rect 222968 309218 223010 309454
rect 223246 309218 223288 309454
rect 222968 309134 223288 309218
rect 222968 308898 223010 309134
rect 223246 308898 223288 309134
rect 222968 308866 223288 308898
rect 233208 309454 233528 309486
rect 233208 309218 233250 309454
rect 233486 309218 233528 309454
rect 233208 309134 233528 309218
rect 233208 308898 233250 309134
rect 233486 308898 233528 309134
rect 233208 308866 233528 308898
rect 243448 309454 243768 309486
rect 243448 309218 243490 309454
rect 243726 309218 243768 309454
rect 243448 309134 243768 309218
rect 243448 308898 243490 309134
rect 243726 308898 243768 309134
rect 243448 308866 243768 308898
rect 253688 309454 254008 309486
rect 253688 309218 253730 309454
rect 253966 309218 254008 309454
rect 253688 309134 254008 309218
rect 253688 308898 253730 309134
rect 253966 308898 254008 309134
rect 253688 308866 254008 308898
rect 263928 309454 264248 309486
rect 263928 309218 263970 309454
rect 264206 309218 264248 309454
rect 263928 309134 264248 309218
rect 263928 308898 263970 309134
rect 264206 308898 264248 309134
rect 263928 308866 264248 308898
rect 274168 309454 274488 309486
rect 274168 309218 274210 309454
rect 274446 309218 274488 309454
rect 274168 309134 274488 309218
rect 274168 308898 274210 309134
rect 274446 308898 274488 309134
rect 274168 308866 274488 308898
rect 284408 309454 284728 309486
rect 284408 309218 284450 309454
rect 284686 309218 284728 309454
rect 284408 309134 284728 309218
rect 284408 308898 284450 309134
rect 284686 308898 284728 309134
rect 284408 308866 284728 308898
rect 294648 309454 294968 309486
rect 294648 309218 294690 309454
rect 294926 309218 294968 309454
rect 294648 309134 294968 309218
rect 294648 308898 294690 309134
rect 294926 308898 294968 309134
rect 294648 308866 294968 308898
rect 304888 309454 305208 309486
rect 304888 309218 304930 309454
rect 305166 309218 305208 309454
rect 304888 309134 305208 309218
rect 304888 308898 304930 309134
rect 305166 308898 305208 309134
rect 304888 308866 305208 308898
rect 315128 309454 315448 309486
rect 315128 309218 315170 309454
rect 315406 309218 315448 309454
rect 315128 309134 315448 309218
rect 315128 308898 315170 309134
rect 315406 308898 315448 309134
rect 315128 308866 315448 308898
rect 325368 309454 325688 309486
rect 325368 309218 325410 309454
rect 325646 309218 325688 309454
rect 325368 309134 325688 309218
rect 325368 308898 325410 309134
rect 325646 308898 325688 309134
rect 325368 308866 325688 308898
rect 335608 309454 335928 309486
rect 335608 309218 335650 309454
rect 335886 309218 335928 309454
rect 335608 309134 335928 309218
rect 335608 308898 335650 309134
rect 335886 308898 335928 309134
rect 335608 308866 335928 308898
rect 345848 309454 346168 309486
rect 345848 309218 345890 309454
rect 346126 309218 346168 309454
rect 345848 309134 346168 309218
rect 345848 308898 345890 309134
rect 346126 308898 346168 309134
rect 345848 308866 346168 308898
rect 356088 309454 356408 309486
rect 356088 309218 356130 309454
rect 356366 309218 356408 309454
rect 356088 309134 356408 309218
rect 356088 308898 356130 309134
rect 356366 308898 356408 309134
rect 356088 308866 356408 308898
rect 366328 309454 366648 309486
rect 366328 309218 366370 309454
rect 366606 309218 366648 309454
rect 366328 309134 366648 309218
rect 366328 308898 366370 309134
rect 366606 308898 366648 309134
rect 366328 308866 366648 308898
rect 376568 309454 376888 309486
rect 376568 309218 376610 309454
rect 376846 309218 376888 309454
rect 376568 309134 376888 309218
rect 376568 308898 376610 309134
rect 376846 308898 376888 309134
rect 376568 308866 376888 308898
rect 386808 309454 387128 309486
rect 386808 309218 386850 309454
rect 387086 309218 387128 309454
rect 386808 309134 387128 309218
rect 386808 308898 386850 309134
rect 387086 308898 387128 309134
rect 386808 308866 387128 308898
rect 397048 309454 397368 309486
rect 397048 309218 397090 309454
rect 397326 309218 397368 309454
rect 397048 309134 397368 309218
rect 397048 308898 397090 309134
rect 397326 308898 397368 309134
rect 397048 308866 397368 308898
rect 407288 309454 407608 309486
rect 407288 309218 407330 309454
rect 407566 309218 407608 309454
rect 407288 309134 407608 309218
rect 407288 308898 407330 309134
rect 407566 308898 407608 309134
rect 407288 308866 407608 308898
rect 417528 309454 417848 309486
rect 417528 309218 417570 309454
rect 417806 309218 417848 309454
rect 417528 309134 417848 309218
rect 417528 308898 417570 309134
rect 417806 308898 417848 309134
rect 417528 308866 417848 308898
rect 427768 309454 428088 309486
rect 427768 309218 427810 309454
rect 428046 309218 428088 309454
rect 427768 309134 428088 309218
rect 427768 308898 427810 309134
rect 428046 308898 428088 309134
rect 427768 308866 428088 308898
rect 438008 309454 438328 309486
rect 438008 309218 438050 309454
rect 438286 309218 438328 309454
rect 438008 309134 438328 309218
rect 438008 308898 438050 309134
rect 438286 308898 438328 309134
rect 438008 308866 438328 308898
rect 448248 309454 448568 309486
rect 448248 309218 448290 309454
rect 448526 309218 448568 309454
rect 448248 309134 448568 309218
rect 448248 308898 448290 309134
rect 448526 308898 448568 309134
rect 448248 308866 448568 308898
rect 458488 309454 458808 309486
rect 458488 309218 458530 309454
rect 458766 309218 458808 309454
rect 458488 309134 458808 309218
rect 458488 308898 458530 309134
rect 458766 308898 458808 309134
rect 458488 308866 458808 308898
rect 468728 309454 469048 309486
rect 468728 309218 468770 309454
rect 469006 309218 469048 309454
rect 468728 309134 469048 309218
rect 468728 308898 468770 309134
rect 469006 308898 469048 309134
rect 468728 308866 469048 308898
rect 478968 309454 479288 309486
rect 478968 309218 479010 309454
rect 479246 309218 479288 309454
rect 478968 309134 479288 309218
rect 478968 308898 479010 309134
rect 479246 308898 479288 309134
rect 478968 308866 479288 308898
rect 489208 309454 489528 309486
rect 489208 309218 489250 309454
rect 489486 309218 489528 309454
rect 489208 309134 489528 309218
rect 489208 308898 489250 309134
rect 489486 308898 489528 309134
rect 489208 308866 489528 308898
rect 499448 309454 499768 309486
rect 499448 309218 499490 309454
rect 499726 309218 499768 309454
rect 499448 309134 499768 309218
rect 499448 308898 499490 309134
rect 499726 308898 499768 309134
rect 499448 308866 499768 308898
rect 509688 309454 510008 309486
rect 509688 309218 509730 309454
rect 509966 309218 510008 309454
rect 509688 309134 510008 309218
rect 509688 308898 509730 309134
rect 509966 308898 510008 309134
rect 509688 308866 510008 308898
rect 519928 309454 520248 309486
rect 519928 309218 519970 309454
rect 520206 309218 520248 309454
rect 519928 309134 520248 309218
rect 519928 308898 519970 309134
rect 520206 308898 520248 309134
rect 519928 308866 520248 308898
rect 530168 309454 530488 309486
rect 530168 309218 530210 309454
rect 530446 309218 530488 309454
rect 530168 309134 530488 309218
rect 530168 308898 530210 309134
rect 530446 308898 530488 309134
rect 530168 308866 530488 308898
rect 15754 294938 15786 295174
rect 16022 294938 16106 295174
rect 16342 294938 16374 295174
rect 15754 294854 16374 294938
rect 15754 294618 15786 294854
rect 16022 294618 16106 294854
rect 16342 294618 16374 294854
rect 15754 259174 16374 294618
rect 541714 298894 542334 334338
rect 541714 298658 541746 298894
rect 541982 298658 542066 298894
rect 542302 298658 542334 298894
rect 541714 298574 542334 298658
rect 541714 298338 541746 298574
rect 541982 298338 542066 298574
rect 542302 298338 542334 298574
rect 23288 291454 23608 291486
rect 23288 291218 23330 291454
rect 23566 291218 23608 291454
rect 23288 291134 23608 291218
rect 23288 290898 23330 291134
rect 23566 290898 23608 291134
rect 23288 290866 23608 290898
rect 33528 291454 33848 291486
rect 33528 291218 33570 291454
rect 33806 291218 33848 291454
rect 33528 291134 33848 291218
rect 33528 290898 33570 291134
rect 33806 290898 33848 291134
rect 33528 290866 33848 290898
rect 43768 291454 44088 291486
rect 43768 291218 43810 291454
rect 44046 291218 44088 291454
rect 43768 291134 44088 291218
rect 43768 290898 43810 291134
rect 44046 290898 44088 291134
rect 43768 290866 44088 290898
rect 54008 291454 54328 291486
rect 54008 291218 54050 291454
rect 54286 291218 54328 291454
rect 54008 291134 54328 291218
rect 54008 290898 54050 291134
rect 54286 290898 54328 291134
rect 54008 290866 54328 290898
rect 64248 291454 64568 291486
rect 64248 291218 64290 291454
rect 64526 291218 64568 291454
rect 64248 291134 64568 291218
rect 64248 290898 64290 291134
rect 64526 290898 64568 291134
rect 64248 290866 64568 290898
rect 74488 291454 74808 291486
rect 74488 291218 74530 291454
rect 74766 291218 74808 291454
rect 74488 291134 74808 291218
rect 74488 290898 74530 291134
rect 74766 290898 74808 291134
rect 74488 290866 74808 290898
rect 84728 291454 85048 291486
rect 84728 291218 84770 291454
rect 85006 291218 85048 291454
rect 84728 291134 85048 291218
rect 84728 290898 84770 291134
rect 85006 290898 85048 291134
rect 84728 290866 85048 290898
rect 94968 291454 95288 291486
rect 94968 291218 95010 291454
rect 95246 291218 95288 291454
rect 94968 291134 95288 291218
rect 94968 290898 95010 291134
rect 95246 290898 95288 291134
rect 94968 290866 95288 290898
rect 105208 291454 105528 291486
rect 105208 291218 105250 291454
rect 105486 291218 105528 291454
rect 105208 291134 105528 291218
rect 105208 290898 105250 291134
rect 105486 290898 105528 291134
rect 105208 290866 105528 290898
rect 115448 291454 115768 291486
rect 115448 291218 115490 291454
rect 115726 291218 115768 291454
rect 115448 291134 115768 291218
rect 115448 290898 115490 291134
rect 115726 290898 115768 291134
rect 115448 290866 115768 290898
rect 125688 291454 126008 291486
rect 125688 291218 125730 291454
rect 125966 291218 126008 291454
rect 125688 291134 126008 291218
rect 125688 290898 125730 291134
rect 125966 290898 126008 291134
rect 125688 290866 126008 290898
rect 135928 291454 136248 291486
rect 135928 291218 135970 291454
rect 136206 291218 136248 291454
rect 135928 291134 136248 291218
rect 135928 290898 135970 291134
rect 136206 290898 136248 291134
rect 135928 290866 136248 290898
rect 146168 291454 146488 291486
rect 146168 291218 146210 291454
rect 146446 291218 146488 291454
rect 146168 291134 146488 291218
rect 146168 290898 146210 291134
rect 146446 290898 146488 291134
rect 146168 290866 146488 290898
rect 156408 291454 156728 291486
rect 156408 291218 156450 291454
rect 156686 291218 156728 291454
rect 156408 291134 156728 291218
rect 156408 290898 156450 291134
rect 156686 290898 156728 291134
rect 156408 290866 156728 290898
rect 166648 291454 166968 291486
rect 166648 291218 166690 291454
rect 166926 291218 166968 291454
rect 166648 291134 166968 291218
rect 166648 290898 166690 291134
rect 166926 290898 166968 291134
rect 166648 290866 166968 290898
rect 176888 291454 177208 291486
rect 176888 291218 176930 291454
rect 177166 291218 177208 291454
rect 176888 291134 177208 291218
rect 176888 290898 176930 291134
rect 177166 290898 177208 291134
rect 176888 290866 177208 290898
rect 187128 291454 187448 291486
rect 187128 291218 187170 291454
rect 187406 291218 187448 291454
rect 187128 291134 187448 291218
rect 187128 290898 187170 291134
rect 187406 290898 187448 291134
rect 187128 290866 187448 290898
rect 197368 291454 197688 291486
rect 197368 291218 197410 291454
rect 197646 291218 197688 291454
rect 197368 291134 197688 291218
rect 197368 290898 197410 291134
rect 197646 290898 197688 291134
rect 197368 290866 197688 290898
rect 207608 291454 207928 291486
rect 207608 291218 207650 291454
rect 207886 291218 207928 291454
rect 207608 291134 207928 291218
rect 207608 290898 207650 291134
rect 207886 290898 207928 291134
rect 207608 290866 207928 290898
rect 217848 291454 218168 291486
rect 217848 291218 217890 291454
rect 218126 291218 218168 291454
rect 217848 291134 218168 291218
rect 217848 290898 217890 291134
rect 218126 290898 218168 291134
rect 217848 290866 218168 290898
rect 228088 291454 228408 291486
rect 228088 291218 228130 291454
rect 228366 291218 228408 291454
rect 228088 291134 228408 291218
rect 228088 290898 228130 291134
rect 228366 290898 228408 291134
rect 228088 290866 228408 290898
rect 238328 291454 238648 291486
rect 238328 291218 238370 291454
rect 238606 291218 238648 291454
rect 238328 291134 238648 291218
rect 238328 290898 238370 291134
rect 238606 290898 238648 291134
rect 238328 290866 238648 290898
rect 248568 291454 248888 291486
rect 248568 291218 248610 291454
rect 248846 291218 248888 291454
rect 248568 291134 248888 291218
rect 248568 290898 248610 291134
rect 248846 290898 248888 291134
rect 248568 290866 248888 290898
rect 258808 291454 259128 291486
rect 258808 291218 258850 291454
rect 259086 291218 259128 291454
rect 258808 291134 259128 291218
rect 258808 290898 258850 291134
rect 259086 290898 259128 291134
rect 258808 290866 259128 290898
rect 269048 291454 269368 291486
rect 269048 291218 269090 291454
rect 269326 291218 269368 291454
rect 269048 291134 269368 291218
rect 269048 290898 269090 291134
rect 269326 290898 269368 291134
rect 269048 290866 269368 290898
rect 279288 291454 279608 291486
rect 279288 291218 279330 291454
rect 279566 291218 279608 291454
rect 279288 291134 279608 291218
rect 279288 290898 279330 291134
rect 279566 290898 279608 291134
rect 279288 290866 279608 290898
rect 289528 291454 289848 291486
rect 289528 291218 289570 291454
rect 289806 291218 289848 291454
rect 289528 291134 289848 291218
rect 289528 290898 289570 291134
rect 289806 290898 289848 291134
rect 289528 290866 289848 290898
rect 299768 291454 300088 291486
rect 299768 291218 299810 291454
rect 300046 291218 300088 291454
rect 299768 291134 300088 291218
rect 299768 290898 299810 291134
rect 300046 290898 300088 291134
rect 299768 290866 300088 290898
rect 310008 291454 310328 291486
rect 310008 291218 310050 291454
rect 310286 291218 310328 291454
rect 310008 291134 310328 291218
rect 310008 290898 310050 291134
rect 310286 290898 310328 291134
rect 310008 290866 310328 290898
rect 320248 291454 320568 291486
rect 320248 291218 320290 291454
rect 320526 291218 320568 291454
rect 320248 291134 320568 291218
rect 320248 290898 320290 291134
rect 320526 290898 320568 291134
rect 320248 290866 320568 290898
rect 330488 291454 330808 291486
rect 330488 291218 330530 291454
rect 330766 291218 330808 291454
rect 330488 291134 330808 291218
rect 330488 290898 330530 291134
rect 330766 290898 330808 291134
rect 330488 290866 330808 290898
rect 340728 291454 341048 291486
rect 340728 291218 340770 291454
rect 341006 291218 341048 291454
rect 340728 291134 341048 291218
rect 340728 290898 340770 291134
rect 341006 290898 341048 291134
rect 340728 290866 341048 290898
rect 350968 291454 351288 291486
rect 350968 291218 351010 291454
rect 351246 291218 351288 291454
rect 350968 291134 351288 291218
rect 350968 290898 351010 291134
rect 351246 290898 351288 291134
rect 350968 290866 351288 290898
rect 361208 291454 361528 291486
rect 361208 291218 361250 291454
rect 361486 291218 361528 291454
rect 361208 291134 361528 291218
rect 361208 290898 361250 291134
rect 361486 290898 361528 291134
rect 361208 290866 361528 290898
rect 371448 291454 371768 291486
rect 371448 291218 371490 291454
rect 371726 291218 371768 291454
rect 371448 291134 371768 291218
rect 371448 290898 371490 291134
rect 371726 290898 371768 291134
rect 371448 290866 371768 290898
rect 381688 291454 382008 291486
rect 381688 291218 381730 291454
rect 381966 291218 382008 291454
rect 381688 291134 382008 291218
rect 381688 290898 381730 291134
rect 381966 290898 382008 291134
rect 381688 290866 382008 290898
rect 391928 291454 392248 291486
rect 391928 291218 391970 291454
rect 392206 291218 392248 291454
rect 391928 291134 392248 291218
rect 391928 290898 391970 291134
rect 392206 290898 392248 291134
rect 391928 290866 392248 290898
rect 402168 291454 402488 291486
rect 402168 291218 402210 291454
rect 402446 291218 402488 291454
rect 402168 291134 402488 291218
rect 402168 290898 402210 291134
rect 402446 290898 402488 291134
rect 402168 290866 402488 290898
rect 412408 291454 412728 291486
rect 412408 291218 412450 291454
rect 412686 291218 412728 291454
rect 412408 291134 412728 291218
rect 412408 290898 412450 291134
rect 412686 290898 412728 291134
rect 412408 290866 412728 290898
rect 422648 291454 422968 291486
rect 422648 291218 422690 291454
rect 422926 291218 422968 291454
rect 422648 291134 422968 291218
rect 422648 290898 422690 291134
rect 422926 290898 422968 291134
rect 422648 290866 422968 290898
rect 432888 291454 433208 291486
rect 432888 291218 432930 291454
rect 433166 291218 433208 291454
rect 432888 291134 433208 291218
rect 432888 290898 432930 291134
rect 433166 290898 433208 291134
rect 432888 290866 433208 290898
rect 443128 291454 443448 291486
rect 443128 291218 443170 291454
rect 443406 291218 443448 291454
rect 443128 291134 443448 291218
rect 443128 290898 443170 291134
rect 443406 290898 443448 291134
rect 443128 290866 443448 290898
rect 453368 291454 453688 291486
rect 453368 291218 453410 291454
rect 453646 291218 453688 291454
rect 453368 291134 453688 291218
rect 453368 290898 453410 291134
rect 453646 290898 453688 291134
rect 453368 290866 453688 290898
rect 463608 291454 463928 291486
rect 463608 291218 463650 291454
rect 463886 291218 463928 291454
rect 463608 291134 463928 291218
rect 463608 290898 463650 291134
rect 463886 290898 463928 291134
rect 463608 290866 463928 290898
rect 473848 291454 474168 291486
rect 473848 291218 473890 291454
rect 474126 291218 474168 291454
rect 473848 291134 474168 291218
rect 473848 290898 473890 291134
rect 474126 290898 474168 291134
rect 473848 290866 474168 290898
rect 484088 291454 484408 291486
rect 484088 291218 484130 291454
rect 484366 291218 484408 291454
rect 484088 291134 484408 291218
rect 484088 290898 484130 291134
rect 484366 290898 484408 291134
rect 484088 290866 484408 290898
rect 494328 291454 494648 291486
rect 494328 291218 494370 291454
rect 494606 291218 494648 291454
rect 494328 291134 494648 291218
rect 494328 290898 494370 291134
rect 494606 290898 494648 291134
rect 494328 290866 494648 290898
rect 504568 291454 504888 291486
rect 504568 291218 504610 291454
rect 504846 291218 504888 291454
rect 504568 291134 504888 291218
rect 504568 290898 504610 291134
rect 504846 290898 504888 291134
rect 504568 290866 504888 290898
rect 514808 291454 515128 291486
rect 514808 291218 514850 291454
rect 515086 291218 515128 291454
rect 514808 291134 515128 291218
rect 514808 290898 514850 291134
rect 515086 290898 515128 291134
rect 514808 290866 515128 290898
rect 525048 291454 525368 291486
rect 525048 291218 525090 291454
rect 525326 291218 525368 291454
rect 525048 291134 525368 291218
rect 525048 290898 525090 291134
rect 525326 290898 525368 291134
rect 525048 290866 525368 290898
rect 535288 291454 535608 291486
rect 535288 291218 535330 291454
rect 535566 291218 535608 291454
rect 535288 291134 535608 291218
rect 535288 290898 535330 291134
rect 535566 290898 535608 291134
rect 535288 290866 535608 290898
rect 28408 273454 28728 273486
rect 28408 273218 28450 273454
rect 28686 273218 28728 273454
rect 28408 273134 28728 273218
rect 28408 272898 28450 273134
rect 28686 272898 28728 273134
rect 28408 272866 28728 272898
rect 38648 273454 38968 273486
rect 38648 273218 38690 273454
rect 38926 273218 38968 273454
rect 38648 273134 38968 273218
rect 38648 272898 38690 273134
rect 38926 272898 38968 273134
rect 38648 272866 38968 272898
rect 48888 273454 49208 273486
rect 48888 273218 48930 273454
rect 49166 273218 49208 273454
rect 48888 273134 49208 273218
rect 48888 272898 48930 273134
rect 49166 272898 49208 273134
rect 48888 272866 49208 272898
rect 59128 273454 59448 273486
rect 59128 273218 59170 273454
rect 59406 273218 59448 273454
rect 59128 273134 59448 273218
rect 59128 272898 59170 273134
rect 59406 272898 59448 273134
rect 59128 272866 59448 272898
rect 69368 273454 69688 273486
rect 69368 273218 69410 273454
rect 69646 273218 69688 273454
rect 69368 273134 69688 273218
rect 69368 272898 69410 273134
rect 69646 272898 69688 273134
rect 69368 272866 69688 272898
rect 79608 273454 79928 273486
rect 79608 273218 79650 273454
rect 79886 273218 79928 273454
rect 79608 273134 79928 273218
rect 79608 272898 79650 273134
rect 79886 272898 79928 273134
rect 79608 272866 79928 272898
rect 89848 273454 90168 273486
rect 89848 273218 89890 273454
rect 90126 273218 90168 273454
rect 89848 273134 90168 273218
rect 89848 272898 89890 273134
rect 90126 272898 90168 273134
rect 89848 272866 90168 272898
rect 100088 273454 100408 273486
rect 100088 273218 100130 273454
rect 100366 273218 100408 273454
rect 100088 273134 100408 273218
rect 100088 272898 100130 273134
rect 100366 272898 100408 273134
rect 100088 272866 100408 272898
rect 110328 273454 110648 273486
rect 110328 273218 110370 273454
rect 110606 273218 110648 273454
rect 110328 273134 110648 273218
rect 110328 272898 110370 273134
rect 110606 272898 110648 273134
rect 110328 272866 110648 272898
rect 120568 273454 120888 273486
rect 120568 273218 120610 273454
rect 120846 273218 120888 273454
rect 120568 273134 120888 273218
rect 120568 272898 120610 273134
rect 120846 272898 120888 273134
rect 120568 272866 120888 272898
rect 130808 273454 131128 273486
rect 130808 273218 130850 273454
rect 131086 273218 131128 273454
rect 130808 273134 131128 273218
rect 130808 272898 130850 273134
rect 131086 272898 131128 273134
rect 130808 272866 131128 272898
rect 141048 273454 141368 273486
rect 141048 273218 141090 273454
rect 141326 273218 141368 273454
rect 141048 273134 141368 273218
rect 141048 272898 141090 273134
rect 141326 272898 141368 273134
rect 141048 272866 141368 272898
rect 151288 273454 151608 273486
rect 151288 273218 151330 273454
rect 151566 273218 151608 273454
rect 151288 273134 151608 273218
rect 151288 272898 151330 273134
rect 151566 272898 151608 273134
rect 151288 272866 151608 272898
rect 161528 273454 161848 273486
rect 161528 273218 161570 273454
rect 161806 273218 161848 273454
rect 161528 273134 161848 273218
rect 161528 272898 161570 273134
rect 161806 272898 161848 273134
rect 161528 272866 161848 272898
rect 171768 273454 172088 273486
rect 171768 273218 171810 273454
rect 172046 273218 172088 273454
rect 171768 273134 172088 273218
rect 171768 272898 171810 273134
rect 172046 272898 172088 273134
rect 171768 272866 172088 272898
rect 182008 273454 182328 273486
rect 182008 273218 182050 273454
rect 182286 273218 182328 273454
rect 182008 273134 182328 273218
rect 182008 272898 182050 273134
rect 182286 272898 182328 273134
rect 182008 272866 182328 272898
rect 192248 273454 192568 273486
rect 192248 273218 192290 273454
rect 192526 273218 192568 273454
rect 192248 273134 192568 273218
rect 192248 272898 192290 273134
rect 192526 272898 192568 273134
rect 192248 272866 192568 272898
rect 202488 273454 202808 273486
rect 202488 273218 202530 273454
rect 202766 273218 202808 273454
rect 202488 273134 202808 273218
rect 202488 272898 202530 273134
rect 202766 272898 202808 273134
rect 202488 272866 202808 272898
rect 212728 273454 213048 273486
rect 212728 273218 212770 273454
rect 213006 273218 213048 273454
rect 212728 273134 213048 273218
rect 212728 272898 212770 273134
rect 213006 272898 213048 273134
rect 212728 272866 213048 272898
rect 222968 273454 223288 273486
rect 222968 273218 223010 273454
rect 223246 273218 223288 273454
rect 222968 273134 223288 273218
rect 222968 272898 223010 273134
rect 223246 272898 223288 273134
rect 222968 272866 223288 272898
rect 233208 273454 233528 273486
rect 233208 273218 233250 273454
rect 233486 273218 233528 273454
rect 233208 273134 233528 273218
rect 233208 272898 233250 273134
rect 233486 272898 233528 273134
rect 233208 272866 233528 272898
rect 243448 273454 243768 273486
rect 243448 273218 243490 273454
rect 243726 273218 243768 273454
rect 243448 273134 243768 273218
rect 243448 272898 243490 273134
rect 243726 272898 243768 273134
rect 243448 272866 243768 272898
rect 253688 273454 254008 273486
rect 253688 273218 253730 273454
rect 253966 273218 254008 273454
rect 253688 273134 254008 273218
rect 253688 272898 253730 273134
rect 253966 272898 254008 273134
rect 253688 272866 254008 272898
rect 263928 273454 264248 273486
rect 263928 273218 263970 273454
rect 264206 273218 264248 273454
rect 263928 273134 264248 273218
rect 263928 272898 263970 273134
rect 264206 272898 264248 273134
rect 263928 272866 264248 272898
rect 274168 273454 274488 273486
rect 274168 273218 274210 273454
rect 274446 273218 274488 273454
rect 274168 273134 274488 273218
rect 274168 272898 274210 273134
rect 274446 272898 274488 273134
rect 274168 272866 274488 272898
rect 284408 273454 284728 273486
rect 284408 273218 284450 273454
rect 284686 273218 284728 273454
rect 284408 273134 284728 273218
rect 284408 272898 284450 273134
rect 284686 272898 284728 273134
rect 284408 272866 284728 272898
rect 294648 273454 294968 273486
rect 294648 273218 294690 273454
rect 294926 273218 294968 273454
rect 294648 273134 294968 273218
rect 294648 272898 294690 273134
rect 294926 272898 294968 273134
rect 294648 272866 294968 272898
rect 304888 273454 305208 273486
rect 304888 273218 304930 273454
rect 305166 273218 305208 273454
rect 304888 273134 305208 273218
rect 304888 272898 304930 273134
rect 305166 272898 305208 273134
rect 304888 272866 305208 272898
rect 315128 273454 315448 273486
rect 315128 273218 315170 273454
rect 315406 273218 315448 273454
rect 315128 273134 315448 273218
rect 315128 272898 315170 273134
rect 315406 272898 315448 273134
rect 315128 272866 315448 272898
rect 325368 273454 325688 273486
rect 325368 273218 325410 273454
rect 325646 273218 325688 273454
rect 325368 273134 325688 273218
rect 325368 272898 325410 273134
rect 325646 272898 325688 273134
rect 325368 272866 325688 272898
rect 335608 273454 335928 273486
rect 335608 273218 335650 273454
rect 335886 273218 335928 273454
rect 335608 273134 335928 273218
rect 335608 272898 335650 273134
rect 335886 272898 335928 273134
rect 335608 272866 335928 272898
rect 345848 273454 346168 273486
rect 345848 273218 345890 273454
rect 346126 273218 346168 273454
rect 345848 273134 346168 273218
rect 345848 272898 345890 273134
rect 346126 272898 346168 273134
rect 345848 272866 346168 272898
rect 356088 273454 356408 273486
rect 356088 273218 356130 273454
rect 356366 273218 356408 273454
rect 356088 273134 356408 273218
rect 356088 272898 356130 273134
rect 356366 272898 356408 273134
rect 356088 272866 356408 272898
rect 366328 273454 366648 273486
rect 366328 273218 366370 273454
rect 366606 273218 366648 273454
rect 366328 273134 366648 273218
rect 366328 272898 366370 273134
rect 366606 272898 366648 273134
rect 366328 272866 366648 272898
rect 376568 273454 376888 273486
rect 376568 273218 376610 273454
rect 376846 273218 376888 273454
rect 376568 273134 376888 273218
rect 376568 272898 376610 273134
rect 376846 272898 376888 273134
rect 376568 272866 376888 272898
rect 386808 273454 387128 273486
rect 386808 273218 386850 273454
rect 387086 273218 387128 273454
rect 386808 273134 387128 273218
rect 386808 272898 386850 273134
rect 387086 272898 387128 273134
rect 386808 272866 387128 272898
rect 397048 273454 397368 273486
rect 397048 273218 397090 273454
rect 397326 273218 397368 273454
rect 397048 273134 397368 273218
rect 397048 272898 397090 273134
rect 397326 272898 397368 273134
rect 397048 272866 397368 272898
rect 407288 273454 407608 273486
rect 407288 273218 407330 273454
rect 407566 273218 407608 273454
rect 407288 273134 407608 273218
rect 407288 272898 407330 273134
rect 407566 272898 407608 273134
rect 407288 272866 407608 272898
rect 417528 273454 417848 273486
rect 417528 273218 417570 273454
rect 417806 273218 417848 273454
rect 417528 273134 417848 273218
rect 417528 272898 417570 273134
rect 417806 272898 417848 273134
rect 417528 272866 417848 272898
rect 427768 273454 428088 273486
rect 427768 273218 427810 273454
rect 428046 273218 428088 273454
rect 427768 273134 428088 273218
rect 427768 272898 427810 273134
rect 428046 272898 428088 273134
rect 427768 272866 428088 272898
rect 438008 273454 438328 273486
rect 438008 273218 438050 273454
rect 438286 273218 438328 273454
rect 438008 273134 438328 273218
rect 438008 272898 438050 273134
rect 438286 272898 438328 273134
rect 438008 272866 438328 272898
rect 448248 273454 448568 273486
rect 448248 273218 448290 273454
rect 448526 273218 448568 273454
rect 448248 273134 448568 273218
rect 448248 272898 448290 273134
rect 448526 272898 448568 273134
rect 448248 272866 448568 272898
rect 458488 273454 458808 273486
rect 458488 273218 458530 273454
rect 458766 273218 458808 273454
rect 458488 273134 458808 273218
rect 458488 272898 458530 273134
rect 458766 272898 458808 273134
rect 458488 272866 458808 272898
rect 468728 273454 469048 273486
rect 468728 273218 468770 273454
rect 469006 273218 469048 273454
rect 468728 273134 469048 273218
rect 468728 272898 468770 273134
rect 469006 272898 469048 273134
rect 468728 272866 469048 272898
rect 478968 273454 479288 273486
rect 478968 273218 479010 273454
rect 479246 273218 479288 273454
rect 478968 273134 479288 273218
rect 478968 272898 479010 273134
rect 479246 272898 479288 273134
rect 478968 272866 479288 272898
rect 489208 273454 489528 273486
rect 489208 273218 489250 273454
rect 489486 273218 489528 273454
rect 489208 273134 489528 273218
rect 489208 272898 489250 273134
rect 489486 272898 489528 273134
rect 489208 272866 489528 272898
rect 499448 273454 499768 273486
rect 499448 273218 499490 273454
rect 499726 273218 499768 273454
rect 499448 273134 499768 273218
rect 499448 272898 499490 273134
rect 499726 272898 499768 273134
rect 499448 272866 499768 272898
rect 509688 273454 510008 273486
rect 509688 273218 509730 273454
rect 509966 273218 510008 273454
rect 509688 273134 510008 273218
rect 509688 272898 509730 273134
rect 509966 272898 510008 273134
rect 509688 272866 510008 272898
rect 519928 273454 520248 273486
rect 519928 273218 519970 273454
rect 520206 273218 520248 273454
rect 519928 273134 520248 273218
rect 519928 272898 519970 273134
rect 520206 272898 520248 273134
rect 519928 272866 520248 272898
rect 530168 273454 530488 273486
rect 530168 273218 530210 273454
rect 530446 273218 530488 273454
rect 530168 273134 530488 273218
rect 530168 272898 530210 273134
rect 530446 272898 530488 273134
rect 530168 272866 530488 272898
rect 15754 258938 15786 259174
rect 16022 258938 16106 259174
rect 16342 258938 16374 259174
rect 15754 258854 16374 258938
rect 15754 258618 15786 258854
rect 16022 258618 16106 258854
rect 16342 258618 16374 258854
rect 15754 223174 16374 258618
rect 541714 262894 542334 298338
rect 541714 262658 541746 262894
rect 541982 262658 542066 262894
rect 542302 262658 542334 262894
rect 541714 262574 542334 262658
rect 541714 262338 541746 262574
rect 541982 262338 542066 262574
rect 542302 262338 542334 262574
rect 23288 255454 23608 255486
rect 23288 255218 23330 255454
rect 23566 255218 23608 255454
rect 23288 255134 23608 255218
rect 23288 254898 23330 255134
rect 23566 254898 23608 255134
rect 23288 254866 23608 254898
rect 33528 255454 33848 255486
rect 33528 255218 33570 255454
rect 33806 255218 33848 255454
rect 33528 255134 33848 255218
rect 33528 254898 33570 255134
rect 33806 254898 33848 255134
rect 33528 254866 33848 254898
rect 43768 255454 44088 255486
rect 43768 255218 43810 255454
rect 44046 255218 44088 255454
rect 43768 255134 44088 255218
rect 43768 254898 43810 255134
rect 44046 254898 44088 255134
rect 43768 254866 44088 254898
rect 54008 255454 54328 255486
rect 54008 255218 54050 255454
rect 54286 255218 54328 255454
rect 54008 255134 54328 255218
rect 54008 254898 54050 255134
rect 54286 254898 54328 255134
rect 54008 254866 54328 254898
rect 64248 255454 64568 255486
rect 64248 255218 64290 255454
rect 64526 255218 64568 255454
rect 64248 255134 64568 255218
rect 64248 254898 64290 255134
rect 64526 254898 64568 255134
rect 64248 254866 64568 254898
rect 74488 255454 74808 255486
rect 74488 255218 74530 255454
rect 74766 255218 74808 255454
rect 74488 255134 74808 255218
rect 74488 254898 74530 255134
rect 74766 254898 74808 255134
rect 74488 254866 74808 254898
rect 84728 255454 85048 255486
rect 84728 255218 84770 255454
rect 85006 255218 85048 255454
rect 84728 255134 85048 255218
rect 84728 254898 84770 255134
rect 85006 254898 85048 255134
rect 84728 254866 85048 254898
rect 94968 255454 95288 255486
rect 94968 255218 95010 255454
rect 95246 255218 95288 255454
rect 94968 255134 95288 255218
rect 94968 254898 95010 255134
rect 95246 254898 95288 255134
rect 94968 254866 95288 254898
rect 105208 255454 105528 255486
rect 105208 255218 105250 255454
rect 105486 255218 105528 255454
rect 105208 255134 105528 255218
rect 105208 254898 105250 255134
rect 105486 254898 105528 255134
rect 105208 254866 105528 254898
rect 115448 255454 115768 255486
rect 115448 255218 115490 255454
rect 115726 255218 115768 255454
rect 115448 255134 115768 255218
rect 115448 254898 115490 255134
rect 115726 254898 115768 255134
rect 115448 254866 115768 254898
rect 125688 255454 126008 255486
rect 125688 255218 125730 255454
rect 125966 255218 126008 255454
rect 125688 255134 126008 255218
rect 125688 254898 125730 255134
rect 125966 254898 126008 255134
rect 125688 254866 126008 254898
rect 135928 255454 136248 255486
rect 135928 255218 135970 255454
rect 136206 255218 136248 255454
rect 135928 255134 136248 255218
rect 135928 254898 135970 255134
rect 136206 254898 136248 255134
rect 135928 254866 136248 254898
rect 146168 255454 146488 255486
rect 146168 255218 146210 255454
rect 146446 255218 146488 255454
rect 146168 255134 146488 255218
rect 146168 254898 146210 255134
rect 146446 254898 146488 255134
rect 146168 254866 146488 254898
rect 156408 255454 156728 255486
rect 156408 255218 156450 255454
rect 156686 255218 156728 255454
rect 156408 255134 156728 255218
rect 156408 254898 156450 255134
rect 156686 254898 156728 255134
rect 156408 254866 156728 254898
rect 166648 255454 166968 255486
rect 166648 255218 166690 255454
rect 166926 255218 166968 255454
rect 166648 255134 166968 255218
rect 166648 254898 166690 255134
rect 166926 254898 166968 255134
rect 166648 254866 166968 254898
rect 176888 255454 177208 255486
rect 176888 255218 176930 255454
rect 177166 255218 177208 255454
rect 176888 255134 177208 255218
rect 176888 254898 176930 255134
rect 177166 254898 177208 255134
rect 176888 254866 177208 254898
rect 187128 255454 187448 255486
rect 187128 255218 187170 255454
rect 187406 255218 187448 255454
rect 187128 255134 187448 255218
rect 187128 254898 187170 255134
rect 187406 254898 187448 255134
rect 187128 254866 187448 254898
rect 197368 255454 197688 255486
rect 197368 255218 197410 255454
rect 197646 255218 197688 255454
rect 197368 255134 197688 255218
rect 197368 254898 197410 255134
rect 197646 254898 197688 255134
rect 197368 254866 197688 254898
rect 207608 255454 207928 255486
rect 207608 255218 207650 255454
rect 207886 255218 207928 255454
rect 207608 255134 207928 255218
rect 207608 254898 207650 255134
rect 207886 254898 207928 255134
rect 207608 254866 207928 254898
rect 217848 255454 218168 255486
rect 217848 255218 217890 255454
rect 218126 255218 218168 255454
rect 217848 255134 218168 255218
rect 217848 254898 217890 255134
rect 218126 254898 218168 255134
rect 217848 254866 218168 254898
rect 228088 255454 228408 255486
rect 228088 255218 228130 255454
rect 228366 255218 228408 255454
rect 228088 255134 228408 255218
rect 228088 254898 228130 255134
rect 228366 254898 228408 255134
rect 228088 254866 228408 254898
rect 238328 255454 238648 255486
rect 238328 255218 238370 255454
rect 238606 255218 238648 255454
rect 238328 255134 238648 255218
rect 238328 254898 238370 255134
rect 238606 254898 238648 255134
rect 238328 254866 238648 254898
rect 248568 255454 248888 255486
rect 248568 255218 248610 255454
rect 248846 255218 248888 255454
rect 248568 255134 248888 255218
rect 248568 254898 248610 255134
rect 248846 254898 248888 255134
rect 248568 254866 248888 254898
rect 258808 255454 259128 255486
rect 258808 255218 258850 255454
rect 259086 255218 259128 255454
rect 258808 255134 259128 255218
rect 258808 254898 258850 255134
rect 259086 254898 259128 255134
rect 258808 254866 259128 254898
rect 269048 255454 269368 255486
rect 269048 255218 269090 255454
rect 269326 255218 269368 255454
rect 269048 255134 269368 255218
rect 269048 254898 269090 255134
rect 269326 254898 269368 255134
rect 269048 254866 269368 254898
rect 279288 255454 279608 255486
rect 279288 255218 279330 255454
rect 279566 255218 279608 255454
rect 279288 255134 279608 255218
rect 279288 254898 279330 255134
rect 279566 254898 279608 255134
rect 279288 254866 279608 254898
rect 289528 255454 289848 255486
rect 289528 255218 289570 255454
rect 289806 255218 289848 255454
rect 289528 255134 289848 255218
rect 289528 254898 289570 255134
rect 289806 254898 289848 255134
rect 289528 254866 289848 254898
rect 299768 255454 300088 255486
rect 299768 255218 299810 255454
rect 300046 255218 300088 255454
rect 299768 255134 300088 255218
rect 299768 254898 299810 255134
rect 300046 254898 300088 255134
rect 299768 254866 300088 254898
rect 310008 255454 310328 255486
rect 310008 255218 310050 255454
rect 310286 255218 310328 255454
rect 310008 255134 310328 255218
rect 310008 254898 310050 255134
rect 310286 254898 310328 255134
rect 310008 254866 310328 254898
rect 320248 255454 320568 255486
rect 320248 255218 320290 255454
rect 320526 255218 320568 255454
rect 320248 255134 320568 255218
rect 320248 254898 320290 255134
rect 320526 254898 320568 255134
rect 320248 254866 320568 254898
rect 330488 255454 330808 255486
rect 330488 255218 330530 255454
rect 330766 255218 330808 255454
rect 330488 255134 330808 255218
rect 330488 254898 330530 255134
rect 330766 254898 330808 255134
rect 330488 254866 330808 254898
rect 340728 255454 341048 255486
rect 340728 255218 340770 255454
rect 341006 255218 341048 255454
rect 340728 255134 341048 255218
rect 340728 254898 340770 255134
rect 341006 254898 341048 255134
rect 340728 254866 341048 254898
rect 350968 255454 351288 255486
rect 350968 255218 351010 255454
rect 351246 255218 351288 255454
rect 350968 255134 351288 255218
rect 350968 254898 351010 255134
rect 351246 254898 351288 255134
rect 350968 254866 351288 254898
rect 361208 255454 361528 255486
rect 361208 255218 361250 255454
rect 361486 255218 361528 255454
rect 361208 255134 361528 255218
rect 361208 254898 361250 255134
rect 361486 254898 361528 255134
rect 361208 254866 361528 254898
rect 371448 255454 371768 255486
rect 371448 255218 371490 255454
rect 371726 255218 371768 255454
rect 371448 255134 371768 255218
rect 371448 254898 371490 255134
rect 371726 254898 371768 255134
rect 371448 254866 371768 254898
rect 381688 255454 382008 255486
rect 381688 255218 381730 255454
rect 381966 255218 382008 255454
rect 381688 255134 382008 255218
rect 381688 254898 381730 255134
rect 381966 254898 382008 255134
rect 381688 254866 382008 254898
rect 391928 255454 392248 255486
rect 391928 255218 391970 255454
rect 392206 255218 392248 255454
rect 391928 255134 392248 255218
rect 391928 254898 391970 255134
rect 392206 254898 392248 255134
rect 391928 254866 392248 254898
rect 402168 255454 402488 255486
rect 402168 255218 402210 255454
rect 402446 255218 402488 255454
rect 402168 255134 402488 255218
rect 402168 254898 402210 255134
rect 402446 254898 402488 255134
rect 402168 254866 402488 254898
rect 412408 255454 412728 255486
rect 412408 255218 412450 255454
rect 412686 255218 412728 255454
rect 412408 255134 412728 255218
rect 412408 254898 412450 255134
rect 412686 254898 412728 255134
rect 412408 254866 412728 254898
rect 422648 255454 422968 255486
rect 422648 255218 422690 255454
rect 422926 255218 422968 255454
rect 422648 255134 422968 255218
rect 422648 254898 422690 255134
rect 422926 254898 422968 255134
rect 422648 254866 422968 254898
rect 432888 255454 433208 255486
rect 432888 255218 432930 255454
rect 433166 255218 433208 255454
rect 432888 255134 433208 255218
rect 432888 254898 432930 255134
rect 433166 254898 433208 255134
rect 432888 254866 433208 254898
rect 443128 255454 443448 255486
rect 443128 255218 443170 255454
rect 443406 255218 443448 255454
rect 443128 255134 443448 255218
rect 443128 254898 443170 255134
rect 443406 254898 443448 255134
rect 443128 254866 443448 254898
rect 453368 255454 453688 255486
rect 453368 255218 453410 255454
rect 453646 255218 453688 255454
rect 453368 255134 453688 255218
rect 453368 254898 453410 255134
rect 453646 254898 453688 255134
rect 453368 254866 453688 254898
rect 463608 255454 463928 255486
rect 463608 255218 463650 255454
rect 463886 255218 463928 255454
rect 463608 255134 463928 255218
rect 463608 254898 463650 255134
rect 463886 254898 463928 255134
rect 463608 254866 463928 254898
rect 473848 255454 474168 255486
rect 473848 255218 473890 255454
rect 474126 255218 474168 255454
rect 473848 255134 474168 255218
rect 473848 254898 473890 255134
rect 474126 254898 474168 255134
rect 473848 254866 474168 254898
rect 484088 255454 484408 255486
rect 484088 255218 484130 255454
rect 484366 255218 484408 255454
rect 484088 255134 484408 255218
rect 484088 254898 484130 255134
rect 484366 254898 484408 255134
rect 484088 254866 484408 254898
rect 494328 255454 494648 255486
rect 494328 255218 494370 255454
rect 494606 255218 494648 255454
rect 494328 255134 494648 255218
rect 494328 254898 494370 255134
rect 494606 254898 494648 255134
rect 494328 254866 494648 254898
rect 504568 255454 504888 255486
rect 504568 255218 504610 255454
rect 504846 255218 504888 255454
rect 504568 255134 504888 255218
rect 504568 254898 504610 255134
rect 504846 254898 504888 255134
rect 504568 254866 504888 254898
rect 514808 255454 515128 255486
rect 514808 255218 514850 255454
rect 515086 255218 515128 255454
rect 514808 255134 515128 255218
rect 514808 254898 514850 255134
rect 515086 254898 515128 255134
rect 514808 254866 515128 254898
rect 525048 255454 525368 255486
rect 525048 255218 525090 255454
rect 525326 255218 525368 255454
rect 525048 255134 525368 255218
rect 525048 254898 525090 255134
rect 525326 254898 525368 255134
rect 525048 254866 525368 254898
rect 535288 255454 535608 255486
rect 535288 255218 535330 255454
rect 535566 255218 535608 255454
rect 535288 255134 535608 255218
rect 535288 254898 535330 255134
rect 535566 254898 535608 255134
rect 535288 254866 535608 254898
rect 28408 237454 28728 237486
rect 28408 237218 28450 237454
rect 28686 237218 28728 237454
rect 28408 237134 28728 237218
rect 28408 236898 28450 237134
rect 28686 236898 28728 237134
rect 28408 236866 28728 236898
rect 38648 237454 38968 237486
rect 38648 237218 38690 237454
rect 38926 237218 38968 237454
rect 38648 237134 38968 237218
rect 38648 236898 38690 237134
rect 38926 236898 38968 237134
rect 38648 236866 38968 236898
rect 48888 237454 49208 237486
rect 48888 237218 48930 237454
rect 49166 237218 49208 237454
rect 48888 237134 49208 237218
rect 48888 236898 48930 237134
rect 49166 236898 49208 237134
rect 48888 236866 49208 236898
rect 59128 237454 59448 237486
rect 59128 237218 59170 237454
rect 59406 237218 59448 237454
rect 59128 237134 59448 237218
rect 59128 236898 59170 237134
rect 59406 236898 59448 237134
rect 59128 236866 59448 236898
rect 69368 237454 69688 237486
rect 69368 237218 69410 237454
rect 69646 237218 69688 237454
rect 69368 237134 69688 237218
rect 69368 236898 69410 237134
rect 69646 236898 69688 237134
rect 69368 236866 69688 236898
rect 79608 237454 79928 237486
rect 79608 237218 79650 237454
rect 79886 237218 79928 237454
rect 79608 237134 79928 237218
rect 79608 236898 79650 237134
rect 79886 236898 79928 237134
rect 79608 236866 79928 236898
rect 89848 237454 90168 237486
rect 89848 237218 89890 237454
rect 90126 237218 90168 237454
rect 89848 237134 90168 237218
rect 89848 236898 89890 237134
rect 90126 236898 90168 237134
rect 89848 236866 90168 236898
rect 100088 237454 100408 237486
rect 100088 237218 100130 237454
rect 100366 237218 100408 237454
rect 100088 237134 100408 237218
rect 100088 236898 100130 237134
rect 100366 236898 100408 237134
rect 100088 236866 100408 236898
rect 110328 237454 110648 237486
rect 110328 237218 110370 237454
rect 110606 237218 110648 237454
rect 110328 237134 110648 237218
rect 110328 236898 110370 237134
rect 110606 236898 110648 237134
rect 110328 236866 110648 236898
rect 120568 237454 120888 237486
rect 120568 237218 120610 237454
rect 120846 237218 120888 237454
rect 120568 237134 120888 237218
rect 120568 236898 120610 237134
rect 120846 236898 120888 237134
rect 120568 236866 120888 236898
rect 130808 237454 131128 237486
rect 130808 237218 130850 237454
rect 131086 237218 131128 237454
rect 130808 237134 131128 237218
rect 130808 236898 130850 237134
rect 131086 236898 131128 237134
rect 130808 236866 131128 236898
rect 141048 237454 141368 237486
rect 141048 237218 141090 237454
rect 141326 237218 141368 237454
rect 141048 237134 141368 237218
rect 141048 236898 141090 237134
rect 141326 236898 141368 237134
rect 141048 236866 141368 236898
rect 151288 237454 151608 237486
rect 151288 237218 151330 237454
rect 151566 237218 151608 237454
rect 151288 237134 151608 237218
rect 151288 236898 151330 237134
rect 151566 236898 151608 237134
rect 151288 236866 151608 236898
rect 161528 237454 161848 237486
rect 161528 237218 161570 237454
rect 161806 237218 161848 237454
rect 161528 237134 161848 237218
rect 161528 236898 161570 237134
rect 161806 236898 161848 237134
rect 161528 236866 161848 236898
rect 171768 237454 172088 237486
rect 171768 237218 171810 237454
rect 172046 237218 172088 237454
rect 171768 237134 172088 237218
rect 171768 236898 171810 237134
rect 172046 236898 172088 237134
rect 171768 236866 172088 236898
rect 182008 237454 182328 237486
rect 182008 237218 182050 237454
rect 182286 237218 182328 237454
rect 182008 237134 182328 237218
rect 182008 236898 182050 237134
rect 182286 236898 182328 237134
rect 182008 236866 182328 236898
rect 192248 237454 192568 237486
rect 192248 237218 192290 237454
rect 192526 237218 192568 237454
rect 192248 237134 192568 237218
rect 192248 236898 192290 237134
rect 192526 236898 192568 237134
rect 192248 236866 192568 236898
rect 202488 237454 202808 237486
rect 202488 237218 202530 237454
rect 202766 237218 202808 237454
rect 202488 237134 202808 237218
rect 202488 236898 202530 237134
rect 202766 236898 202808 237134
rect 202488 236866 202808 236898
rect 212728 237454 213048 237486
rect 212728 237218 212770 237454
rect 213006 237218 213048 237454
rect 212728 237134 213048 237218
rect 212728 236898 212770 237134
rect 213006 236898 213048 237134
rect 212728 236866 213048 236898
rect 222968 237454 223288 237486
rect 222968 237218 223010 237454
rect 223246 237218 223288 237454
rect 222968 237134 223288 237218
rect 222968 236898 223010 237134
rect 223246 236898 223288 237134
rect 222968 236866 223288 236898
rect 233208 237454 233528 237486
rect 233208 237218 233250 237454
rect 233486 237218 233528 237454
rect 233208 237134 233528 237218
rect 233208 236898 233250 237134
rect 233486 236898 233528 237134
rect 233208 236866 233528 236898
rect 243448 237454 243768 237486
rect 243448 237218 243490 237454
rect 243726 237218 243768 237454
rect 243448 237134 243768 237218
rect 243448 236898 243490 237134
rect 243726 236898 243768 237134
rect 243448 236866 243768 236898
rect 253688 237454 254008 237486
rect 253688 237218 253730 237454
rect 253966 237218 254008 237454
rect 253688 237134 254008 237218
rect 253688 236898 253730 237134
rect 253966 236898 254008 237134
rect 253688 236866 254008 236898
rect 263928 237454 264248 237486
rect 263928 237218 263970 237454
rect 264206 237218 264248 237454
rect 263928 237134 264248 237218
rect 263928 236898 263970 237134
rect 264206 236898 264248 237134
rect 263928 236866 264248 236898
rect 274168 237454 274488 237486
rect 274168 237218 274210 237454
rect 274446 237218 274488 237454
rect 274168 237134 274488 237218
rect 274168 236898 274210 237134
rect 274446 236898 274488 237134
rect 274168 236866 274488 236898
rect 284408 237454 284728 237486
rect 284408 237218 284450 237454
rect 284686 237218 284728 237454
rect 284408 237134 284728 237218
rect 284408 236898 284450 237134
rect 284686 236898 284728 237134
rect 284408 236866 284728 236898
rect 294648 237454 294968 237486
rect 294648 237218 294690 237454
rect 294926 237218 294968 237454
rect 294648 237134 294968 237218
rect 294648 236898 294690 237134
rect 294926 236898 294968 237134
rect 294648 236866 294968 236898
rect 304888 237454 305208 237486
rect 304888 237218 304930 237454
rect 305166 237218 305208 237454
rect 304888 237134 305208 237218
rect 304888 236898 304930 237134
rect 305166 236898 305208 237134
rect 304888 236866 305208 236898
rect 315128 237454 315448 237486
rect 315128 237218 315170 237454
rect 315406 237218 315448 237454
rect 315128 237134 315448 237218
rect 315128 236898 315170 237134
rect 315406 236898 315448 237134
rect 315128 236866 315448 236898
rect 325368 237454 325688 237486
rect 325368 237218 325410 237454
rect 325646 237218 325688 237454
rect 325368 237134 325688 237218
rect 325368 236898 325410 237134
rect 325646 236898 325688 237134
rect 325368 236866 325688 236898
rect 335608 237454 335928 237486
rect 335608 237218 335650 237454
rect 335886 237218 335928 237454
rect 335608 237134 335928 237218
rect 335608 236898 335650 237134
rect 335886 236898 335928 237134
rect 335608 236866 335928 236898
rect 345848 237454 346168 237486
rect 345848 237218 345890 237454
rect 346126 237218 346168 237454
rect 345848 237134 346168 237218
rect 345848 236898 345890 237134
rect 346126 236898 346168 237134
rect 345848 236866 346168 236898
rect 356088 237454 356408 237486
rect 356088 237218 356130 237454
rect 356366 237218 356408 237454
rect 356088 237134 356408 237218
rect 356088 236898 356130 237134
rect 356366 236898 356408 237134
rect 356088 236866 356408 236898
rect 366328 237454 366648 237486
rect 366328 237218 366370 237454
rect 366606 237218 366648 237454
rect 366328 237134 366648 237218
rect 366328 236898 366370 237134
rect 366606 236898 366648 237134
rect 366328 236866 366648 236898
rect 376568 237454 376888 237486
rect 376568 237218 376610 237454
rect 376846 237218 376888 237454
rect 376568 237134 376888 237218
rect 376568 236898 376610 237134
rect 376846 236898 376888 237134
rect 376568 236866 376888 236898
rect 386808 237454 387128 237486
rect 386808 237218 386850 237454
rect 387086 237218 387128 237454
rect 386808 237134 387128 237218
rect 386808 236898 386850 237134
rect 387086 236898 387128 237134
rect 386808 236866 387128 236898
rect 397048 237454 397368 237486
rect 397048 237218 397090 237454
rect 397326 237218 397368 237454
rect 397048 237134 397368 237218
rect 397048 236898 397090 237134
rect 397326 236898 397368 237134
rect 397048 236866 397368 236898
rect 407288 237454 407608 237486
rect 407288 237218 407330 237454
rect 407566 237218 407608 237454
rect 407288 237134 407608 237218
rect 407288 236898 407330 237134
rect 407566 236898 407608 237134
rect 407288 236866 407608 236898
rect 417528 237454 417848 237486
rect 417528 237218 417570 237454
rect 417806 237218 417848 237454
rect 417528 237134 417848 237218
rect 417528 236898 417570 237134
rect 417806 236898 417848 237134
rect 417528 236866 417848 236898
rect 427768 237454 428088 237486
rect 427768 237218 427810 237454
rect 428046 237218 428088 237454
rect 427768 237134 428088 237218
rect 427768 236898 427810 237134
rect 428046 236898 428088 237134
rect 427768 236866 428088 236898
rect 438008 237454 438328 237486
rect 438008 237218 438050 237454
rect 438286 237218 438328 237454
rect 438008 237134 438328 237218
rect 438008 236898 438050 237134
rect 438286 236898 438328 237134
rect 438008 236866 438328 236898
rect 448248 237454 448568 237486
rect 448248 237218 448290 237454
rect 448526 237218 448568 237454
rect 448248 237134 448568 237218
rect 448248 236898 448290 237134
rect 448526 236898 448568 237134
rect 448248 236866 448568 236898
rect 458488 237454 458808 237486
rect 458488 237218 458530 237454
rect 458766 237218 458808 237454
rect 458488 237134 458808 237218
rect 458488 236898 458530 237134
rect 458766 236898 458808 237134
rect 458488 236866 458808 236898
rect 468728 237454 469048 237486
rect 468728 237218 468770 237454
rect 469006 237218 469048 237454
rect 468728 237134 469048 237218
rect 468728 236898 468770 237134
rect 469006 236898 469048 237134
rect 468728 236866 469048 236898
rect 478968 237454 479288 237486
rect 478968 237218 479010 237454
rect 479246 237218 479288 237454
rect 478968 237134 479288 237218
rect 478968 236898 479010 237134
rect 479246 236898 479288 237134
rect 478968 236866 479288 236898
rect 489208 237454 489528 237486
rect 489208 237218 489250 237454
rect 489486 237218 489528 237454
rect 489208 237134 489528 237218
rect 489208 236898 489250 237134
rect 489486 236898 489528 237134
rect 489208 236866 489528 236898
rect 499448 237454 499768 237486
rect 499448 237218 499490 237454
rect 499726 237218 499768 237454
rect 499448 237134 499768 237218
rect 499448 236898 499490 237134
rect 499726 236898 499768 237134
rect 499448 236866 499768 236898
rect 509688 237454 510008 237486
rect 509688 237218 509730 237454
rect 509966 237218 510008 237454
rect 509688 237134 510008 237218
rect 509688 236898 509730 237134
rect 509966 236898 510008 237134
rect 509688 236866 510008 236898
rect 519928 237454 520248 237486
rect 519928 237218 519970 237454
rect 520206 237218 520248 237454
rect 519928 237134 520248 237218
rect 519928 236898 519970 237134
rect 520206 236898 520248 237134
rect 519928 236866 520248 236898
rect 530168 237454 530488 237486
rect 530168 237218 530210 237454
rect 530446 237218 530488 237454
rect 530168 237134 530488 237218
rect 530168 236898 530210 237134
rect 530446 236898 530488 237134
rect 530168 236866 530488 236898
rect 15754 222938 15786 223174
rect 16022 222938 16106 223174
rect 16342 222938 16374 223174
rect 15754 222854 16374 222938
rect 15754 222618 15786 222854
rect 16022 222618 16106 222854
rect 16342 222618 16374 222854
rect 15754 187174 16374 222618
rect 541714 226894 542334 262338
rect 541714 226658 541746 226894
rect 541982 226658 542066 226894
rect 542302 226658 542334 226894
rect 541714 226574 542334 226658
rect 541714 226338 541746 226574
rect 541982 226338 542066 226574
rect 542302 226338 542334 226574
rect 23288 219454 23608 219486
rect 23288 219218 23330 219454
rect 23566 219218 23608 219454
rect 23288 219134 23608 219218
rect 23288 218898 23330 219134
rect 23566 218898 23608 219134
rect 23288 218866 23608 218898
rect 33528 219454 33848 219486
rect 33528 219218 33570 219454
rect 33806 219218 33848 219454
rect 33528 219134 33848 219218
rect 33528 218898 33570 219134
rect 33806 218898 33848 219134
rect 33528 218866 33848 218898
rect 43768 219454 44088 219486
rect 43768 219218 43810 219454
rect 44046 219218 44088 219454
rect 43768 219134 44088 219218
rect 43768 218898 43810 219134
rect 44046 218898 44088 219134
rect 43768 218866 44088 218898
rect 54008 219454 54328 219486
rect 54008 219218 54050 219454
rect 54286 219218 54328 219454
rect 54008 219134 54328 219218
rect 54008 218898 54050 219134
rect 54286 218898 54328 219134
rect 54008 218866 54328 218898
rect 64248 219454 64568 219486
rect 64248 219218 64290 219454
rect 64526 219218 64568 219454
rect 64248 219134 64568 219218
rect 64248 218898 64290 219134
rect 64526 218898 64568 219134
rect 64248 218866 64568 218898
rect 74488 219454 74808 219486
rect 74488 219218 74530 219454
rect 74766 219218 74808 219454
rect 74488 219134 74808 219218
rect 74488 218898 74530 219134
rect 74766 218898 74808 219134
rect 74488 218866 74808 218898
rect 84728 219454 85048 219486
rect 84728 219218 84770 219454
rect 85006 219218 85048 219454
rect 84728 219134 85048 219218
rect 84728 218898 84770 219134
rect 85006 218898 85048 219134
rect 84728 218866 85048 218898
rect 94968 219454 95288 219486
rect 94968 219218 95010 219454
rect 95246 219218 95288 219454
rect 94968 219134 95288 219218
rect 94968 218898 95010 219134
rect 95246 218898 95288 219134
rect 94968 218866 95288 218898
rect 105208 219454 105528 219486
rect 105208 219218 105250 219454
rect 105486 219218 105528 219454
rect 105208 219134 105528 219218
rect 105208 218898 105250 219134
rect 105486 218898 105528 219134
rect 105208 218866 105528 218898
rect 115448 219454 115768 219486
rect 115448 219218 115490 219454
rect 115726 219218 115768 219454
rect 115448 219134 115768 219218
rect 115448 218898 115490 219134
rect 115726 218898 115768 219134
rect 115448 218866 115768 218898
rect 125688 219454 126008 219486
rect 125688 219218 125730 219454
rect 125966 219218 126008 219454
rect 125688 219134 126008 219218
rect 125688 218898 125730 219134
rect 125966 218898 126008 219134
rect 125688 218866 126008 218898
rect 135928 219454 136248 219486
rect 135928 219218 135970 219454
rect 136206 219218 136248 219454
rect 135928 219134 136248 219218
rect 135928 218898 135970 219134
rect 136206 218898 136248 219134
rect 135928 218866 136248 218898
rect 146168 219454 146488 219486
rect 146168 219218 146210 219454
rect 146446 219218 146488 219454
rect 146168 219134 146488 219218
rect 146168 218898 146210 219134
rect 146446 218898 146488 219134
rect 146168 218866 146488 218898
rect 156408 219454 156728 219486
rect 156408 219218 156450 219454
rect 156686 219218 156728 219454
rect 156408 219134 156728 219218
rect 156408 218898 156450 219134
rect 156686 218898 156728 219134
rect 156408 218866 156728 218898
rect 166648 219454 166968 219486
rect 166648 219218 166690 219454
rect 166926 219218 166968 219454
rect 166648 219134 166968 219218
rect 166648 218898 166690 219134
rect 166926 218898 166968 219134
rect 166648 218866 166968 218898
rect 176888 219454 177208 219486
rect 176888 219218 176930 219454
rect 177166 219218 177208 219454
rect 176888 219134 177208 219218
rect 176888 218898 176930 219134
rect 177166 218898 177208 219134
rect 176888 218866 177208 218898
rect 187128 219454 187448 219486
rect 187128 219218 187170 219454
rect 187406 219218 187448 219454
rect 187128 219134 187448 219218
rect 187128 218898 187170 219134
rect 187406 218898 187448 219134
rect 187128 218866 187448 218898
rect 197368 219454 197688 219486
rect 197368 219218 197410 219454
rect 197646 219218 197688 219454
rect 197368 219134 197688 219218
rect 197368 218898 197410 219134
rect 197646 218898 197688 219134
rect 197368 218866 197688 218898
rect 207608 219454 207928 219486
rect 207608 219218 207650 219454
rect 207886 219218 207928 219454
rect 207608 219134 207928 219218
rect 207608 218898 207650 219134
rect 207886 218898 207928 219134
rect 207608 218866 207928 218898
rect 217848 219454 218168 219486
rect 217848 219218 217890 219454
rect 218126 219218 218168 219454
rect 217848 219134 218168 219218
rect 217848 218898 217890 219134
rect 218126 218898 218168 219134
rect 217848 218866 218168 218898
rect 228088 219454 228408 219486
rect 228088 219218 228130 219454
rect 228366 219218 228408 219454
rect 228088 219134 228408 219218
rect 228088 218898 228130 219134
rect 228366 218898 228408 219134
rect 228088 218866 228408 218898
rect 238328 219454 238648 219486
rect 238328 219218 238370 219454
rect 238606 219218 238648 219454
rect 238328 219134 238648 219218
rect 238328 218898 238370 219134
rect 238606 218898 238648 219134
rect 238328 218866 238648 218898
rect 248568 219454 248888 219486
rect 248568 219218 248610 219454
rect 248846 219218 248888 219454
rect 248568 219134 248888 219218
rect 248568 218898 248610 219134
rect 248846 218898 248888 219134
rect 248568 218866 248888 218898
rect 258808 219454 259128 219486
rect 258808 219218 258850 219454
rect 259086 219218 259128 219454
rect 258808 219134 259128 219218
rect 258808 218898 258850 219134
rect 259086 218898 259128 219134
rect 258808 218866 259128 218898
rect 269048 219454 269368 219486
rect 269048 219218 269090 219454
rect 269326 219218 269368 219454
rect 269048 219134 269368 219218
rect 269048 218898 269090 219134
rect 269326 218898 269368 219134
rect 269048 218866 269368 218898
rect 279288 219454 279608 219486
rect 279288 219218 279330 219454
rect 279566 219218 279608 219454
rect 279288 219134 279608 219218
rect 279288 218898 279330 219134
rect 279566 218898 279608 219134
rect 279288 218866 279608 218898
rect 289528 219454 289848 219486
rect 289528 219218 289570 219454
rect 289806 219218 289848 219454
rect 289528 219134 289848 219218
rect 289528 218898 289570 219134
rect 289806 218898 289848 219134
rect 289528 218866 289848 218898
rect 299768 219454 300088 219486
rect 299768 219218 299810 219454
rect 300046 219218 300088 219454
rect 299768 219134 300088 219218
rect 299768 218898 299810 219134
rect 300046 218898 300088 219134
rect 299768 218866 300088 218898
rect 310008 219454 310328 219486
rect 310008 219218 310050 219454
rect 310286 219218 310328 219454
rect 310008 219134 310328 219218
rect 310008 218898 310050 219134
rect 310286 218898 310328 219134
rect 310008 218866 310328 218898
rect 320248 219454 320568 219486
rect 320248 219218 320290 219454
rect 320526 219218 320568 219454
rect 320248 219134 320568 219218
rect 320248 218898 320290 219134
rect 320526 218898 320568 219134
rect 320248 218866 320568 218898
rect 330488 219454 330808 219486
rect 330488 219218 330530 219454
rect 330766 219218 330808 219454
rect 330488 219134 330808 219218
rect 330488 218898 330530 219134
rect 330766 218898 330808 219134
rect 330488 218866 330808 218898
rect 340728 219454 341048 219486
rect 340728 219218 340770 219454
rect 341006 219218 341048 219454
rect 340728 219134 341048 219218
rect 340728 218898 340770 219134
rect 341006 218898 341048 219134
rect 340728 218866 341048 218898
rect 350968 219454 351288 219486
rect 350968 219218 351010 219454
rect 351246 219218 351288 219454
rect 350968 219134 351288 219218
rect 350968 218898 351010 219134
rect 351246 218898 351288 219134
rect 350968 218866 351288 218898
rect 361208 219454 361528 219486
rect 361208 219218 361250 219454
rect 361486 219218 361528 219454
rect 361208 219134 361528 219218
rect 361208 218898 361250 219134
rect 361486 218898 361528 219134
rect 361208 218866 361528 218898
rect 371448 219454 371768 219486
rect 371448 219218 371490 219454
rect 371726 219218 371768 219454
rect 371448 219134 371768 219218
rect 371448 218898 371490 219134
rect 371726 218898 371768 219134
rect 371448 218866 371768 218898
rect 381688 219454 382008 219486
rect 381688 219218 381730 219454
rect 381966 219218 382008 219454
rect 381688 219134 382008 219218
rect 381688 218898 381730 219134
rect 381966 218898 382008 219134
rect 381688 218866 382008 218898
rect 391928 219454 392248 219486
rect 391928 219218 391970 219454
rect 392206 219218 392248 219454
rect 391928 219134 392248 219218
rect 391928 218898 391970 219134
rect 392206 218898 392248 219134
rect 391928 218866 392248 218898
rect 402168 219454 402488 219486
rect 402168 219218 402210 219454
rect 402446 219218 402488 219454
rect 402168 219134 402488 219218
rect 402168 218898 402210 219134
rect 402446 218898 402488 219134
rect 402168 218866 402488 218898
rect 412408 219454 412728 219486
rect 412408 219218 412450 219454
rect 412686 219218 412728 219454
rect 412408 219134 412728 219218
rect 412408 218898 412450 219134
rect 412686 218898 412728 219134
rect 412408 218866 412728 218898
rect 422648 219454 422968 219486
rect 422648 219218 422690 219454
rect 422926 219218 422968 219454
rect 422648 219134 422968 219218
rect 422648 218898 422690 219134
rect 422926 218898 422968 219134
rect 422648 218866 422968 218898
rect 432888 219454 433208 219486
rect 432888 219218 432930 219454
rect 433166 219218 433208 219454
rect 432888 219134 433208 219218
rect 432888 218898 432930 219134
rect 433166 218898 433208 219134
rect 432888 218866 433208 218898
rect 443128 219454 443448 219486
rect 443128 219218 443170 219454
rect 443406 219218 443448 219454
rect 443128 219134 443448 219218
rect 443128 218898 443170 219134
rect 443406 218898 443448 219134
rect 443128 218866 443448 218898
rect 453368 219454 453688 219486
rect 453368 219218 453410 219454
rect 453646 219218 453688 219454
rect 453368 219134 453688 219218
rect 453368 218898 453410 219134
rect 453646 218898 453688 219134
rect 453368 218866 453688 218898
rect 463608 219454 463928 219486
rect 463608 219218 463650 219454
rect 463886 219218 463928 219454
rect 463608 219134 463928 219218
rect 463608 218898 463650 219134
rect 463886 218898 463928 219134
rect 463608 218866 463928 218898
rect 473848 219454 474168 219486
rect 473848 219218 473890 219454
rect 474126 219218 474168 219454
rect 473848 219134 474168 219218
rect 473848 218898 473890 219134
rect 474126 218898 474168 219134
rect 473848 218866 474168 218898
rect 484088 219454 484408 219486
rect 484088 219218 484130 219454
rect 484366 219218 484408 219454
rect 484088 219134 484408 219218
rect 484088 218898 484130 219134
rect 484366 218898 484408 219134
rect 484088 218866 484408 218898
rect 494328 219454 494648 219486
rect 494328 219218 494370 219454
rect 494606 219218 494648 219454
rect 494328 219134 494648 219218
rect 494328 218898 494370 219134
rect 494606 218898 494648 219134
rect 494328 218866 494648 218898
rect 504568 219454 504888 219486
rect 504568 219218 504610 219454
rect 504846 219218 504888 219454
rect 504568 219134 504888 219218
rect 504568 218898 504610 219134
rect 504846 218898 504888 219134
rect 504568 218866 504888 218898
rect 514808 219454 515128 219486
rect 514808 219218 514850 219454
rect 515086 219218 515128 219454
rect 514808 219134 515128 219218
rect 514808 218898 514850 219134
rect 515086 218898 515128 219134
rect 514808 218866 515128 218898
rect 525048 219454 525368 219486
rect 525048 219218 525090 219454
rect 525326 219218 525368 219454
rect 525048 219134 525368 219218
rect 525048 218898 525090 219134
rect 525326 218898 525368 219134
rect 525048 218866 525368 218898
rect 535288 219454 535608 219486
rect 535288 219218 535330 219454
rect 535566 219218 535608 219454
rect 535288 219134 535608 219218
rect 535288 218898 535330 219134
rect 535566 218898 535608 219134
rect 535288 218866 535608 218898
rect 28408 201454 28728 201486
rect 28408 201218 28450 201454
rect 28686 201218 28728 201454
rect 28408 201134 28728 201218
rect 28408 200898 28450 201134
rect 28686 200898 28728 201134
rect 28408 200866 28728 200898
rect 38648 201454 38968 201486
rect 38648 201218 38690 201454
rect 38926 201218 38968 201454
rect 38648 201134 38968 201218
rect 38648 200898 38690 201134
rect 38926 200898 38968 201134
rect 38648 200866 38968 200898
rect 48888 201454 49208 201486
rect 48888 201218 48930 201454
rect 49166 201218 49208 201454
rect 48888 201134 49208 201218
rect 48888 200898 48930 201134
rect 49166 200898 49208 201134
rect 48888 200866 49208 200898
rect 59128 201454 59448 201486
rect 59128 201218 59170 201454
rect 59406 201218 59448 201454
rect 59128 201134 59448 201218
rect 59128 200898 59170 201134
rect 59406 200898 59448 201134
rect 59128 200866 59448 200898
rect 69368 201454 69688 201486
rect 69368 201218 69410 201454
rect 69646 201218 69688 201454
rect 69368 201134 69688 201218
rect 69368 200898 69410 201134
rect 69646 200898 69688 201134
rect 69368 200866 69688 200898
rect 79608 201454 79928 201486
rect 79608 201218 79650 201454
rect 79886 201218 79928 201454
rect 79608 201134 79928 201218
rect 79608 200898 79650 201134
rect 79886 200898 79928 201134
rect 79608 200866 79928 200898
rect 89848 201454 90168 201486
rect 89848 201218 89890 201454
rect 90126 201218 90168 201454
rect 89848 201134 90168 201218
rect 89848 200898 89890 201134
rect 90126 200898 90168 201134
rect 89848 200866 90168 200898
rect 100088 201454 100408 201486
rect 100088 201218 100130 201454
rect 100366 201218 100408 201454
rect 100088 201134 100408 201218
rect 100088 200898 100130 201134
rect 100366 200898 100408 201134
rect 100088 200866 100408 200898
rect 110328 201454 110648 201486
rect 110328 201218 110370 201454
rect 110606 201218 110648 201454
rect 110328 201134 110648 201218
rect 110328 200898 110370 201134
rect 110606 200898 110648 201134
rect 110328 200866 110648 200898
rect 120568 201454 120888 201486
rect 120568 201218 120610 201454
rect 120846 201218 120888 201454
rect 120568 201134 120888 201218
rect 120568 200898 120610 201134
rect 120846 200898 120888 201134
rect 120568 200866 120888 200898
rect 130808 201454 131128 201486
rect 130808 201218 130850 201454
rect 131086 201218 131128 201454
rect 130808 201134 131128 201218
rect 130808 200898 130850 201134
rect 131086 200898 131128 201134
rect 130808 200866 131128 200898
rect 141048 201454 141368 201486
rect 141048 201218 141090 201454
rect 141326 201218 141368 201454
rect 141048 201134 141368 201218
rect 141048 200898 141090 201134
rect 141326 200898 141368 201134
rect 141048 200866 141368 200898
rect 151288 201454 151608 201486
rect 151288 201218 151330 201454
rect 151566 201218 151608 201454
rect 151288 201134 151608 201218
rect 151288 200898 151330 201134
rect 151566 200898 151608 201134
rect 151288 200866 151608 200898
rect 161528 201454 161848 201486
rect 161528 201218 161570 201454
rect 161806 201218 161848 201454
rect 161528 201134 161848 201218
rect 161528 200898 161570 201134
rect 161806 200898 161848 201134
rect 161528 200866 161848 200898
rect 171768 201454 172088 201486
rect 171768 201218 171810 201454
rect 172046 201218 172088 201454
rect 171768 201134 172088 201218
rect 171768 200898 171810 201134
rect 172046 200898 172088 201134
rect 171768 200866 172088 200898
rect 182008 201454 182328 201486
rect 182008 201218 182050 201454
rect 182286 201218 182328 201454
rect 182008 201134 182328 201218
rect 182008 200898 182050 201134
rect 182286 200898 182328 201134
rect 182008 200866 182328 200898
rect 192248 201454 192568 201486
rect 192248 201218 192290 201454
rect 192526 201218 192568 201454
rect 192248 201134 192568 201218
rect 192248 200898 192290 201134
rect 192526 200898 192568 201134
rect 192248 200866 192568 200898
rect 202488 201454 202808 201486
rect 202488 201218 202530 201454
rect 202766 201218 202808 201454
rect 202488 201134 202808 201218
rect 202488 200898 202530 201134
rect 202766 200898 202808 201134
rect 202488 200866 202808 200898
rect 212728 201454 213048 201486
rect 212728 201218 212770 201454
rect 213006 201218 213048 201454
rect 212728 201134 213048 201218
rect 212728 200898 212770 201134
rect 213006 200898 213048 201134
rect 212728 200866 213048 200898
rect 222968 201454 223288 201486
rect 222968 201218 223010 201454
rect 223246 201218 223288 201454
rect 222968 201134 223288 201218
rect 222968 200898 223010 201134
rect 223246 200898 223288 201134
rect 222968 200866 223288 200898
rect 233208 201454 233528 201486
rect 233208 201218 233250 201454
rect 233486 201218 233528 201454
rect 233208 201134 233528 201218
rect 233208 200898 233250 201134
rect 233486 200898 233528 201134
rect 233208 200866 233528 200898
rect 243448 201454 243768 201486
rect 243448 201218 243490 201454
rect 243726 201218 243768 201454
rect 243448 201134 243768 201218
rect 243448 200898 243490 201134
rect 243726 200898 243768 201134
rect 243448 200866 243768 200898
rect 253688 201454 254008 201486
rect 253688 201218 253730 201454
rect 253966 201218 254008 201454
rect 253688 201134 254008 201218
rect 253688 200898 253730 201134
rect 253966 200898 254008 201134
rect 253688 200866 254008 200898
rect 263928 201454 264248 201486
rect 263928 201218 263970 201454
rect 264206 201218 264248 201454
rect 263928 201134 264248 201218
rect 263928 200898 263970 201134
rect 264206 200898 264248 201134
rect 263928 200866 264248 200898
rect 274168 201454 274488 201486
rect 274168 201218 274210 201454
rect 274446 201218 274488 201454
rect 274168 201134 274488 201218
rect 274168 200898 274210 201134
rect 274446 200898 274488 201134
rect 274168 200866 274488 200898
rect 284408 201454 284728 201486
rect 284408 201218 284450 201454
rect 284686 201218 284728 201454
rect 284408 201134 284728 201218
rect 284408 200898 284450 201134
rect 284686 200898 284728 201134
rect 284408 200866 284728 200898
rect 294648 201454 294968 201486
rect 294648 201218 294690 201454
rect 294926 201218 294968 201454
rect 294648 201134 294968 201218
rect 294648 200898 294690 201134
rect 294926 200898 294968 201134
rect 294648 200866 294968 200898
rect 304888 201454 305208 201486
rect 304888 201218 304930 201454
rect 305166 201218 305208 201454
rect 304888 201134 305208 201218
rect 304888 200898 304930 201134
rect 305166 200898 305208 201134
rect 304888 200866 305208 200898
rect 315128 201454 315448 201486
rect 315128 201218 315170 201454
rect 315406 201218 315448 201454
rect 315128 201134 315448 201218
rect 315128 200898 315170 201134
rect 315406 200898 315448 201134
rect 315128 200866 315448 200898
rect 325368 201454 325688 201486
rect 325368 201218 325410 201454
rect 325646 201218 325688 201454
rect 325368 201134 325688 201218
rect 325368 200898 325410 201134
rect 325646 200898 325688 201134
rect 325368 200866 325688 200898
rect 335608 201454 335928 201486
rect 335608 201218 335650 201454
rect 335886 201218 335928 201454
rect 335608 201134 335928 201218
rect 335608 200898 335650 201134
rect 335886 200898 335928 201134
rect 335608 200866 335928 200898
rect 345848 201454 346168 201486
rect 345848 201218 345890 201454
rect 346126 201218 346168 201454
rect 345848 201134 346168 201218
rect 345848 200898 345890 201134
rect 346126 200898 346168 201134
rect 345848 200866 346168 200898
rect 356088 201454 356408 201486
rect 356088 201218 356130 201454
rect 356366 201218 356408 201454
rect 356088 201134 356408 201218
rect 356088 200898 356130 201134
rect 356366 200898 356408 201134
rect 356088 200866 356408 200898
rect 366328 201454 366648 201486
rect 366328 201218 366370 201454
rect 366606 201218 366648 201454
rect 366328 201134 366648 201218
rect 366328 200898 366370 201134
rect 366606 200898 366648 201134
rect 366328 200866 366648 200898
rect 376568 201454 376888 201486
rect 376568 201218 376610 201454
rect 376846 201218 376888 201454
rect 376568 201134 376888 201218
rect 376568 200898 376610 201134
rect 376846 200898 376888 201134
rect 376568 200866 376888 200898
rect 386808 201454 387128 201486
rect 386808 201218 386850 201454
rect 387086 201218 387128 201454
rect 386808 201134 387128 201218
rect 386808 200898 386850 201134
rect 387086 200898 387128 201134
rect 386808 200866 387128 200898
rect 397048 201454 397368 201486
rect 397048 201218 397090 201454
rect 397326 201218 397368 201454
rect 397048 201134 397368 201218
rect 397048 200898 397090 201134
rect 397326 200898 397368 201134
rect 397048 200866 397368 200898
rect 407288 201454 407608 201486
rect 407288 201218 407330 201454
rect 407566 201218 407608 201454
rect 407288 201134 407608 201218
rect 407288 200898 407330 201134
rect 407566 200898 407608 201134
rect 407288 200866 407608 200898
rect 417528 201454 417848 201486
rect 417528 201218 417570 201454
rect 417806 201218 417848 201454
rect 417528 201134 417848 201218
rect 417528 200898 417570 201134
rect 417806 200898 417848 201134
rect 417528 200866 417848 200898
rect 427768 201454 428088 201486
rect 427768 201218 427810 201454
rect 428046 201218 428088 201454
rect 427768 201134 428088 201218
rect 427768 200898 427810 201134
rect 428046 200898 428088 201134
rect 427768 200866 428088 200898
rect 438008 201454 438328 201486
rect 438008 201218 438050 201454
rect 438286 201218 438328 201454
rect 438008 201134 438328 201218
rect 438008 200898 438050 201134
rect 438286 200898 438328 201134
rect 438008 200866 438328 200898
rect 448248 201454 448568 201486
rect 448248 201218 448290 201454
rect 448526 201218 448568 201454
rect 448248 201134 448568 201218
rect 448248 200898 448290 201134
rect 448526 200898 448568 201134
rect 448248 200866 448568 200898
rect 458488 201454 458808 201486
rect 458488 201218 458530 201454
rect 458766 201218 458808 201454
rect 458488 201134 458808 201218
rect 458488 200898 458530 201134
rect 458766 200898 458808 201134
rect 458488 200866 458808 200898
rect 468728 201454 469048 201486
rect 468728 201218 468770 201454
rect 469006 201218 469048 201454
rect 468728 201134 469048 201218
rect 468728 200898 468770 201134
rect 469006 200898 469048 201134
rect 468728 200866 469048 200898
rect 478968 201454 479288 201486
rect 478968 201218 479010 201454
rect 479246 201218 479288 201454
rect 478968 201134 479288 201218
rect 478968 200898 479010 201134
rect 479246 200898 479288 201134
rect 478968 200866 479288 200898
rect 489208 201454 489528 201486
rect 489208 201218 489250 201454
rect 489486 201218 489528 201454
rect 489208 201134 489528 201218
rect 489208 200898 489250 201134
rect 489486 200898 489528 201134
rect 489208 200866 489528 200898
rect 499448 201454 499768 201486
rect 499448 201218 499490 201454
rect 499726 201218 499768 201454
rect 499448 201134 499768 201218
rect 499448 200898 499490 201134
rect 499726 200898 499768 201134
rect 499448 200866 499768 200898
rect 509688 201454 510008 201486
rect 509688 201218 509730 201454
rect 509966 201218 510008 201454
rect 509688 201134 510008 201218
rect 509688 200898 509730 201134
rect 509966 200898 510008 201134
rect 509688 200866 510008 200898
rect 519928 201454 520248 201486
rect 519928 201218 519970 201454
rect 520206 201218 520248 201454
rect 519928 201134 520248 201218
rect 519928 200898 519970 201134
rect 520206 200898 520248 201134
rect 519928 200866 520248 200898
rect 530168 201454 530488 201486
rect 530168 201218 530210 201454
rect 530446 201218 530488 201454
rect 530168 201134 530488 201218
rect 530168 200898 530210 201134
rect 530446 200898 530488 201134
rect 530168 200866 530488 200898
rect 15754 186938 15786 187174
rect 16022 186938 16106 187174
rect 16342 186938 16374 187174
rect 15754 186854 16374 186938
rect 15754 186618 15786 186854
rect 16022 186618 16106 186854
rect 16342 186618 16374 186854
rect 15754 151174 16374 186618
rect 541714 190894 542334 226338
rect 541714 190658 541746 190894
rect 541982 190658 542066 190894
rect 542302 190658 542334 190894
rect 541714 190574 542334 190658
rect 541714 190338 541746 190574
rect 541982 190338 542066 190574
rect 542302 190338 542334 190574
rect 23288 183454 23608 183486
rect 23288 183218 23330 183454
rect 23566 183218 23608 183454
rect 23288 183134 23608 183218
rect 23288 182898 23330 183134
rect 23566 182898 23608 183134
rect 23288 182866 23608 182898
rect 33528 183454 33848 183486
rect 33528 183218 33570 183454
rect 33806 183218 33848 183454
rect 33528 183134 33848 183218
rect 33528 182898 33570 183134
rect 33806 182898 33848 183134
rect 33528 182866 33848 182898
rect 43768 183454 44088 183486
rect 43768 183218 43810 183454
rect 44046 183218 44088 183454
rect 43768 183134 44088 183218
rect 43768 182898 43810 183134
rect 44046 182898 44088 183134
rect 43768 182866 44088 182898
rect 54008 183454 54328 183486
rect 54008 183218 54050 183454
rect 54286 183218 54328 183454
rect 54008 183134 54328 183218
rect 54008 182898 54050 183134
rect 54286 182898 54328 183134
rect 54008 182866 54328 182898
rect 64248 183454 64568 183486
rect 64248 183218 64290 183454
rect 64526 183218 64568 183454
rect 64248 183134 64568 183218
rect 64248 182898 64290 183134
rect 64526 182898 64568 183134
rect 64248 182866 64568 182898
rect 74488 183454 74808 183486
rect 74488 183218 74530 183454
rect 74766 183218 74808 183454
rect 74488 183134 74808 183218
rect 74488 182898 74530 183134
rect 74766 182898 74808 183134
rect 74488 182866 74808 182898
rect 84728 183454 85048 183486
rect 84728 183218 84770 183454
rect 85006 183218 85048 183454
rect 84728 183134 85048 183218
rect 84728 182898 84770 183134
rect 85006 182898 85048 183134
rect 84728 182866 85048 182898
rect 94968 183454 95288 183486
rect 94968 183218 95010 183454
rect 95246 183218 95288 183454
rect 94968 183134 95288 183218
rect 94968 182898 95010 183134
rect 95246 182898 95288 183134
rect 94968 182866 95288 182898
rect 105208 183454 105528 183486
rect 105208 183218 105250 183454
rect 105486 183218 105528 183454
rect 105208 183134 105528 183218
rect 105208 182898 105250 183134
rect 105486 182898 105528 183134
rect 105208 182866 105528 182898
rect 115448 183454 115768 183486
rect 115448 183218 115490 183454
rect 115726 183218 115768 183454
rect 115448 183134 115768 183218
rect 115448 182898 115490 183134
rect 115726 182898 115768 183134
rect 115448 182866 115768 182898
rect 125688 183454 126008 183486
rect 125688 183218 125730 183454
rect 125966 183218 126008 183454
rect 125688 183134 126008 183218
rect 125688 182898 125730 183134
rect 125966 182898 126008 183134
rect 125688 182866 126008 182898
rect 135928 183454 136248 183486
rect 135928 183218 135970 183454
rect 136206 183218 136248 183454
rect 135928 183134 136248 183218
rect 135928 182898 135970 183134
rect 136206 182898 136248 183134
rect 135928 182866 136248 182898
rect 146168 183454 146488 183486
rect 146168 183218 146210 183454
rect 146446 183218 146488 183454
rect 146168 183134 146488 183218
rect 146168 182898 146210 183134
rect 146446 182898 146488 183134
rect 146168 182866 146488 182898
rect 156408 183454 156728 183486
rect 156408 183218 156450 183454
rect 156686 183218 156728 183454
rect 156408 183134 156728 183218
rect 156408 182898 156450 183134
rect 156686 182898 156728 183134
rect 156408 182866 156728 182898
rect 166648 183454 166968 183486
rect 166648 183218 166690 183454
rect 166926 183218 166968 183454
rect 166648 183134 166968 183218
rect 166648 182898 166690 183134
rect 166926 182898 166968 183134
rect 166648 182866 166968 182898
rect 176888 183454 177208 183486
rect 176888 183218 176930 183454
rect 177166 183218 177208 183454
rect 176888 183134 177208 183218
rect 176888 182898 176930 183134
rect 177166 182898 177208 183134
rect 176888 182866 177208 182898
rect 187128 183454 187448 183486
rect 187128 183218 187170 183454
rect 187406 183218 187448 183454
rect 187128 183134 187448 183218
rect 187128 182898 187170 183134
rect 187406 182898 187448 183134
rect 187128 182866 187448 182898
rect 197368 183454 197688 183486
rect 197368 183218 197410 183454
rect 197646 183218 197688 183454
rect 197368 183134 197688 183218
rect 197368 182898 197410 183134
rect 197646 182898 197688 183134
rect 197368 182866 197688 182898
rect 207608 183454 207928 183486
rect 207608 183218 207650 183454
rect 207886 183218 207928 183454
rect 207608 183134 207928 183218
rect 207608 182898 207650 183134
rect 207886 182898 207928 183134
rect 207608 182866 207928 182898
rect 217848 183454 218168 183486
rect 217848 183218 217890 183454
rect 218126 183218 218168 183454
rect 217848 183134 218168 183218
rect 217848 182898 217890 183134
rect 218126 182898 218168 183134
rect 217848 182866 218168 182898
rect 228088 183454 228408 183486
rect 228088 183218 228130 183454
rect 228366 183218 228408 183454
rect 228088 183134 228408 183218
rect 228088 182898 228130 183134
rect 228366 182898 228408 183134
rect 228088 182866 228408 182898
rect 238328 183454 238648 183486
rect 238328 183218 238370 183454
rect 238606 183218 238648 183454
rect 238328 183134 238648 183218
rect 238328 182898 238370 183134
rect 238606 182898 238648 183134
rect 238328 182866 238648 182898
rect 248568 183454 248888 183486
rect 248568 183218 248610 183454
rect 248846 183218 248888 183454
rect 248568 183134 248888 183218
rect 248568 182898 248610 183134
rect 248846 182898 248888 183134
rect 248568 182866 248888 182898
rect 258808 183454 259128 183486
rect 258808 183218 258850 183454
rect 259086 183218 259128 183454
rect 258808 183134 259128 183218
rect 258808 182898 258850 183134
rect 259086 182898 259128 183134
rect 258808 182866 259128 182898
rect 269048 183454 269368 183486
rect 269048 183218 269090 183454
rect 269326 183218 269368 183454
rect 269048 183134 269368 183218
rect 269048 182898 269090 183134
rect 269326 182898 269368 183134
rect 269048 182866 269368 182898
rect 279288 183454 279608 183486
rect 279288 183218 279330 183454
rect 279566 183218 279608 183454
rect 279288 183134 279608 183218
rect 279288 182898 279330 183134
rect 279566 182898 279608 183134
rect 279288 182866 279608 182898
rect 289528 183454 289848 183486
rect 289528 183218 289570 183454
rect 289806 183218 289848 183454
rect 289528 183134 289848 183218
rect 289528 182898 289570 183134
rect 289806 182898 289848 183134
rect 289528 182866 289848 182898
rect 299768 183454 300088 183486
rect 299768 183218 299810 183454
rect 300046 183218 300088 183454
rect 299768 183134 300088 183218
rect 299768 182898 299810 183134
rect 300046 182898 300088 183134
rect 299768 182866 300088 182898
rect 310008 183454 310328 183486
rect 310008 183218 310050 183454
rect 310286 183218 310328 183454
rect 310008 183134 310328 183218
rect 310008 182898 310050 183134
rect 310286 182898 310328 183134
rect 310008 182866 310328 182898
rect 320248 183454 320568 183486
rect 320248 183218 320290 183454
rect 320526 183218 320568 183454
rect 320248 183134 320568 183218
rect 320248 182898 320290 183134
rect 320526 182898 320568 183134
rect 320248 182866 320568 182898
rect 330488 183454 330808 183486
rect 330488 183218 330530 183454
rect 330766 183218 330808 183454
rect 330488 183134 330808 183218
rect 330488 182898 330530 183134
rect 330766 182898 330808 183134
rect 330488 182866 330808 182898
rect 340728 183454 341048 183486
rect 340728 183218 340770 183454
rect 341006 183218 341048 183454
rect 340728 183134 341048 183218
rect 340728 182898 340770 183134
rect 341006 182898 341048 183134
rect 340728 182866 341048 182898
rect 350968 183454 351288 183486
rect 350968 183218 351010 183454
rect 351246 183218 351288 183454
rect 350968 183134 351288 183218
rect 350968 182898 351010 183134
rect 351246 182898 351288 183134
rect 350968 182866 351288 182898
rect 361208 183454 361528 183486
rect 361208 183218 361250 183454
rect 361486 183218 361528 183454
rect 361208 183134 361528 183218
rect 361208 182898 361250 183134
rect 361486 182898 361528 183134
rect 361208 182866 361528 182898
rect 371448 183454 371768 183486
rect 371448 183218 371490 183454
rect 371726 183218 371768 183454
rect 371448 183134 371768 183218
rect 371448 182898 371490 183134
rect 371726 182898 371768 183134
rect 371448 182866 371768 182898
rect 381688 183454 382008 183486
rect 381688 183218 381730 183454
rect 381966 183218 382008 183454
rect 381688 183134 382008 183218
rect 381688 182898 381730 183134
rect 381966 182898 382008 183134
rect 381688 182866 382008 182898
rect 391928 183454 392248 183486
rect 391928 183218 391970 183454
rect 392206 183218 392248 183454
rect 391928 183134 392248 183218
rect 391928 182898 391970 183134
rect 392206 182898 392248 183134
rect 391928 182866 392248 182898
rect 402168 183454 402488 183486
rect 402168 183218 402210 183454
rect 402446 183218 402488 183454
rect 402168 183134 402488 183218
rect 402168 182898 402210 183134
rect 402446 182898 402488 183134
rect 402168 182866 402488 182898
rect 412408 183454 412728 183486
rect 412408 183218 412450 183454
rect 412686 183218 412728 183454
rect 412408 183134 412728 183218
rect 412408 182898 412450 183134
rect 412686 182898 412728 183134
rect 412408 182866 412728 182898
rect 422648 183454 422968 183486
rect 422648 183218 422690 183454
rect 422926 183218 422968 183454
rect 422648 183134 422968 183218
rect 422648 182898 422690 183134
rect 422926 182898 422968 183134
rect 422648 182866 422968 182898
rect 432888 183454 433208 183486
rect 432888 183218 432930 183454
rect 433166 183218 433208 183454
rect 432888 183134 433208 183218
rect 432888 182898 432930 183134
rect 433166 182898 433208 183134
rect 432888 182866 433208 182898
rect 443128 183454 443448 183486
rect 443128 183218 443170 183454
rect 443406 183218 443448 183454
rect 443128 183134 443448 183218
rect 443128 182898 443170 183134
rect 443406 182898 443448 183134
rect 443128 182866 443448 182898
rect 453368 183454 453688 183486
rect 453368 183218 453410 183454
rect 453646 183218 453688 183454
rect 453368 183134 453688 183218
rect 453368 182898 453410 183134
rect 453646 182898 453688 183134
rect 453368 182866 453688 182898
rect 463608 183454 463928 183486
rect 463608 183218 463650 183454
rect 463886 183218 463928 183454
rect 463608 183134 463928 183218
rect 463608 182898 463650 183134
rect 463886 182898 463928 183134
rect 463608 182866 463928 182898
rect 473848 183454 474168 183486
rect 473848 183218 473890 183454
rect 474126 183218 474168 183454
rect 473848 183134 474168 183218
rect 473848 182898 473890 183134
rect 474126 182898 474168 183134
rect 473848 182866 474168 182898
rect 484088 183454 484408 183486
rect 484088 183218 484130 183454
rect 484366 183218 484408 183454
rect 484088 183134 484408 183218
rect 484088 182898 484130 183134
rect 484366 182898 484408 183134
rect 484088 182866 484408 182898
rect 494328 183454 494648 183486
rect 494328 183218 494370 183454
rect 494606 183218 494648 183454
rect 494328 183134 494648 183218
rect 494328 182898 494370 183134
rect 494606 182898 494648 183134
rect 494328 182866 494648 182898
rect 504568 183454 504888 183486
rect 504568 183218 504610 183454
rect 504846 183218 504888 183454
rect 504568 183134 504888 183218
rect 504568 182898 504610 183134
rect 504846 182898 504888 183134
rect 504568 182866 504888 182898
rect 514808 183454 515128 183486
rect 514808 183218 514850 183454
rect 515086 183218 515128 183454
rect 514808 183134 515128 183218
rect 514808 182898 514850 183134
rect 515086 182898 515128 183134
rect 514808 182866 515128 182898
rect 525048 183454 525368 183486
rect 525048 183218 525090 183454
rect 525326 183218 525368 183454
rect 525048 183134 525368 183218
rect 525048 182898 525090 183134
rect 525326 182898 525368 183134
rect 525048 182866 525368 182898
rect 535288 183454 535608 183486
rect 535288 183218 535330 183454
rect 535566 183218 535608 183454
rect 535288 183134 535608 183218
rect 535288 182898 535330 183134
rect 535566 182898 535608 183134
rect 535288 182866 535608 182898
rect 28408 165454 28728 165486
rect 28408 165218 28450 165454
rect 28686 165218 28728 165454
rect 28408 165134 28728 165218
rect 28408 164898 28450 165134
rect 28686 164898 28728 165134
rect 28408 164866 28728 164898
rect 38648 165454 38968 165486
rect 38648 165218 38690 165454
rect 38926 165218 38968 165454
rect 38648 165134 38968 165218
rect 38648 164898 38690 165134
rect 38926 164898 38968 165134
rect 38648 164866 38968 164898
rect 48888 165454 49208 165486
rect 48888 165218 48930 165454
rect 49166 165218 49208 165454
rect 48888 165134 49208 165218
rect 48888 164898 48930 165134
rect 49166 164898 49208 165134
rect 48888 164866 49208 164898
rect 59128 165454 59448 165486
rect 59128 165218 59170 165454
rect 59406 165218 59448 165454
rect 59128 165134 59448 165218
rect 59128 164898 59170 165134
rect 59406 164898 59448 165134
rect 59128 164866 59448 164898
rect 69368 165454 69688 165486
rect 69368 165218 69410 165454
rect 69646 165218 69688 165454
rect 69368 165134 69688 165218
rect 69368 164898 69410 165134
rect 69646 164898 69688 165134
rect 69368 164866 69688 164898
rect 79608 165454 79928 165486
rect 79608 165218 79650 165454
rect 79886 165218 79928 165454
rect 79608 165134 79928 165218
rect 79608 164898 79650 165134
rect 79886 164898 79928 165134
rect 79608 164866 79928 164898
rect 89848 165454 90168 165486
rect 89848 165218 89890 165454
rect 90126 165218 90168 165454
rect 89848 165134 90168 165218
rect 89848 164898 89890 165134
rect 90126 164898 90168 165134
rect 89848 164866 90168 164898
rect 100088 165454 100408 165486
rect 100088 165218 100130 165454
rect 100366 165218 100408 165454
rect 100088 165134 100408 165218
rect 100088 164898 100130 165134
rect 100366 164898 100408 165134
rect 100088 164866 100408 164898
rect 110328 165454 110648 165486
rect 110328 165218 110370 165454
rect 110606 165218 110648 165454
rect 110328 165134 110648 165218
rect 110328 164898 110370 165134
rect 110606 164898 110648 165134
rect 110328 164866 110648 164898
rect 120568 165454 120888 165486
rect 120568 165218 120610 165454
rect 120846 165218 120888 165454
rect 120568 165134 120888 165218
rect 120568 164898 120610 165134
rect 120846 164898 120888 165134
rect 120568 164866 120888 164898
rect 130808 165454 131128 165486
rect 130808 165218 130850 165454
rect 131086 165218 131128 165454
rect 130808 165134 131128 165218
rect 130808 164898 130850 165134
rect 131086 164898 131128 165134
rect 130808 164866 131128 164898
rect 141048 165454 141368 165486
rect 141048 165218 141090 165454
rect 141326 165218 141368 165454
rect 141048 165134 141368 165218
rect 141048 164898 141090 165134
rect 141326 164898 141368 165134
rect 141048 164866 141368 164898
rect 151288 165454 151608 165486
rect 151288 165218 151330 165454
rect 151566 165218 151608 165454
rect 151288 165134 151608 165218
rect 151288 164898 151330 165134
rect 151566 164898 151608 165134
rect 151288 164866 151608 164898
rect 161528 165454 161848 165486
rect 161528 165218 161570 165454
rect 161806 165218 161848 165454
rect 161528 165134 161848 165218
rect 161528 164898 161570 165134
rect 161806 164898 161848 165134
rect 161528 164866 161848 164898
rect 171768 165454 172088 165486
rect 171768 165218 171810 165454
rect 172046 165218 172088 165454
rect 171768 165134 172088 165218
rect 171768 164898 171810 165134
rect 172046 164898 172088 165134
rect 171768 164866 172088 164898
rect 182008 165454 182328 165486
rect 182008 165218 182050 165454
rect 182286 165218 182328 165454
rect 182008 165134 182328 165218
rect 182008 164898 182050 165134
rect 182286 164898 182328 165134
rect 182008 164866 182328 164898
rect 192248 165454 192568 165486
rect 192248 165218 192290 165454
rect 192526 165218 192568 165454
rect 192248 165134 192568 165218
rect 192248 164898 192290 165134
rect 192526 164898 192568 165134
rect 192248 164866 192568 164898
rect 202488 165454 202808 165486
rect 202488 165218 202530 165454
rect 202766 165218 202808 165454
rect 202488 165134 202808 165218
rect 202488 164898 202530 165134
rect 202766 164898 202808 165134
rect 202488 164866 202808 164898
rect 212728 165454 213048 165486
rect 212728 165218 212770 165454
rect 213006 165218 213048 165454
rect 212728 165134 213048 165218
rect 212728 164898 212770 165134
rect 213006 164898 213048 165134
rect 212728 164866 213048 164898
rect 222968 165454 223288 165486
rect 222968 165218 223010 165454
rect 223246 165218 223288 165454
rect 222968 165134 223288 165218
rect 222968 164898 223010 165134
rect 223246 164898 223288 165134
rect 222968 164866 223288 164898
rect 233208 165454 233528 165486
rect 233208 165218 233250 165454
rect 233486 165218 233528 165454
rect 233208 165134 233528 165218
rect 233208 164898 233250 165134
rect 233486 164898 233528 165134
rect 233208 164866 233528 164898
rect 243448 165454 243768 165486
rect 243448 165218 243490 165454
rect 243726 165218 243768 165454
rect 243448 165134 243768 165218
rect 243448 164898 243490 165134
rect 243726 164898 243768 165134
rect 243448 164866 243768 164898
rect 253688 165454 254008 165486
rect 253688 165218 253730 165454
rect 253966 165218 254008 165454
rect 253688 165134 254008 165218
rect 253688 164898 253730 165134
rect 253966 164898 254008 165134
rect 253688 164866 254008 164898
rect 263928 165454 264248 165486
rect 263928 165218 263970 165454
rect 264206 165218 264248 165454
rect 263928 165134 264248 165218
rect 263928 164898 263970 165134
rect 264206 164898 264248 165134
rect 263928 164866 264248 164898
rect 274168 165454 274488 165486
rect 274168 165218 274210 165454
rect 274446 165218 274488 165454
rect 274168 165134 274488 165218
rect 274168 164898 274210 165134
rect 274446 164898 274488 165134
rect 274168 164866 274488 164898
rect 284408 165454 284728 165486
rect 284408 165218 284450 165454
rect 284686 165218 284728 165454
rect 284408 165134 284728 165218
rect 284408 164898 284450 165134
rect 284686 164898 284728 165134
rect 284408 164866 284728 164898
rect 294648 165454 294968 165486
rect 294648 165218 294690 165454
rect 294926 165218 294968 165454
rect 294648 165134 294968 165218
rect 294648 164898 294690 165134
rect 294926 164898 294968 165134
rect 294648 164866 294968 164898
rect 304888 165454 305208 165486
rect 304888 165218 304930 165454
rect 305166 165218 305208 165454
rect 304888 165134 305208 165218
rect 304888 164898 304930 165134
rect 305166 164898 305208 165134
rect 304888 164866 305208 164898
rect 315128 165454 315448 165486
rect 315128 165218 315170 165454
rect 315406 165218 315448 165454
rect 315128 165134 315448 165218
rect 315128 164898 315170 165134
rect 315406 164898 315448 165134
rect 315128 164866 315448 164898
rect 325368 165454 325688 165486
rect 325368 165218 325410 165454
rect 325646 165218 325688 165454
rect 325368 165134 325688 165218
rect 325368 164898 325410 165134
rect 325646 164898 325688 165134
rect 325368 164866 325688 164898
rect 335608 165454 335928 165486
rect 335608 165218 335650 165454
rect 335886 165218 335928 165454
rect 335608 165134 335928 165218
rect 335608 164898 335650 165134
rect 335886 164898 335928 165134
rect 335608 164866 335928 164898
rect 345848 165454 346168 165486
rect 345848 165218 345890 165454
rect 346126 165218 346168 165454
rect 345848 165134 346168 165218
rect 345848 164898 345890 165134
rect 346126 164898 346168 165134
rect 345848 164866 346168 164898
rect 356088 165454 356408 165486
rect 356088 165218 356130 165454
rect 356366 165218 356408 165454
rect 356088 165134 356408 165218
rect 356088 164898 356130 165134
rect 356366 164898 356408 165134
rect 356088 164866 356408 164898
rect 366328 165454 366648 165486
rect 366328 165218 366370 165454
rect 366606 165218 366648 165454
rect 366328 165134 366648 165218
rect 366328 164898 366370 165134
rect 366606 164898 366648 165134
rect 366328 164866 366648 164898
rect 376568 165454 376888 165486
rect 376568 165218 376610 165454
rect 376846 165218 376888 165454
rect 376568 165134 376888 165218
rect 376568 164898 376610 165134
rect 376846 164898 376888 165134
rect 376568 164866 376888 164898
rect 386808 165454 387128 165486
rect 386808 165218 386850 165454
rect 387086 165218 387128 165454
rect 386808 165134 387128 165218
rect 386808 164898 386850 165134
rect 387086 164898 387128 165134
rect 386808 164866 387128 164898
rect 397048 165454 397368 165486
rect 397048 165218 397090 165454
rect 397326 165218 397368 165454
rect 397048 165134 397368 165218
rect 397048 164898 397090 165134
rect 397326 164898 397368 165134
rect 397048 164866 397368 164898
rect 407288 165454 407608 165486
rect 407288 165218 407330 165454
rect 407566 165218 407608 165454
rect 407288 165134 407608 165218
rect 407288 164898 407330 165134
rect 407566 164898 407608 165134
rect 407288 164866 407608 164898
rect 417528 165454 417848 165486
rect 417528 165218 417570 165454
rect 417806 165218 417848 165454
rect 417528 165134 417848 165218
rect 417528 164898 417570 165134
rect 417806 164898 417848 165134
rect 417528 164866 417848 164898
rect 427768 165454 428088 165486
rect 427768 165218 427810 165454
rect 428046 165218 428088 165454
rect 427768 165134 428088 165218
rect 427768 164898 427810 165134
rect 428046 164898 428088 165134
rect 427768 164866 428088 164898
rect 438008 165454 438328 165486
rect 438008 165218 438050 165454
rect 438286 165218 438328 165454
rect 438008 165134 438328 165218
rect 438008 164898 438050 165134
rect 438286 164898 438328 165134
rect 438008 164866 438328 164898
rect 448248 165454 448568 165486
rect 448248 165218 448290 165454
rect 448526 165218 448568 165454
rect 448248 165134 448568 165218
rect 448248 164898 448290 165134
rect 448526 164898 448568 165134
rect 448248 164866 448568 164898
rect 458488 165454 458808 165486
rect 458488 165218 458530 165454
rect 458766 165218 458808 165454
rect 458488 165134 458808 165218
rect 458488 164898 458530 165134
rect 458766 164898 458808 165134
rect 458488 164866 458808 164898
rect 468728 165454 469048 165486
rect 468728 165218 468770 165454
rect 469006 165218 469048 165454
rect 468728 165134 469048 165218
rect 468728 164898 468770 165134
rect 469006 164898 469048 165134
rect 468728 164866 469048 164898
rect 478968 165454 479288 165486
rect 478968 165218 479010 165454
rect 479246 165218 479288 165454
rect 478968 165134 479288 165218
rect 478968 164898 479010 165134
rect 479246 164898 479288 165134
rect 478968 164866 479288 164898
rect 489208 165454 489528 165486
rect 489208 165218 489250 165454
rect 489486 165218 489528 165454
rect 489208 165134 489528 165218
rect 489208 164898 489250 165134
rect 489486 164898 489528 165134
rect 489208 164866 489528 164898
rect 499448 165454 499768 165486
rect 499448 165218 499490 165454
rect 499726 165218 499768 165454
rect 499448 165134 499768 165218
rect 499448 164898 499490 165134
rect 499726 164898 499768 165134
rect 499448 164866 499768 164898
rect 509688 165454 510008 165486
rect 509688 165218 509730 165454
rect 509966 165218 510008 165454
rect 509688 165134 510008 165218
rect 509688 164898 509730 165134
rect 509966 164898 510008 165134
rect 509688 164866 510008 164898
rect 519928 165454 520248 165486
rect 519928 165218 519970 165454
rect 520206 165218 520248 165454
rect 519928 165134 520248 165218
rect 519928 164898 519970 165134
rect 520206 164898 520248 165134
rect 519928 164866 520248 164898
rect 530168 165454 530488 165486
rect 530168 165218 530210 165454
rect 530446 165218 530488 165454
rect 530168 165134 530488 165218
rect 530168 164898 530210 165134
rect 530446 164898 530488 165134
rect 530168 164866 530488 164898
rect 15754 150938 15786 151174
rect 16022 150938 16106 151174
rect 16342 150938 16374 151174
rect 15754 150854 16374 150938
rect 15754 150618 15786 150854
rect 16022 150618 16106 150854
rect 16342 150618 16374 150854
rect 15754 115174 16374 150618
rect 541714 154894 542334 190338
rect 541714 154658 541746 154894
rect 541982 154658 542066 154894
rect 542302 154658 542334 154894
rect 541714 154574 542334 154658
rect 541714 154338 541746 154574
rect 541982 154338 542066 154574
rect 542302 154338 542334 154574
rect 23288 147454 23608 147486
rect 23288 147218 23330 147454
rect 23566 147218 23608 147454
rect 23288 147134 23608 147218
rect 23288 146898 23330 147134
rect 23566 146898 23608 147134
rect 23288 146866 23608 146898
rect 33528 147454 33848 147486
rect 33528 147218 33570 147454
rect 33806 147218 33848 147454
rect 33528 147134 33848 147218
rect 33528 146898 33570 147134
rect 33806 146898 33848 147134
rect 33528 146866 33848 146898
rect 43768 147454 44088 147486
rect 43768 147218 43810 147454
rect 44046 147218 44088 147454
rect 43768 147134 44088 147218
rect 43768 146898 43810 147134
rect 44046 146898 44088 147134
rect 43768 146866 44088 146898
rect 54008 147454 54328 147486
rect 54008 147218 54050 147454
rect 54286 147218 54328 147454
rect 54008 147134 54328 147218
rect 54008 146898 54050 147134
rect 54286 146898 54328 147134
rect 54008 146866 54328 146898
rect 64248 147454 64568 147486
rect 64248 147218 64290 147454
rect 64526 147218 64568 147454
rect 64248 147134 64568 147218
rect 64248 146898 64290 147134
rect 64526 146898 64568 147134
rect 64248 146866 64568 146898
rect 74488 147454 74808 147486
rect 74488 147218 74530 147454
rect 74766 147218 74808 147454
rect 74488 147134 74808 147218
rect 74488 146898 74530 147134
rect 74766 146898 74808 147134
rect 74488 146866 74808 146898
rect 84728 147454 85048 147486
rect 84728 147218 84770 147454
rect 85006 147218 85048 147454
rect 84728 147134 85048 147218
rect 84728 146898 84770 147134
rect 85006 146898 85048 147134
rect 84728 146866 85048 146898
rect 94968 147454 95288 147486
rect 94968 147218 95010 147454
rect 95246 147218 95288 147454
rect 94968 147134 95288 147218
rect 94968 146898 95010 147134
rect 95246 146898 95288 147134
rect 94968 146866 95288 146898
rect 105208 147454 105528 147486
rect 105208 147218 105250 147454
rect 105486 147218 105528 147454
rect 105208 147134 105528 147218
rect 105208 146898 105250 147134
rect 105486 146898 105528 147134
rect 105208 146866 105528 146898
rect 115448 147454 115768 147486
rect 115448 147218 115490 147454
rect 115726 147218 115768 147454
rect 115448 147134 115768 147218
rect 115448 146898 115490 147134
rect 115726 146898 115768 147134
rect 115448 146866 115768 146898
rect 125688 147454 126008 147486
rect 125688 147218 125730 147454
rect 125966 147218 126008 147454
rect 125688 147134 126008 147218
rect 125688 146898 125730 147134
rect 125966 146898 126008 147134
rect 125688 146866 126008 146898
rect 135928 147454 136248 147486
rect 135928 147218 135970 147454
rect 136206 147218 136248 147454
rect 135928 147134 136248 147218
rect 135928 146898 135970 147134
rect 136206 146898 136248 147134
rect 135928 146866 136248 146898
rect 146168 147454 146488 147486
rect 146168 147218 146210 147454
rect 146446 147218 146488 147454
rect 146168 147134 146488 147218
rect 146168 146898 146210 147134
rect 146446 146898 146488 147134
rect 146168 146866 146488 146898
rect 156408 147454 156728 147486
rect 156408 147218 156450 147454
rect 156686 147218 156728 147454
rect 156408 147134 156728 147218
rect 156408 146898 156450 147134
rect 156686 146898 156728 147134
rect 156408 146866 156728 146898
rect 166648 147454 166968 147486
rect 166648 147218 166690 147454
rect 166926 147218 166968 147454
rect 166648 147134 166968 147218
rect 166648 146898 166690 147134
rect 166926 146898 166968 147134
rect 166648 146866 166968 146898
rect 176888 147454 177208 147486
rect 176888 147218 176930 147454
rect 177166 147218 177208 147454
rect 176888 147134 177208 147218
rect 176888 146898 176930 147134
rect 177166 146898 177208 147134
rect 176888 146866 177208 146898
rect 187128 147454 187448 147486
rect 187128 147218 187170 147454
rect 187406 147218 187448 147454
rect 187128 147134 187448 147218
rect 187128 146898 187170 147134
rect 187406 146898 187448 147134
rect 187128 146866 187448 146898
rect 197368 147454 197688 147486
rect 197368 147218 197410 147454
rect 197646 147218 197688 147454
rect 197368 147134 197688 147218
rect 197368 146898 197410 147134
rect 197646 146898 197688 147134
rect 197368 146866 197688 146898
rect 207608 147454 207928 147486
rect 207608 147218 207650 147454
rect 207886 147218 207928 147454
rect 207608 147134 207928 147218
rect 207608 146898 207650 147134
rect 207886 146898 207928 147134
rect 207608 146866 207928 146898
rect 217848 147454 218168 147486
rect 217848 147218 217890 147454
rect 218126 147218 218168 147454
rect 217848 147134 218168 147218
rect 217848 146898 217890 147134
rect 218126 146898 218168 147134
rect 217848 146866 218168 146898
rect 228088 147454 228408 147486
rect 228088 147218 228130 147454
rect 228366 147218 228408 147454
rect 228088 147134 228408 147218
rect 228088 146898 228130 147134
rect 228366 146898 228408 147134
rect 228088 146866 228408 146898
rect 238328 147454 238648 147486
rect 238328 147218 238370 147454
rect 238606 147218 238648 147454
rect 238328 147134 238648 147218
rect 238328 146898 238370 147134
rect 238606 146898 238648 147134
rect 238328 146866 238648 146898
rect 248568 147454 248888 147486
rect 248568 147218 248610 147454
rect 248846 147218 248888 147454
rect 248568 147134 248888 147218
rect 248568 146898 248610 147134
rect 248846 146898 248888 147134
rect 248568 146866 248888 146898
rect 258808 147454 259128 147486
rect 258808 147218 258850 147454
rect 259086 147218 259128 147454
rect 258808 147134 259128 147218
rect 258808 146898 258850 147134
rect 259086 146898 259128 147134
rect 258808 146866 259128 146898
rect 269048 147454 269368 147486
rect 269048 147218 269090 147454
rect 269326 147218 269368 147454
rect 269048 147134 269368 147218
rect 269048 146898 269090 147134
rect 269326 146898 269368 147134
rect 269048 146866 269368 146898
rect 279288 147454 279608 147486
rect 279288 147218 279330 147454
rect 279566 147218 279608 147454
rect 279288 147134 279608 147218
rect 279288 146898 279330 147134
rect 279566 146898 279608 147134
rect 279288 146866 279608 146898
rect 289528 147454 289848 147486
rect 289528 147218 289570 147454
rect 289806 147218 289848 147454
rect 289528 147134 289848 147218
rect 289528 146898 289570 147134
rect 289806 146898 289848 147134
rect 289528 146866 289848 146898
rect 299768 147454 300088 147486
rect 299768 147218 299810 147454
rect 300046 147218 300088 147454
rect 299768 147134 300088 147218
rect 299768 146898 299810 147134
rect 300046 146898 300088 147134
rect 299768 146866 300088 146898
rect 310008 147454 310328 147486
rect 310008 147218 310050 147454
rect 310286 147218 310328 147454
rect 310008 147134 310328 147218
rect 310008 146898 310050 147134
rect 310286 146898 310328 147134
rect 310008 146866 310328 146898
rect 320248 147454 320568 147486
rect 320248 147218 320290 147454
rect 320526 147218 320568 147454
rect 320248 147134 320568 147218
rect 320248 146898 320290 147134
rect 320526 146898 320568 147134
rect 320248 146866 320568 146898
rect 330488 147454 330808 147486
rect 330488 147218 330530 147454
rect 330766 147218 330808 147454
rect 330488 147134 330808 147218
rect 330488 146898 330530 147134
rect 330766 146898 330808 147134
rect 330488 146866 330808 146898
rect 340728 147454 341048 147486
rect 340728 147218 340770 147454
rect 341006 147218 341048 147454
rect 340728 147134 341048 147218
rect 340728 146898 340770 147134
rect 341006 146898 341048 147134
rect 340728 146866 341048 146898
rect 350968 147454 351288 147486
rect 350968 147218 351010 147454
rect 351246 147218 351288 147454
rect 350968 147134 351288 147218
rect 350968 146898 351010 147134
rect 351246 146898 351288 147134
rect 350968 146866 351288 146898
rect 361208 147454 361528 147486
rect 361208 147218 361250 147454
rect 361486 147218 361528 147454
rect 361208 147134 361528 147218
rect 361208 146898 361250 147134
rect 361486 146898 361528 147134
rect 361208 146866 361528 146898
rect 371448 147454 371768 147486
rect 371448 147218 371490 147454
rect 371726 147218 371768 147454
rect 371448 147134 371768 147218
rect 371448 146898 371490 147134
rect 371726 146898 371768 147134
rect 371448 146866 371768 146898
rect 381688 147454 382008 147486
rect 381688 147218 381730 147454
rect 381966 147218 382008 147454
rect 381688 147134 382008 147218
rect 381688 146898 381730 147134
rect 381966 146898 382008 147134
rect 381688 146866 382008 146898
rect 391928 147454 392248 147486
rect 391928 147218 391970 147454
rect 392206 147218 392248 147454
rect 391928 147134 392248 147218
rect 391928 146898 391970 147134
rect 392206 146898 392248 147134
rect 391928 146866 392248 146898
rect 402168 147454 402488 147486
rect 402168 147218 402210 147454
rect 402446 147218 402488 147454
rect 402168 147134 402488 147218
rect 402168 146898 402210 147134
rect 402446 146898 402488 147134
rect 402168 146866 402488 146898
rect 412408 147454 412728 147486
rect 412408 147218 412450 147454
rect 412686 147218 412728 147454
rect 412408 147134 412728 147218
rect 412408 146898 412450 147134
rect 412686 146898 412728 147134
rect 412408 146866 412728 146898
rect 422648 147454 422968 147486
rect 422648 147218 422690 147454
rect 422926 147218 422968 147454
rect 422648 147134 422968 147218
rect 422648 146898 422690 147134
rect 422926 146898 422968 147134
rect 422648 146866 422968 146898
rect 432888 147454 433208 147486
rect 432888 147218 432930 147454
rect 433166 147218 433208 147454
rect 432888 147134 433208 147218
rect 432888 146898 432930 147134
rect 433166 146898 433208 147134
rect 432888 146866 433208 146898
rect 443128 147454 443448 147486
rect 443128 147218 443170 147454
rect 443406 147218 443448 147454
rect 443128 147134 443448 147218
rect 443128 146898 443170 147134
rect 443406 146898 443448 147134
rect 443128 146866 443448 146898
rect 453368 147454 453688 147486
rect 453368 147218 453410 147454
rect 453646 147218 453688 147454
rect 453368 147134 453688 147218
rect 453368 146898 453410 147134
rect 453646 146898 453688 147134
rect 453368 146866 453688 146898
rect 463608 147454 463928 147486
rect 463608 147218 463650 147454
rect 463886 147218 463928 147454
rect 463608 147134 463928 147218
rect 463608 146898 463650 147134
rect 463886 146898 463928 147134
rect 463608 146866 463928 146898
rect 473848 147454 474168 147486
rect 473848 147218 473890 147454
rect 474126 147218 474168 147454
rect 473848 147134 474168 147218
rect 473848 146898 473890 147134
rect 474126 146898 474168 147134
rect 473848 146866 474168 146898
rect 484088 147454 484408 147486
rect 484088 147218 484130 147454
rect 484366 147218 484408 147454
rect 484088 147134 484408 147218
rect 484088 146898 484130 147134
rect 484366 146898 484408 147134
rect 484088 146866 484408 146898
rect 494328 147454 494648 147486
rect 494328 147218 494370 147454
rect 494606 147218 494648 147454
rect 494328 147134 494648 147218
rect 494328 146898 494370 147134
rect 494606 146898 494648 147134
rect 494328 146866 494648 146898
rect 504568 147454 504888 147486
rect 504568 147218 504610 147454
rect 504846 147218 504888 147454
rect 504568 147134 504888 147218
rect 504568 146898 504610 147134
rect 504846 146898 504888 147134
rect 504568 146866 504888 146898
rect 514808 147454 515128 147486
rect 514808 147218 514850 147454
rect 515086 147218 515128 147454
rect 514808 147134 515128 147218
rect 514808 146898 514850 147134
rect 515086 146898 515128 147134
rect 514808 146866 515128 146898
rect 525048 147454 525368 147486
rect 525048 147218 525090 147454
rect 525326 147218 525368 147454
rect 525048 147134 525368 147218
rect 525048 146898 525090 147134
rect 525326 146898 525368 147134
rect 525048 146866 525368 146898
rect 535288 147454 535608 147486
rect 535288 147218 535330 147454
rect 535566 147218 535608 147454
rect 535288 147134 535608 147218
rect 535288 146898 535330 147134
rect 535566 146898 535608 147134
rect 535288 146866 535608 146898
rect 28408 129454 28728 129486
rect 28408 129218 28450 129454
rect 28686 129218 28728 129454
rect 28408 129134 28728 129218
rect 28408 128898 28450 129134
rect 28686 128898 28728 129134
rect 28408 128866 28728 128898
rect 38648 129454 38968 129486
rect 38648 129218 38690 129454
rect 38926 129218 38968 129454
rect 38648 129134 38968 129218
rect 38648 128898 38690 129134
rect 38926 128898 38968 129134
rect 38648 128866 38968 128898
rect 48888 129454 49208 129486
rect 48888 129218 48930 129454
rect 49166 129218 49208 129454
rect 48888 129134 49208 129218
rect 48888 128898 48930 129134
rect 49166 128898 49208 129134
rect 48888 128866 49208 128898
rect 59128 129454 59448 129486
rect 59128 129218 59170 129454
rect 59406 129218 59448 129454
rect 59128 129134 59448 129218
rect 59128 128898 59170 129134
rect 59406 128898 59448 129134
rect 59128 128866 59448 128898
rect 69368 129454 69688 129486
rect 69368 129218 69410 129454
rect 69646 129218 69688 129454
rect 69368 129134 69688 129218
rect 69368 128898 69410 129134
rect 69646 128898 69688 129134
rect 69368 128866 69688 128898
rect 79608 129454 79928 129486
rect 79608 129218 79650 129454
rect 79886 129218 79928 129454
rect 79608 129134 79928 129218
rect 79608 128898 79650 129134
rect 79886 128898 79928 129134
rect 79608 128866 79928 128898
rect 89848 129454 90168 129486
rect 89848 129218 89890 129454
rect 90126 129218 90168 129454
rect 89848 129134 90168 129218
rect 89848 128898 89890 129134
rect 90126 128898 90168 129134
rect 89848 128866 90168 128898
rect 100088 129454 100408 129486
rect 100088 129218 100130 129454
rect 100366 129218 100408 129454
rect 100088 129134 100408 129218
rect 100088 128898 100130 129134
rect 100366 128898 100408 129134
rect 100088 128866 100408 128898
rect 110328 129454 110648 129486
rect 110328 129218 110370 129454
rect 110606 129218 110648 129454
rect 110328 129134 110648 129218
rect 110328 128898 110370 129134
rect 110606 128898 110648 129134
rect 110328 128866 110648 128898
rect 120568 129454 120888 129486
rect 120568 129218 120610 129454
rect 120846 129218 120888 129454
rect 120568 129134 120888 129218
rect 120568 128898 120610 129134
rect 120846 128898 120888 129134
rect 120568 128866 120888 128898
rect 130808 129454 131128 129486
rect 130808 129218 130850 129454
rect 131086 129218 131128 129454
rect 130808 129134 131128 129218
rect 130808 128898 130850 129134
rect 131086 128898 131128 129134
rect 130808 128866 131128 128898
rect 141048 129454 141368 129486
rect 141048 129218 141090 129454
rect 141326 129218 141368 129454
rect 141048 129134 141368 129218
rect 141048 128898 141090 129134
rect 141326 128898 141368 129134
rect 141048 128866 141368 128898
rect 151288 129454 151608 129486
rect 151288 129218 151330 129454
rect 151566 129218 151608 129454
rect 151288 129134 151608 129218
rect 151288 128898 151330 129134
rect 151566 128898 151608 129134
rect 151288 128866 151608 128898
rect 161528 129454 161848 129486
rect 161528 129218 161570 129454
rect 161806 129218 161848 129454
rect 161528 129134 161848 129218
rect 161528 128898 161570 129134
rect 161806 128898 161848 129134
rect 161528 128866 161848 128898
rect 171768 129454 172088 129486
rect 171768 129218 171810 129454
rect 172046 129218 172088 129454
rect 171768 129134 172088 129218
rect 171768 128898 171810 129134
rect 172046 128898 172088 129134
rect 171768 128866 172088 128898
rect 182008 129454 182328 129486
rect 182008 129218 182050 129454
rect 182286 129218 182328 129454
rect 182008 129134 182328 129218
rect 182008 128898 182050 129134
rect 182286 128898 182328 129134
rect 182008 128866 182328 128898
rect 192248 129454 192568 129486
rect 192248 129218 192290 129454
rect 192526 129218 192568 129454
rect 192248 129134 192568 129218
rect 192248 128898 192290 129134
rect 192526 128898 192568 129134
rect 192248 128866 192568 128898
rect 202488 129454 202808 129486
rect 202488 129218 202530 129454
rect 202766 129218 202808 129454
rect 202488 129134 202808 129218
rect 202488 128898 202530 129134
rect 202766 128898 202808 129134
rect 202488 128866 202808 128898
rect 212728 129454 213048 129486
rect 212728 129218 212770 129454
rect 213006 129218 213048 129454
rect 212728 129134 213048 129218
rect 212728 128898 212770 129134
rect 213006 128898 213048 129134
rect 212728 128866 213048 128898
rect 222968 129454 223288 129486
rect 222968 129218 223010 129454
rect 223246 129218 223288 129454
rect 222968 129134 223288 129218
rect 222968 128898 223010 129134
rect 223246 128898 223288 129134
rect 222968 128866 223288 128898
rect 233208 129454 233528 129486
rect 233208 129218 233250 129454
rect 233486 129218 233528 129454
rect 233208 129134 233528 129218
rect 233208 128898 233250 129134
rect 233486 128898 233528 129134
rect 233208 128866 233528 128898
rect 243448 129454 243768 129486
rect 243448 129218 243490 129454
rect 243726 129218 243768 129454
rect 243448 129134 243768 129218
rect 243448 128898 243490 129134
rect 243726 128898 243768 129134
rect 243448 128866 243768 128898
rect 253688 129454 254008 129486
rect 253688 129218 253730 129454
rect 253966 129218 254008 129454
rect 253688 129134 254008 129218
rect 253688 128898 253730 129134
rect 253966 128898 254008 129134
rect 253688 128866 254008 128898
rect 263928 129454 264248 129486
rect 263928 129218 263970 129454
rect 264206 129218 264248 129454
rect 263928 129134 264248 129218
rect 263928 128898 263970 129134
rect 264206 128898 264248 129134
rect 263928 128866 264248 128898
rect 274168 129454 274488 129486
rect 274168 129218 274210 129454
rect 274446 129218 274488 129454
rect 274168 129134 274488 129218
rect 274168 128898 274210 129134
rect 274446 128898 274488 129134
rect 274168 128866 274488 128898
rect 284408 129454 284728 129486
rect 284408 129218 284450 129454
rect 284686 129218 284728 129454
rect 284408 129134 284728 129218
rect 284408 128898 284450 129134
rect 284686 128898 284728 129134
rect 284408 128866 284728 128898
rect 294648 129454 294968 129486
rect 294648 129218 294690 129454
rect 294926 129218 294968 129454
rect 294648 129134 294968 129218
rect 294648 128898 294690 129134
rect 294926 128898 294968 129134
rect 294648 128866 294968 128898
rect 304888 129454 305208 129486
rect 304888 129218 304930 129454
rect 305166 129218 305208 129454
rect 304888 129134 305208 129218
rect 304888 128898 304930 129134
rect 305166 128898 305208 129134
rect 304888 128866 305208 128898
rect 315128 129454 315448 129486
rect 315128 129218 315170 129454
rect 315406 129218 315448 129454
rect 315128 129134 315448 129218
rect 315128 128898 315170 129134
rect 315406 128898 315448 129134
rect 315128 128866 315448 128898
rect 325368 129454 325688 129486
rect 325368 129218 325410 129454
rect 325646 129218 325688 129454
rect 325368 129134 325688 129218
rect 325368 128898 325410 129134
rect 325646 128898 325688 129134
rect 325368 128866 325688 128898
rect 335608 129454 335928 129486
rect 335608 129218 335650 129454
rect 335886 129218 335928 129454
rect 335608 129134 335928 129218
rect 335608 128898 335650 129134
rect 335886 128898 335928 129134
rect 335608 128866 335928 128898
rect 345848 129454 346168 129486
rect 345848 129218 345890 129454
rect 346126 129218 346168 129454
rect 345848 129134 346168 129218
rect 345848 128898 345890 129134
rect 346126 128898 346168 129134
rect 345848 128866 346168 128898
rect 356088 129454 356408 129486
rect 356088 129218 356130 129454
rect 356366 129218 356408 129454
rect 356088 129134 356408 129218
rect 356088 128898 356130 129134
rect 356366 128898 356408 129134
rect 356088 128866 356408 128898
rect 366328 129454 366648 129486
rect 366328 129218 366370 129454
rect 366606 129218 366648 129454
rect 366328 129134 366648 129218
rect 366328 128898 366370 129134
rect 366606 128898 366648 129134
rect 366328 128866 366648 128898
rect 376568 129454 376888 129486
rect 376568 129218 376610 129454
rect 376846 129218 376888 129454
rect 376568 129134 376888 129218
rect 376568 128898 376610 129134
rect 376846 128898 376888 129134
rect 376568 128866 376888 128898
rect 386808 129454 387128 129486
rect 386808 129218 386850 129454
rect 387086 129218 387128 129454
rect 386808 129134 387128 129218
rect 386808 128898 386850 129134
rect 387086 128898 387128 129134
rect 386808 128866 387128 128898
rect 397048 129454 397368 129486
rect 397048 129218 397090 129454
rect 397326 129218 397368 129454
rect 397048 129134 397368 129218
rect 397048 128898 397090 129134
rect 397326 128898 397368 129134
rect 397048 128866 397368 128898
rect 407288 129454 407608 129486
rect 407288 129218 407330 129454
rect 407566 129218 407608 129454
rect 407288 129134 407608 129218
rect 407288 128898 407330 129134
rect 407566 128898 407608 129134
rect 407288 128866 407608 128898
rect 417528 129454 417848 129486
rect 417528 129218 417570 129454
rect 417806 129218 417848 129454
rect 417528 129134 417848 129218
rect 417528 128898 417570 129134
rect 417806 128898 417848 129134
rect 417528 128866 417848 128898
rect 427768 129454 428088 129486
rect 427768 129218 427810 129454
rect 428046 129218 428088 129454
rect 427768 129134 428088 129218
rect 427768 128898 427810 129134
rect 428046 128898 428088 129134
rect 427768 128866 428088 128898
rect 438008 129454 438328 129486
rect 438008 129218 438050 129454
rect 438286 129218 438328 129454
rect 438008 129134 438328 129218
rect 438008 128898 438050 129134
rect 438286 128898 438328 129134
rect 438008 128866 438328 128898
rect 448248 129454 448568 129486
rect 448248 129218 448290 129454
rect 448526 129218 448568 129454
rect 448248 129134 448568 129218
rect 448248 128898 448290 129134
rect 448526 128898 448568 129134
rect 448248 128866 448568 128898
rect 458488 129454 458808 129486
rect 458488 129218 458530 129454
rect 458766 129218 458808 129454
rect 458488 129134 458808 129218
rect 458488 128898 458530 129134
rect 458766 128898 458808 129134
rect 458488 128866 458808 128898
rect 468728 129454 469048 129486
rect 468728 129218 468770 129454
rect 469006 129218 469048 129454
rect 468728 129134 469048 129218
rect 468728 128898 468770 129134
rect 469006 128898 469048 129134
rect 468728 128866 469048 128898
rect 478968 129454 479288 129486
rect 478968 129218 479010 129454
rect 479246 129218 479288 129454
rect 478968 129134 479288 129218
rect 478968 128898 479010 129134
rect 479246 128898 479288 129134
rect 478968 128866 479288 128898
rect 489208 129454 489528 129486
rect 489208 129218 489250 129454
rect 489486 129218 489528 129454
rect 489208 129134 489528 129218
rect 489208 128898 489250 129134
rect 489486 128898 489528 129134
rect 489208 128866 489528 128898
rect 499448 129454 499768 129486
rect 499448 129218 499490 129454
rect 499726 129218 499768 129454
rect 499448 129134 499768 129218
rect 499448 128898 499490 129134
rect 499726 128898 499768 129134
rect 499448 128866 499768 128898
rect 509688 129454 510008 129486
rect 509688 129218 509730 129454
rect 509966 129218 510008 129454
rect 509688 129134 510008 129218
rect 509688 128898 509730 129134
rect 509966 128898 510008 129134
rect 509688 128866 510008 128898
rect 519928 129454 520248 129486
rect 519928 129218 519970 129454
rect 520206 129218 520248 129454
rect 519928 129134 520248 129218
rect 519928 128898 519970 129134
rect 520206 128898 520248 129134
rect 519928 128866 520248 128898
rect 530168 129454 530488 129486
rect 530168 129218 530210 129454
rect 530446 129218 530488 129454
rect 530168 129134 530488 129218
rect 530168 128898 530210 129134
rect 530446 128898 530488 129134
rect 530168 128866 530488 128898
rect 15754 114938 15786 115174
rect 16022 114938 16106 115174
rect 16342 114938 16374 115174
rect 15754 114854 16374 114938
rect 15754 114618 15786 114854
rect 16022 114618 16106 114854
rect 16342 114618 16374 114854
rect 15754 79174 16374 114618
rect 541714 118894 542334 154338
rect 541714 118658 541746 118894
rect 541982 118658 542066 118894
rect 542302 118658 542334 118894
rect 541714 118574 542334 118658
rect 541714 118338 541746 118574
rect 541982 118338 542066 118574
rect 542302 118338 542334 118574
rect 23288 111454 23608 111486
rect 23288 111218 23330 111454
rect 23566 111218 23608 111454
rect 23288 111134 23608 111218
rect 23288 110898 23330 111134
rect 23566 110898 23608 111134
rect 23288 110866 23608 110898
rect 33528 111454 33848 111486
rect 33528 111218 33570 111454
rect 33806 111218 33848 111454
rect 33528 111134 33848 111218
rect 33528 110898 33570 111134
rect 33806 110898 33848 111134
rect 33528 110866 33848 110898
rect 43768 111454 44088 111486
rect 43768 111218 43810 111454
rect 44046 111218 44088 111454
rect 43768 111134 44088 111218
rect 43768 110898 43810 111134
rect 44046 110898 44088 111134
rect 43768 110866 44088 110898
rect 54008 111454 54328 111486
rect 54008 111218 54050 111454
rect 54286 111218 54328 111454
rect 54008 111134 54328 111218
rect 54008 110898 54050 111134
rect 54286 110898 54328 111134
rect 54008 110866 54328 110898
rect 64248 111454 64568 111486
rect 64248 111218 64290 111454
rect 64526 111218 64568 111454
rect 64248 111134 64568 111218
rect 64248 110898 64290 111134
rect 64526 110898 64568 111134
rect 64248 110866 64568 110898
rect 74488 111454 74808 111486
rect 74488 111218 74530 111454
rect 74766 111218 74808 111454
rect 74488 111134 74808 111218
rect 74488 110898 74530 111134
rect 74766 110898 74808 111134
rect 74488 110866 74808 110898
rect 84728 111454 85048 111486
rect 84728 111218 84770 111454
rect 85006 111218 85048 111454
rect 84728 111134 85048 111218
rect 84728 110898 84770 111134
rect 85006 110898 85048 111134
rect 84728 110866 85048 110898
rect 94968 111454 95288 111486
rect 94968 111218 95010 111454
rect 95246 111218 95288 111454
rect 94968 111134 95288 111218
rect 94968 110898 95010 111134
rect 95246 110898 95288 111134
rect 94968 110866 95288 110898
rect 105208 111454 105528 111486
rect 105208 111218 105250 111454
rect 105486 111218 105528 111454
rect 105208 111134 105528 111218
rect 105208 110898 105250 111134
rect 105486 110898 105528 111134
rect 105208 110866 105528 110898
rect 115448 111454 115768 111486
rect 115448 111218 115490 111454
rect 115726 111218 115768 111454
rect 115448 111134 115768 111218
rect 115448 110898 115490 111134
rect 115726 110898 115768 111134
rect 115448 110866 115768 110898
rect 125688 111454 126008 111486
rect 125688 111218 125730 111454
rect 125966 111218 126008 111454
rect 125688 111134 126008 111218
rect 125688 110898 125730 111134
rect 125966 110898 126008 111134
rect 125688 110866 126008 110898
rect 135928 111454 136248 111486
rect 135928 111218 135970 111454
rect 136206 111218 136248 111454
rect 135928 111134 136248 111218
rect 135928 110898 135970 111134
rect 136206 110898 136248 111134
rect 135928 110866 136248 110898
rect 146168 111454 146488 111486
rect 146168 111218 146210 111454
rect 146446 111218 146488 111454
rect 146168 111134 146488 111218
rect 146168 110898 146210 111134
rect 146446 110898 146488 111134
rect 146168 110866 146488 110898
rect 156408 111454 156728 111486
rect 156408 111218 156450 111454
rect 156686 111218 156728 111454
rect 156408 111134 156728 111218
rect 156408 110898 156450 111134
rect 156686 110898 156728 111134
rect 156408 110866 156728 110898
rect 166648 111454 166968 111486
rect 166648 111218 166690 111454
rect 166926 111218 166968 111454
rect 166648 111134 166968 111218
rect 166648 110898 166690 111134
rect 166926 110898 166968 111134
rect 166648 110866 166968 110898
rect 176888 111454 177208 111486
rect 176888 111218 176930 111454
rect 177166 111218 177208 111454
rect 176888 111134 177208 111218
rect 176888 110898 176930 111134
rect 177166 110898 177208 111134
rect 176888 110866 177208 110898
rect 187128 111454 187448 111486
rect 187128 111218 187170 111454
rect 187406 111218 187448 111454
rect 187128 111134 187448 111218
rect 187128 110898 187170 111134
rect 187406 110898 187448 111134
rect 187128 110866 187448 110898
rect 197368 111454 197688 111486
rect 197368 111218 197410 111454
rect 197646 111218 197688 111454
rect 197368 111134 197688 111218
rect 197368 110898 197410 111134
rect 197646 110898 197688 111134
rect 197368 110866 197688 110898
rect 207608 111454 207928 111486
rect 207608 111218 207650 111454
rect 207886 111218 207928 111454
rect 207608 111134 207928 111218
rect 207608 110898 207650 111134
rect 207886 110898 207928 111134
rect 207608 110866 207928 110898
rect 217848 111454 218168 111486
rect 217848 111218 217890 111454
rect 218126 111218 218168 111454
rect 217848 111134 218168 111218
rect 217848 110898 217890 111134
rect 218126 110898 218168 111134
rect 217848 110866 218168 110898
rect 228088 111454 228408 111486
rect 228088 111218 228130 111454
rect 228366 111218 228408 111454
rect 228088 111134 228408 111218
rect 228088 110898 228130 111134
rect 228366 110898 228408 111134
rect 228088 110866 228408 110898
rect 238328 111454 238648 111486
rect 238328 111218 238370 111454
rect 238606 111218 238648 111454
rect 238328 111134 238648 111218
rect 238328 110898 238370 111134
rect 238606 110898 238648 111134
rect 238328 110866 238648 110898
rect 248568 111454 248888 111486
rect 248568 111218 248610 111454
rect 248846 111218 248888 111454
rect 248568 111134 248888 111218
rect 248568 110898 248610 111134
rect 248846 110898 248888 111134
rect 248568 110866 248888 110898
rect 258808 111454 259128 111486
rect 258808 111218 258850 111454
rect 259086 111218 259128 111454
rect 258808 111134 259128 111218
rect 258808 110898 258850 111134
rect 259086 110898 259128 111134
rect 258808 110866 259128 110898
rect 269048 111454 269368 111486
rect 269048 111218 269090 111454
rect 269326 111218 269368 111454
rect 269048 111134 269368 111218
rect 269048 110898 269090 111134
rect 269326 110898 269368 111134
rect 269048 110866 269368 110898
rect 279288 111454 279608 111486
rect 279288 111218 279330 111454
rect 279566 111218 279608 111454
rect 279288 111134 279608 111218
rect 279288 110898 279330 111134
rect 279566 110898 279608 111134
rect 279288 110866 279608 110898
rect 289528 111454 289848 111486
rect 289528 111218 289570 111454
rect 289806 111218 289848 111454
rect 289528 111134 289848 111218
rect 289528 110898 289570 111134
rect 289806 110898 289848 111134
rect 289528 110866 289848 110898
rect 299768 111454 300088 111486
rect 299768 111218 299810 111454
rect 300046 111218 300088 111454
rect 299768 111134 300088 111218
rect 299768 110898 299810 111134
rect 300046 110898 300088 111134
rect 299768 110866 300088 110898
rect 310008 111454 310328 111486
rect 310008 111218 310050 111454
rect 310286 111218 310328 111454
rect 310008 111134 310328 111218
rect 310008 110898 310050 111134
rect 310286 110898 310328 111134
rect 310008 110866 310328 110898
rect 320248 111454 320568 111486
rect 320248 111218 320290 111454
rect 320526 111218 320568 111454
rect 320248 111134 320568 111218
rect 320248 110898 320290 111134
rect 320526 110898 320568 111134
rect 320248 110866 320568 110898
rect 330488 111454 330808 111486
rect 330488 111218 330530 111454
rect 330766 111218 330808 111454
rect 330488 111134 330808 111218
rect 330488 110898 330530 111134
rect 330766 110898 330808 111134
rect 330488 110866 330808 110898
rect 340728 111454 341048 111486
rect 340728 111218 340770 111454
rect 341006 111218 341048 111454
rect 340728 111134 341048 111218
rect 340728 110898 340770 111134
rect 341006 110898 341048 111134
rect 340728 110866 341048 110898
rect 350968 111454 351288 111486
rect 350968 111218 351010 111454
rect 351246 111218 351288 111454
rect 350968 111134 351288 111218
rect 350968 110898 351010 111134
rect 351246 110898 351288 111134
rect 350968 110866 351288 110898
rect 361208 111454 361528 111486
rect 361208 111218 361250 111454
rect 361486 111218 361528 111454
rect 361208 111134 361528 111218
rect 361208 110898 361250 111134
rect 361486 110898 361528 111134
rect 361208 110866 361528 110898
rect 371448 111454 371768 111486
rect 371448 111218 371490 111454
rect 371726 111218 371768 111454
rect 371448 111134 371768 111218
rect 371448 110898 371490 111134
rect 371726 110898 371768 111134
rect 371448 110866 371768 110898
rect 381688 111454 382008 111486
rect 381688 111218 381730 111454
rect 381966 111218 382008 111454
rect 381688 111134 382008 111218
rect 381688 110898 381730 111134
rect 381966 110898 382008 111134
rect 381688 110866 382008 110898
rect 391928 111454 392248 111486
rect 391928 111218 391970 111454
rect 392206 111218 392248 111454
rect 391928 111134 392248 111218
rect 391928 110898 391970 111134
rect 392206 110898 392248 111134
rect 391928 110866 392248 110898
rect 402168 111454 402488 111486
rect 402168 111218 402210 111454
rect 402446 111218 402488 111454
rect 402168 111134 402488 111218
rect 402168 110898 402210 111134
rect 402446 110898 402488 111134
rect 402168 110866 402488 110898
rect 412408 111454 412728 111486
rect 412408 111218 412450 111454
rect 412686 111218 412728 111454
rect 412408 111134 412728 111218
rect 412408 110898 412450 111134
rect 412686 110898 412728 111134
rect 412408 110866 412728 110898
rect 422648 111454 422968 111486
rect 422648 111218 422690 111454
rect 422926 111218 422968 111454
rect 422648 111134 422968 111218
rect 422648 110898 422690 111134
rect 422926 110898 422968 111134
rect 422648 110866 422968 110898
rect 432888 111454 433208 111486
rect 432888 111218 432930 111454
rect 433166 111218 433208 111454
rect 432888 111134 433208 111218
rect 432888 110898 432930 111134
rect 433166 110898 433208 111134
rect 432888 110866 433208 110898
rect 443128 111454 443448 111486
rect 443128 111218 443170 111454
rect 443406 111218 443448 111454
rect 443128 111134 443448 111218
rect 443128 110898 443170 111134
rect 443406 110898 443448 111134
rect 443128 110866 443448 110898
rect 453368 111454 453688 111486
rect 453368 111218 453410 111454
rect 453646 111218 453688 111454
rect 453368 111134 453688 111218
rect 453368 110898 453410 111134
rect 453646 110898 453688 111134
rect 453368 110866 453688 110898
rect 463608 111454 463928 111486
rect 463608 111218 463650 111454
rect 463886 111218 463928 111454
rect 463608 111134 463928 111218
rect 463608 110898 463650 111134
rect 463886 110898 463928 111134
rect 463608 110866 463928 110898
rect 473848 111454 474168 111486
rect 473848 111218 473890 111454
rect 474126 111218 474168 111454
rect 473848 111134 474168 111218
rect 473848 110898 473890 111134
rect 474126 110898 474168 111134
rect 473848 110866 474168 110898
rect 484088 111454 484408 111486
rect 484088 111218 484130 111454
rect 484366 111218 484408 111454
rect 484088 111134 484408 111218
rect 484088 110898 484130 111134
rect 484366 110898 484408 111134
rect 484088 110866 484408 110898
rect 494328 111454 494648 111486
rect 494328 111218 494370 111454
rect 494606 111218 494648 111454
rect 494328 111134 494648 111218
rect 494328 110898 494370 111134
rect 494606 110898 494648 111134
rect 494328 110866 494648 110898
rect 504568 111454 504888 111486
rect 504568 111218 504610 111454
rect 504846 111218 504888 111454
rect 504568 111134 504888 111218
rect 504568 110898 504610 111134
rect 504846 110898 504888 111134
rect 504568 110866 504888 110898
rect 514808 111454 515128 111486
rect 514808 111218 514850 111454
rect 515086 111218 515128 111454
rect 514808 111134 515128 111218
rect 514808 110898 514850 111134
rect 515086 110898 515128 111134
rect 514808 110866 515128 110898
rect 525048 111454 525368 111486
rect 525048 111218 525090 111454
rect 525326 111218 525368 111454
rect 525048 111134 525368 111218
rect 525048 110898 525090 111134
rect 525326 110898 525368 111134
rect 525048 110866 525368 110898
rect 535288 111454 535608 111486
rect 535288 111218 535330 111454
rect 535566 111218 535608 111454
rect 535288 111134 535608 111218
rect 535288 110898 535330 111134
rect 535566 110898 535608 111134
rect 535288 110866 535608 110898
rect 28408 93454 28728 93486
rect 28408 93218 28450 93454
rect 28686 93218 28728 93454
rect 28408 93134 28728 93218
rect 28408 92898 28450 93134
rect 28686 92898 28728 93134
rect 28408 92866 28728 92898
rect 38648 93454 38968 93486
rect 38648 93218 38690 93454
rect 38926 93218 38968 93454
rect 38648 93134 38968 93218
rect 38648 92898 38690 93134
rect 38926 92898 38968 93134
rect 38648 92866 38968 92898
rect 48888 93454 49208 93486
rect 48888 93218 48930 93454
rect 49166 93218 49208 93454
rect 48888 93134 49208 93218
rect 48888 92898 48930 93134
rect 49166 92898 49208 93134
rect 48888 92866 49208 92898
rect 59128 93454 59448 93486
rect 59128 93218 59170 93454
rect 59406 93218 59448 93454
rect 59128 93134 59448 93218
rect 59128 92898 59170 93134
rect 59406 92898 59448 93134
rect 59128 92866 59448 92898
rect 69368 93454 69688 93486
rect 69368 93218 69410 93454
rect 69646 93218 69688 93454
rect 69368 93134 69688 93218
rect 69368 92898 69410 93134
rect 69646 92898 69688 93134
rect 69368 92866 69688 92898
rect 79608 93454 79928 93486
rect 79608 93218 79650 93454
rect 79886 93218 79928 93454
rect 79608 93134 79928 93218
rect 79608 92898 79650 93134
rect 79886 92898 79928 93134
rect 79608 92866 79928 92898
rect 89848 93454 90168 93486
rect 89848 93218 89890 93454
rect 90126 93218 90168 93454
rect 89848 93134 90168 93218
rect 89848 92898 89890 93134
rect 90126 92898 90168 93134
rect 89848 92866 90168 92898
rect 100088 93454 100408 93486
rect 100088 93218 100130 93454
rect 100366 93218 100408 93454
rect 100088 93134 100408 93218
rect 100088 92898 100130 93134
rect 100366 92898 100408 93134
rect 100088 92866 100408 92898
rect 110328 93454 110648 93486
rect 110328 93218 110370 93454
rect 110606 93218 110648 93454
rect 110328 93134 110648 93218
rect 110328 92898 110370 93134
rect 110606 92898 110648 93134
rect 110328 92866 110648 92898
rect 120568 93454 120888 93486
rect 120568 93218 120610 93454
rect 120846 93218 120888 93454
rect 120568 93134 120888 93218
rect 120568 92898 120610 93134
rect 120846 92898 120888 93134
rect 120568 92866 120888 92898
rect 130808 93454 131128 93486
rect 130808 93218 130850 93454
rect 131086 93218 131128 93454
rect 130808 93134 131128 93218
rect 130808 92898 130850 93134
rect 131086 92898 131128 93134
rect 130808 92866 131128 92898
rect 141048 93454 141368 93486
rect 141048 93218 141090 93454
rect 141326 93218 141368 93454
rect 141048 93134 141368 93218
rect 141048 92898 141090 93134
rect 141326 92898 141368 93134
rect 141048 92866 141368 92898
rect 151288 93454 151608 93486
rect 151288 93218 151330 93454
rect 151566 93218 151608 93454
rect 151288 93134 151608 93218
rect 151288 92898 151330 93134
rect 151566 92898 151608 93134
rect 151288 92866 151608 92898
rect 161528 93454 161848 93486
rect 161528 93218 161570 93454
rect 161806 93218 161848 93454
rect 161528 93134 161848 93218
rect 161528 92898 161570 93134
rect 161806 92898 161848 93134
rect 161528 92866 161848 92898
rect 171768 93454 172088 93486
rect 171768 93218 171810 93454
rect 172046 93218 172088 93454
rect 171768 93134 172088 93218
rect 171768 92898 171810 93134
rect 172046 92898 172088 93134
rect 171768 92866 172088 92898
rect 182008 93454 182328 93486
rect 182008 93218 182050 93454
rect 182286 93218 182328 93454
rect 182008 93134 182328 93218
rect 182008 92898 182050 93134
rect 182286 92898 182328 93134
rect 182008 92866 182328 92898
rect 192248 93454 192568 93486
rect 192248 93218 192290 93454
rect 192526 93218 192568 93454
rect 192248 93134 192568 93218
rect 192248 92898 192290 93134
rect 192526 92898 192568 93134
rect 192248 92866 192568 92898
rect 202488 93454 202808 93486
rect 202488 93218 202530 93454
rect 202766 93218 202808 93454
rect 202488 93134 202808 93218
rect 202488 92898 202530 93134
rect 202766 92898 202808 93134
rect 202488 92866 202808 92898
rect 212728 93454 213048 93486
rect 212728 93218 212770 93454
rect 213006 93218 213048 93454
rect 212728 93134 213048 93218
rect 212728 92898 212770 93134
rect 213006 92898 213048 93134
rect 212728 92866 213048 92898
rect 222968 93454 223288 93486
rect 222968 93218 223010 93454
rect 223246 93218 223288 93454
rect 222968 93134 223288 93218
rect 222968 92898 223010 93134
rect 223246 92898 223288 93134
rect 222968 92866 223288 92898
rect 233208 93454 233528 93486
rect 233208 93218 233250 93454
rect 233486 93218 233528 93454
rect 233208 93134 233528 93218
rect 233208 92898 233250 93134
rect 233486 92898 233528 93134
rect 233208 92866 233528 92898
rect 243448 93454 243768 93486
rect 243448 93218 243490 93454
rect 243726 93218 243768 93454
rect 243448 93134 243768 93218
rect 243448 92898 243490 93134
rect 243726 92898 243768 93134
rect 243448 92866 243768 92898
rect 253688 93454 254008 93486
rect 253688 93218 253730 93454
rect 253966 93218 254008 93454
rect 253688 93134 254008 93218
rect 253688 92898 253730 93134
rect 253966 92898 254008 93134
rect 253688 92866 254008 92898
rect 263928 93454 264248 93486
rect 263928 93218 263970 93454
rect 264206 93218 264248 93454
rect 263928 93134 264248 93218
rect 263928 92898 263970 93134
rect 264206 92898 264248 93134
rect 263928 92866 264248 92898
rect 274168 93454 274488 93486
rect 274168 93218 274210 93454
rect 274446 93218 274488 93454
rect 274168 93134 274488 93218
rect 274168 92898 274210 93134
rect 274446 92898 274488 93134
rect 274168 92866 274488 92898
rect 284408 93454 284728 93486
rect 284408 93218 284450 93454
rect 284686 93218 284728 93454
rect 284408 93134 284728 93218
rect 284408 92898 284450 93134
rect 284686 92898 284728 93134
rect 284408 92866 284728 92898
rect 294648 93454 294968 93486
rect 294648 93218 294690 93454
rect 294926 93218 294968 93454
rect 294648 93134 294968 93218
rect 294648 92898 294690 93134
rect 294926 92898 294968 93134
rect 294648 92866 294968 92898
rect 304888 93454 305208 93486
rect 304888 93218 304930 93454
rect 305166 93218 305208 93454
rect 304888 93134 305208 93218
rect 304888 92898 304930 93134
rect 305166 92898 305208 93134
rect 304888 92866 305208 92898
rect 315128 93454 315448 93486
rect 315128 93218 315170 93454
rect 315406 93218 315448 93454
rect 315128 93134 315448 93218
rect 315128 92898 315170 93134
rect 315406 92898 315448 93134
rect 315128 92866 315448 92898
rect 325368 93454 325688 93486
rect 325368 93218 325410 93454
rect 325646 93218 325688 93454
rect 325368 93134 325688 93218
rect 325368 92898 325410 93134
rect 325646 92898 325688 93134
rect 325368 92866 325688 92898
rect 335608 93454 335928 93486
rect 335608 93218 335650 93454
rect 335886 93218 335928 93454
rect 335608 93134 335928 93218
rect 335608 92898 335650 93134
rect 335886 92898 335928 93134
rect 335608 92866 335928 92898
rect 345848 93454 346168 93486
rect 345848 93218 345890 93454
rect 346126 93218 346168 93454
rect 345848 93134 346168 93218
rect 345848 92898 345890 93134
rect 346126 92898 346168 93134
rect 345848 92866 346168 92898
rect 356088 93454 356408 93486
rect 356088 93218 356130 93454
rect 356366 93218 356408 93454
rect 356088 93134 356408 93218
rect 356088 92898 356130 93134
rect 356366 92898 356408 93134
rect 356088 92866 356408 92898
rect 366328 93454 366648 93486
rect 366328 93218 366370 93454
rect 366606 93218 366648 93454
rect 366328 93134 366648 93218
rect 366328 92898 366370 93134
rect 366606 92898 366648 93134
rect 366328 92866 366648 92898
rect 376568 93454 376888 93486
rect 376568 93218 376610 93454
rect 376846 93218 376888 93454
rect 376568 93134 376888 93218
rect 376568 92898 376610 93134
rect 376846 92898 376888 93134
rect 376568 92866 376888 92898
rect 386808 93454 387128 93486
rect 386808 93218 386850 93454
rect 387086 93218 387128 93454
rect 386808 93134 387128 93218
rect 386808 92898 386850 93134
rect 387086 92898 387128 93134
rect 386808 92866 387128 92898
rect 397048 93454 397368 93486
rect 397048 93218 397090 93454
rect 397326 93218 397368 93454
rect 397048 93134 397368 93218
rect 397048 92898 397090 93134
rect 397326 92898 397368 93134
rect 397048 92866 397368 92898
rect 407288 93454 407608 93486
rect 407288 93218 407330 93454
rect 407566 93218 407608 93454
rect 407288 93134 407608 93218
rect 407288 92898 407330 93134
rect 407566 92898 407608 93134
rect 407288 92866 407608 92898
rect 417528 93454 417848 93486
rect 417528 93218 417570 93454
rect 417806 93218 417848 93454
rect 417528 93134 417848 93218
rect 417528 92898 417570 93134
rect 417806 92898 417848 93134
rect 417528 92866 417848 92898
rect 427768 93454 428088 93486
rect 427768 93218 427810 93454
rect 428046 93218 428088 93454
rect 427768 93134 428088 93218
rect 427768 92898 427810 93134
rect 428046 92898 428088 93134
rect 427768 92866 428088 92898
rect 438008 93454 438328 93486
rect 438008 93218 438050 93454
rect 438286 93218 438328 93454
rect 438008 93134 438328 93218
rect 438008 92898 438050 93134
rect 438286 92898 438328 93134
rect 438008 92866 438328 92898
rect 448248 93454 448568 93486
rect 448248 93218 448290 93454
rect 448526 93218 448568 93454
rect 448248 93134 448568 93218
rect 448248 92898 448290 93134
rect 448526 92898 448568 93134
rect 448248 92866 448568 92898
rect 458488 93454 458808 93486
rect 458488 93218 458530 93454
rect 458766 93218 458808 93454
rect 458488 93134 458808 93218
rect 458488 92898 458530 93134
rect 458766 92898 458808 93134
rect 458488 92866 458808 92898
rect 468728 93454 469048 93486
rect 468728 93218 468770 93454
rect 469006 93218 469048 93454
rect 468728 93134 469048 93218
rect 468728 92898 468770 93134
rect 469006 92898 469048 93134
rect 468728 92866 469048 92898
rect 478968 93454 479288 93486
rect 478968 93218 479010 93454
rect 479246 93218 479288 93454
rect 478968 93134 479288 93218
rect 478968 92898 479010 93134
rect 479246 92898 479288 93134
rect 478968 92866 479288 92898
rect 489208 93454 489528 93486
rect 489208 93218 489250 93454
rect 489486 93218 489528 93454
rect 489208 93134 489528 93218
rect 489208 92898 489250 93134
rect 489486 92898 489528 93134
rect 489208 92866 489528 92898
rect 499448 93454 499768 93486
rect 499448 93218 499490 93454
rect 499726 93218 499768 93454
rect 499448 93134 499768 93218
rect 499448 92898 499490 93134
rect 499726 92898 499768 93134
rect 499448 92866 499768 92898
rect 509688 93454 510008 93486
rect 509688 93218 509730 93454
rect 509966 93218 510008 93454
rect 509688 93134 510008 93218
rect 509688 92898 509730 93134
rect 509966 92898 510008 93134
rect 509688 92866 510008 92898
rect 519928 93454 520248 93486
rect 519928 93218 519970 93454
rect 520206 93218 520248 93454
rect 519928 93134 520248 93218
rect 519928 92898 519970 93134
rect 520206 92898 520248 93134
rect 519928 92866 520248 92898
rect 530168 93454 530488 93486
rect 530168 93218 530210 93454
rect 530446 93218 530488 93454
rect 530168 93134 530488 93218
rect 530168 92898 530210 93134
rect 530446 92898 530488 93134
rect 530168 92866 530488 92898
rect 15754 78938 15786 79174
rect 16022 78938 16106 79174
rect 16342 78938 16374 79174
rect 15754 78854 16374 78938
rect 15754 78618 15786 78854
rect 16022 78618 16106 78854
rect 16342 78618 16374 78854
rect 15754 43174 16374 78618
rect 541714 82894 542334 118338
rect 541714 82658 541746 82894
rect 541982 82658 542066 82894
rect 542302 82658 542334 82894
rect 541714 82574 542334 82658
rect 541714 82338 541746 82574
rect 541982 82338 542066 82574
rect 542302 82338 542334 82574
rect 23288 75454 23608 75486
rect 23288 75218 23330 75454
rect 23566 75218 23608 75454
rect 23288 75134 23608 75218
rect 23288 74898 23330 75134
rect 23566 74898 23608 75134
rect 23288 74866 23608 74898
rect 33528 75454 33848 75486
rect 33528 75218 33570 75454
rect 33806 75218 33848 75454
rect 33528 75134 33848 75218
rect 33528 74898 33570 75134
rect 33806 74898 33848 75134
rect 33528 74866 33848 74898
rect 43768 75454 44088 75486
rect 43768 75218 43810 75454
rect 44046 75218 44088 75454
rect 43768 75134 44088 75218
rect 43768 74898 43810 75134
rect 44046 74898 44088 75134
rect 43768 74866 44088 74898
rect 54008 75454 54328 75486
rect 54008 75218 54050 75454
rect 54286 75218 54328 75454
rect 54008 75134 54328 75218
rect 54008 74898 54050 75134
rect 54286 74898 54328 75134
rect 54008 74866 54328 74898
rect 64248 75454 64568 75486
rect 64248 75218 64290 75454
rect 64526 75218 64568 75454
rect 64248 75134 64568 75218
rect 64248 74898 64290 75134
rect 64526 74898 64568 75134
rect 64248 74866 64568 74898
rect 74488 75454 74808 75486
rect 74488 75218 74530 75454
rect 74766 75218 74808 75454
rect 74488 75134 74808 75218
rect 74488 74898 74530 75134
rect 74766 74898 74808 75134
rect 74488 74866 74808 74898
rect 84728 75454 85048 75486
rect 84728 75218 84770 75454
rect 85006 75218 85048 75454
rect 84728 75134 85048 75218
rect 84728 74898 84770 75134
rect 85006 74898 85048 75134
rect 84728 74866 85048 74898
rect 94968 75454 95288 75486
rect 94968 75218 95010 75454
rect 95246 75218 95288 75454
rect 94968 75134 95288 75218
rect 94968 74898 95010 75134
rect 95246 74898 95288 75134
rect 94968 74866 95288 74898
rect 105208 75454 105528 75486
rect 105208 75218 105250 75454
rect 105486 75218 105528 75454
rect 105208 75134 105528 75218
rect 105208 74898 105250 75134
rect 105486 74898 105528 75134
rect 105208 74866 105528 74898
rect 115448 75454 115768 75486
rect 115448 75218 115490 75454
rect 115726 75218 115768 75454
rect 115448 75134 115768 75218
rect 115448 74898 115490 75134
rect 115726 74898 115768 75134
rect 115448 74866 115768 74898
rect 125688 75454 126008 75486
rect 125688 75218 125730 75454
rect 125966 75218 126008 75454
rect 125688 75134 126008 75218
rect 125688 74898 125730 75134
rect 125966 74898 126008 75134
rect 125688 74866 126008 74898
rect 135928 75454 136248 75486
rect 135928 75218 135970 75454
rect 136206 75218 136248 75454
rect 135928 75134 136248 75218
rect 135928 74898 135970 75134
rect 136206 74898 136248 75134
rect 135928 74866 136248 74898
rect 146168 75454 146488 75486
rect 146168 75218 146210 75454
rect 146446 75218 146488 75454
rect 146168 75134 146488 75218
rect 146168 74898 146210 75134
rect 146446 74898 146488 75134
rect 146168 74866 146488 74898
rect 156408 75454 156728 75486
rect 156408 75218 156450 75454
rect 156686 75218 156728 75454
rect 156408 75134 156728 75218
rect 156408 74898 156450 75134
rect 156686 74898 156728 75134
rect 156408 74866 156728 74898
rect 166648 75454 166968 75486
rect 166648 75218 166690 75454
rect 166926 75218 166968 75454
rect 166648 75134 166968 75218
rect 166648 74898 166690 75134
rect 166926 74898 166968 75134
rect 166648 74866 166968 74898
rect 176888 75454 177208 75486
rect 176888 75218 176930 75454
rect 177166 75218 177208 75454
rect 176888 75134 177208 75218
rect 176888 74898 176930 75134
rect 177166 74898 177208 75134
rect 176888 74866 177208 74898
rect 187128 75454 187448 75486
rect 187128 75218 187170 75454
rect 187406 75218 187448 75454
rect 187128 75134 187448 75218
rect 187128 74898 187170 75134
rect 187406 74898 187448 75134
rect 187128 74866 187448 74898
rect 197368 75454 197688 75486
rect 197368 75218 197410 75454
rect 197646 75218 197688 75454
rect 197368 75134 197688 75218
rect 197368 74898 197410 75134
rect 197646 74898 197688 75134
rect 197368 74866 197688 74898
rect 207608 75454 207928 75486
rect 207608 75218 207650 75454
rect 207886 75218 207928 75454
rect 207608 75134 207928 75218
rect 207608 74898 207650 75134
rect 207886 74898 207928 75134
rect 207608 74866 207928 74898
rect 217848 75454 218168 75486
rect 217848 75218 217890 75454
rect 218126 75218 218168 75454
rect 217848 75134 218168 75218
rect 217848 74898 217890 75134
rect 218126 74898 218168 75134
rect 217848 74866 218168 74898
rect 228088 75454 228408 75486
rect 228088 75218 228130 75454
rect 228366 75218 228408 75454
rect 228088 75134 228408 75218
rect 228088 74898 228130 75134
rect 228366 74898 228408 75134
rect 228088 74866 228408 74898
rect 238328 75454 238648 75486
rect 238328 75218 238370 75454
rect 238606 75218 238648 75454
rect 238328 75134 238648 75218
rect 238328 74898 238370 75134
rect 238606 74898 238648 75134
rect 238328 74866 238648 74898
rect 248568 75454 248888 75486
rect 248568 75218 248610 75454
rect 248846 75218 248888 75454
rect 248568 75134 248888 75218
rect 248568 74898 248610 75134
rect 248846 74898 248888 75134
rect 248568 74866 248888 74898
rect 258808 75454 259128 75486
rect 258808 75218 258850 75454
rect 259086 75218 259128 75454
rect 258808 75134 259128 75218
rect 258808 74898 258850 75134
rect 259086 74898 259128 75134
rect 258808 74866 259128 74898
rect 269048 75454 269368 75486
rect 269048 75218 269090 75454
rect 269326 75218 269368 75454
rect 269048 75134 269368 75218
rect 269048 74898 269090 75134
rect 269326 74898 269368 75134
rect 269048 74866 269368 74898
rect 279288 75454 279608 75486
rect 279288 75218 279330 75454
rect 279566 75218 279608 75454
rect 279288 75134 279608 75218
rect 279288 74898 279330 75134
rect 279566 74898 279608 75134
rect 279288 74866 279608 74898
rect 289528 75454 289848 75486
rect 289528 75218 289570 75454
rect 289806 75218 289848 75454
rect 289528 75134 289848 75218
rect 289528 74898 289570 75134
rect 289806 74898 289848 75134
rect 289528 74866 289848 74898
rect 299768 75454 300088 75486
rect 299768 75218 299810 75454
rect 300046 75218 300088 75454
rect 299768 75134 300088 75218
rect 299768 74898 299810 75134
rect 300046 74898 300088 75134
rect 299768 74866 300088 74898
rect 310008 75454 310328 75486
rect 310008 75218 310050 75454
rect 310286 75218 310328 75454
rect 310008 75134 310328 75218
rect 310008 74898 310050 75134
rect 310286 74898 310328 75134
rect 310008 74866 310328 74898
rect 320248 75454 320568 75486
rect 320248 75218 320290 75454
rect 320526 75218 320568 75454
rect 320248 75134 320568 75218
rect 320248 74898 320290 75134
rect 320526 74898 320568 75134
rect 320248 74866 320568 74898
rect 330488 75454 330808 75486
rect 330488 75218 330530 75454
rect 330766 75218 330808 75454
rect 330488 75134 330808 75218
rect 330488 74898 330530 75134
rect 330766 74898 330808 75134
rect 330488 74866 330808 74898
rect 340728 75454 341048 75486
rect 340728 75218 340770 75454
rect 341006 75218 341048 75454
rect 340728 75134 341048 75218
rect 340728 74898 340770 75134
rect 341006 74898 341048 75134
rect 340728 74866 341048 74898
rect 350968 75454 351288 75486
rect 350968 75218 351010 75454
rect 351246 75218 351288 75454
rect 350968 75134 351288 75218
rect 350968 74898 351010 75134
rect 351246 74898 351288 75134
rect 350968 74866 351288 74898
rect 361208 75454 361528 75486
rect 361208 75218 361250 75454
rect 361486 75218 361528 75454
rect 361208 75134 361528 75218
rect 361208 74898 361250 75134
rect 361486 74898 361528 75134
rect 361208 74866 361528 74898
rect 371448 75454 371768 75486
rect 371448 75218 371490 75454
rect 371726 75218 371768 75454
rect 371448 75134 371768 75218
rect 371448 74898 371490 75134
rect 371726 74898 371768 75134
rect 371448 74866 371768 74898
rect 381688 75454 382008 75486
rect 381688 75218 381730 75454
rect 381966 75218 382008 75454
rect 381688 75134 382008 75218
rect 381688 74898 381730 75134
rect 381966 74898 382008 75134
rect 381688 74866 382008 74898
rect 391928 75454 392248 75486
rect 391928 75218 391970 75454
rect 392206 75218 392248 75454
rect 391928 75134 392248 75218
rect 391928 74898 391970 75134
rect 392206 74898 392248 75134
rect 391928 74866 392248 74898
rect 402168 75454 402488 75486
rect 402168 75218 402210 75454
rect 402446 75218 402488 75454
rect 402168 75134 402488 75218
rect 402168 74898 402210 75134
rect 402446 74898 402488 75134
rect 402168 74866 402488 74898
rect 412408 75454 412728 75486
rect 412408 75218 412450 75454
rect 412686 75218 412728 75454
rect 412408 75134 412728 75218
rect 412408 74898 412450 75134
rect 412686 74898 412728 75134
rect 412408 74866 412728 74898
rect 422648 75454 422968 75486
rect 422648 75218 422690 75454
rect 422926 75218 422968 75454
rect 422648 75134 422968 75218
rect 422648 74898 422690 75134
rect 422926 74898 422968 75134
rect 422648 74866 422968 74898
rect 432888 75454 433208 75486
rect 432888 75218 432930 75454
rect 433166 75218 433208 75454
rect 432888 75134 433208 75218
rect 432888 74898 432930 75134
rect 433166 74898 433208 75134
rect 432888 74866 433208 74898
rect 443128 75454 443448 75486
rect 443128 75218 443170 75454
rect 443406 75218 443448 75454
rect 443128 75134 443448 75218
rect 443128 74898 443170 75134
rect 443406 74898 443448 75134
rect 443128 74866 443448 74898
rect 453368 75454 453688 75486
rect 453368 75218 453410 75454
rect 453646 75218 453688 75454
rect 453368 75134 453688 75218
rect 453368 74898 453410 75134
rect 453646 74898 453688 75134
rect 453368 74866 453688 74898
rect 463608 75454 463928 75486
rect 463608 75218 463650 75454
rect 463886 75218 463928 75454
rect 463608 75134 463928 75218
rect 463608 74898 463650 75134
rect 463886 74898 463928 75134
rect 463608 74866 463928 74898
rect 473848 75454 474168 75486
rect 473848 75218 473890 75454
rect 474126 75218 474168 75454
rect 473848 75134 474168 75218
rect 473848 74898 473890 75134
rect 474126 74898 474168 75134
rect 473848 74866 474168 74898
rect 484088 75454 484408 75486
rect 484088 75218 484130 75454
rect 484366 75218 484408 75454
rect 484088 75134 484408 75218
rect 484088 74898 484130 75134
rect 484366 74898 484408 75134
rect 484088 74866 484408 74898
rect 494328 75454 494648 75486
rect 494328 75218 494370 75454
rect 494606 75218 494648 75454
rect 494328 75134 494648 75218
rect 494328 74898 494370 75134
rect 494606 74898 494648 75134
rect 494328 74866 494648 74898
rect 504568 75454 504888 75486
rect 504568 75218 504610 75454
rect 504846 75218 504888 75454
rect 504568 75134 504888 75218
rect 504568 74898 504610 75134
rect 504846 74898 504888 75134
rect 504568 74866 504888 74898
rect 514808 75454 515128 75486
rect 514808 75218 514850 75454
rect 515086 75218 515128 75454
rect 514808 75134 515128 75218
rect 514808 74898 514850 75134
rect 515086 74898 515128 75134
rect 514808 74866 515128 74898
rect 525048 75454 525368 75486
rect 525048 75218 525090 75454
rect 525326 75218 525368 75454
rect 525048 75134 525368 75218
rect 525048 74898 525090 75134
rect 525326 74898 525368 75134
rect 525048 74866 525368 74898
rect 535288 75454 535608 75486
rect 535288 75218 535330 75454
rect 535566 75218 535608 75454
rect 535288 75134 535608 75218
rect 535288 74898 535330 75134
rect 535566 74898 535608 75134
rect 535288 74866 535608 74898
rect 28408 57454 28728 57486
rect 28408 57218 28450 57454
rect 28686 57218 28728 57454
rect 28408 57134 28728 57218
rect 28408 56898 28450 57134
rect 28686 56898 28728 57134
rect 28408 56866 28728 56898
rect 38648 57454 38968 57486
rect 38648 57218 38690 57454
rect 38926 57218 38968 57454
rect 38648 57134 38968 57218
rect 38648 56898 38690 57134
rect 38926 56898 38968 57134
rect 38648 56866 38968 56898
rect 48888 57454 49208 57486
rect 48888 57218 48930 57454
rect 49166 57218 49208 57454
rect 48888 57134 49208 57218
rect 48888 56898 48930 57134
rect 49166 56898 49208 57134
rect 48888 56866 49208 56898
rect 59128 57454 59448 57486
rect 59128 57218 59170 57454
rect 59406 57218 59448 57454
rect 59128 57134 59448 57218
rect 59128 56898 59170 57134
rect 59406 56898 59448 57134
rect 59128 56866 59448 56898
rect 69368 57454 69688 57486
rect 69368 57218 69410 57454
rect 69646 57218 69688 57454
rect 69368 57134 69688 57218
rect 69368 56898 69410 57134
rect 69646 56898 69688 57134
rect 69368 56866 69688 56898
rect 79608 57454 79928 57486
rect 79608 57218 79650 57454
rect 79886 57218 79928 57454
rect 79608 57134 79928 57218
rect 79608 56898 79650 57134
rect 79886 56898 79928 57134
rect 79608 56866 79928 56898
rect 89848 57454 90168 57486
rect 89848 57218 89890 57454
rect 90126 57218 90168 57454
rect 89848 57134 90168 57218
rect 89848 56898 89890 57134
rect 90126 56898 90168 57134
rect 89848 56866 90168 56898
rect 100088 57454 100408 57486
rect 100088 57218 100130 57454
rect 100366 57218 100408 57454
rect 100088 57134 100408 57218
rect 100088 56898 100130 57134
rect 100366 56898 100408 57134
rect 100088 56866 100408 56898
rect 110328 57454 110648 57486
rect 110328 57218 110370 57454
rect 110606 57218 110648 57454
rect 110328 57134 110648 57218
rect 110328 56898 110370 57134
rect 110606 56898 110648 57134
rect 110328 56866 110648 56898
rect 120568 57454 120888 57486
rect 120568 57218 120610 57454
rect 120846 57218 120888 57454
rect 120568 57134 120888 57218
rect 120568 56898 120610 57134
rect 120846 56898 120888 57134
rect 120568 56866 120888 56898
rect 130808 57454 131128 57486
rect 130808 57218 130850 57454
rect 131086 57218 131128 57454
rect 130808 57134 131128 57218
rect 130808 56898 130850 57134
rect 131086 56898 131128 57134
rect 130808 56866 131128 56898
rect 141048 57454 141368 57486
rect 141048 57218 141090 57454
rect 141326 57218 141368 57454
rect 141048 57134 141368 57218
rect 141048 56898 141090 57134
rect 141326 56898 141368 57134
rect 141048 56866 141368 56898
rect 151288 57454 151608 57486
rect 151288 57218 151330 57454
rect 151566 57218 151608 57454
rect 151288 57134 151608 57218
rect 151288 56898 151330 57134
rect 151566 56898 151608 57134
rect 151288 56866 151608 56898
rect 161528 57454 161848 57486
rect 161528 57218 161570 57454
rect 161806 57218 161848 57454
rect 161528 57134 161848 57218
rect 161528 56898 161570 57134
rect 161806 56898 161848 57134
rect 161528 56866 161848 56898
rect 171768 57454 172088 57486
rect 171768 57218 171810 57454
rect 172046 57218 172088 57454
rect 171768 57134 172088 57218
rect 171768 56898 171810 57134
rect 172046 56898 172088 57134
rect 171768 56866 172088 56898
rect 182008 57454 182328 57486
rect 182008 57218 182050 57454
rect 182286 57218 182328 57454
rect 182008 57134 182328 57218
rect 182008 56898 182050 57134
rect 182286 56898 182328 57134
rect 182008 56866 182328 56898
rect 192248 57454 192568 57486
rect 192248 57218 192290 57454
rect 192526 57218 192568 57454
rect 192248 57134 192568 57218
rect 192248 56898 192290 57134
rect 192526 56898 192568 57134
rect 192248 56866 192568 56898
rect 202488 57454 202808 57486
rect 202488 57218 202530 57454
rect 202766 57218 202808 57454
rect 202488 57134 202808 57218
rect 202488 56898 202530 57134
rect 202766 56898 202808 57134
rect 202488 56866 202808 56898
rect 212728 57454 213048 57486
rect 212728 57218 212770 57454
rect 213006 57218 213048 57454
rect 212728 57134 213048 57218
rect 212728 56898 212770 57134
rect 213006 56898 213048 57134
rect 212728 56866 213048 56898
rect 222968 57454 223288 57486
rect 222968 57218 223010 57454
rect 223246 57218 223288 57454
rect 222968 57134 223288 57218
rect 222968 56898 223010 57134
rect 223246 56898 223288 57134
rect 222968 56866 223288 56898
rect 233208 57454 233528 57486
rect 233208 57218 233250 57454
rect 233486 57218 233528 57454
rect 233208 57134 233528 57218
rect 233208 56898 233250 57134
rect 233486 56898 233528 57134
rect 233208 56866 233528 56898
rect 243448 57454 243768 57486
rect 243448 57218 243490 57454
rect 243726 57218 243768 57454
rect 243448 57134 243768 57218
rect 243448 56898 243490 57134
rect 243726 56898 243768 57134
rect 243448 56866 243768 56898
rect 253688 57454 254008 57486
rect 253688 57218 253730 57454
rect 253966 57218 254008 57454
rect 253688 57134 254008 57218
rect 253688 56898 253730 57134
rect 253966 56898 254008 57134
rect 253688 56866 254008 56898
rect 263928 57454 264248 57486
rect 263928 57218 263970 57454
rect 264206 57218 264248 57454
rect 263928 57134 264248 57218
rect 263928 56898 263970 57134
rect 264206 56898 264248 57134
rect 263928 56866 264248 56898
rect 274168 57454 274488 57486
rect 274168 57218 274210 57454
rect 274446 57218 274488 57454
rect 274168 57134 274488 57218
rect 274168 56898 274210 57134
rect 274446 56898 274488 57134
rect 274168 56866 274488 56898
rect 284408 57454 284728 57486
rect 284408 57218 284450 57454
rect 284686 57218 284728 57454
rect 284408 57134 284728 57218
rect 284408 56898 284450 57134
rect 284686 56898 284728 57134
rect 284408 56866 284728 56898
rect 294648 57454 294968 57486
rect 294648 57218 294690 57454
rect 294926 57218 294968 57454
rect 294648 57134 294968 57218
rect 294648 56898 294690 57134
rect 294926 56898 294968 57134
rect 294648 56866 294968 56898
rect 304888 57454 305208 57486
rect 304888 57218 304930 57454
rect 305166 57218 305208 57454
rect 304888 57134 305208 57218
rect 304888 56898 304930 57134
rect 305166 56898 305208 57134
rect 304888 56866 305208 56898
rect 315128 57454 315448 57486
rect 315128 57218 315170 57454
rect 315406 57218 315448 57454
rect 315128 57134 315448 57218
rect 315128 56898 315170 57134
rect 315406 56898 315448 57134
rect 315128 56866 315448 56898
rect 325368 57454 325688 57486
rect 325368 57218 325410 57454
rect 325646 57218 325688 57454
rect 325368 57134 325688 57218
rect 325368 56898 325410 57134
rect 325646 56898 325688 57134
rect 325368 56866 325688 56898
rect 335608 57454 335928 57486
rect 335608 57218 335650 57454
rect 335886 57218 335928 57454
rect 335608 57134 335928 57218
rect 335608 56898 335650 57134
rect 335886 56898 335928 57134
rect 335608 56866 335928 56898
rect 345848 57454 346168 57486
rect 345848 57218 345890 57454
rect 346126 57218 346168 57454
rect 345848 57134 346168 57218
rect 345848 56898 345890 57134
rect 346126 56898 346168 57134
rect 345848 56866 346168 56898
rect 356088 57454 356408 57486
rect 356088 57218 356130 57454
rect 356366 57218 356408 57454
rect 356088 57134 356408 57218
rect 356088 56898 356130 57134
rect 356366 56898 356408 57134
rect 356088 56866 356408 56898
rect 366328 57454 366648 57486
rect 366328 57218 366370 57454
rect 366606 57218 366648 57454
rect 366328 57134 366648 57218
rect 366328 56898 366370 57134
rect 366606 56898 366648 57134
rect 366328 56866 366648 56898
rect 376568 57454 376888 57486
rect 376568 57218 376610 57454
rect 376846 57218 376888 57454
rect 376568 57134 376888 57218
rect 376568 56898 376610 57134
rect 376846 56898 376888 57134
rect 376568 56866 376888 56898
rect 386808 57454 387128 57486
rect 386808 57218 386850 57454
rect 387086 57218 387128 57454
rect 386808 57134 387128 57218
rect 386808 56898 386850 57134
rect 387086 56898 387128 57134
rect 386808 56866 387128 56898
rect 397048 57454 397368 57486
rect 397048 57218 397090 57454
rect 397326 57218 397368 57454
rect 397048 57134 397368 57218
rect 397048 56898 397090 57134
rect 397326 56898 397368 57134
rect 397048 56866 397368 56898
rect 407288 57454 407608 57486
rect 407288 57218 407330 57454
rect 407566 57218 407608 57454
rect 407288 57134 407608 57218
rect 407288 56898 407330 57134
rect 407566 56898 407608 57134
rect 407288 56866 407608 56898
rect 417528 57454 417848 57486
rect 417528 57218 417570 57454
rect 417806 57218 417848 57454
rect 417528 57134 417848 57218
rect 417528 56898 417570 57134
rect 417806 56898 417848 57134
rect 417528 56866 417848 56898
rect 427768 57454 428088 57486
rect 427768 57218 427810 57454
rect 428046 57218 428088 57454
rect 427768 57134 428088 57218
rect 427768 56898 427810 57134
rect 428046 56898 428088 57134
rect 427768 56866 428088 56898
rect 438008 57454 438328 57486
rect 438008 57218 438050 57454
rect 438286 57218 438328 57454
rect 438008 57134 438328 57218
rect 438008 56898 438050 57134
rect 438286 56898 438328 57134
rect 438008 56866 438328 56898
rect 448248 57454 448568 57486
rect 448248 57218 448290 57454
rect 448526 57218 448568 57454
rect 448248 57134 448568 57218
rect 448248 56898 448290 57134
rect 448526 56898 448568 57134
rect 448248 56866 448568 56898
rect 458488 57454 458808 57486
rect 458488 57218 458530 57454
rect 458766 57218 458808 57454
rect 458488 57134 458808 57218
rect 458488 56898 458530 57134
rect 458766 56898 458808 57134
rect 458488 56866 458808 56898
rect 468728 57454 469048 57486
rect 468728 57218 468770 57454
rect 469006 57218 469048 57454
rect 468728 57134 469048 57218
rect 468728 56898 468770 57134
rect 469006 56898 469048 57134
rect 468728 56866 469048 56898
rect 478968 57454 479288 57486
rect 478968 57218 479010 57454
rect 479246 57218 479288 57454
rect 478968 57134 479288 57218
rect 478968 56898 479010 57134
rect 479246 56898 479288 57134
rect 478968 56866 479288 56898
rect 489208 57454 489528 57486
rect 489208 57218 489250 57454
rect 489486 57218 489528 57454
rect 489208 57134 489528 57218
rect 489208 56898 489250 57134
rect 489486 56898 489528 57134
rect 489208 56866 489528 56898
rect 499448 57454 499768 57486
rect 499448 57218 499490 57454
rect 499726 57218 499768 57454
rect 499448 57134 499768 57218
rect 499448 56898 499490 57134
rect 499726 56898 499768 57134
rect 499448 56866 499768 56898
rect 509688 57454 510008 57486
rect 509688 57218 509730 57454
rect 509966 57218 510008 57454
rect 509688 57134 510008 57218
rect 509688 56898 509730 57134
rect 509966 56898 510008 57134
rect 509688 56866 510008 56898
rect 519928 57454 520248 57486
rect 519928 57218 519970 57454
rect 520206 57218 520248 57454
rect 519928 57134 520248 57218
rect 519928 56898 519970 57134
rect 520206 56898 520248 57134
rect 519928 56866 520248 56898
rect 530168 57454 530488 57486
rect 530168 57218 530210 57454
rect 530446 57218 530488 57454
rect 530168 57134 530488 57218
rect 530168 56898 530210 57134
rect 530446 56898 530488 57134
rect 530168 56866 530488 56898
rect 15754 42938 15786 43174
rect 16022 42938 16106 43174
rect 16342 42938 16374 43174
rect 15754 42854 16374 42938
rect 15754 42618 15786 42854
rect 16022 42618 16106 42854
rect 16342 42618 16374 42854
rect 15754 7174 16374 42618
rect 541714 46894 542334 82338
rect 541714 46658 541746 46894
rect 541982 46658 542066 46894
rect 542302 46658 542334 46894
rect 541714 46574 542334 46658
rect 541714 46338 541746 46574
rect 541982 46338 542066 46574
rect 542302 46338 542334 46574
rect 23288 39454 23608 39486
rect 23288 39218 23330 39454
rect 23566 39218 23608 39454
rect 23288 39134 23608 39218
rect 23288 38898 23330 39134
rect 23566 38898 23608 39134
rect 23288 38866 23608 38898
rect 33528 39454 33848 39486
rect 33528 39218 33570 39454
rect 33806 39218 33848 39454
rect 33528 39134 33848 39218
rect 33528 38898 33570 39134
rect 33806 38898 33848 39134
rect 33528 38866 33848 38898
rect 43768 39454 44088 39486
rect 43768 39218 43810 39454
rect 44046 39218 44088 39454
rect 43768 39134 44088 39218
rect 43768 38898 43810 39134
rect 44046 38898 44088 39134
rect 43768 38866 44088 38898
rect 54008 39454 54328 39486
rect 54008 39218 54050 39454
rect 54286 39218 54328 39454
rect 54008 39134 54328 39218
rect 54008 38898 54050 39134
rect 54286 38898 54328 39134
rect 54008 38866 54328 38898
rect 64248 39454 64568 39486
rect 64248 39218 64290 39454
rect 64526 39218 64568 39454
rect 64248 39134 64568 39218
rect 64248 38898 64290 39134
rect 64526 38898 64568 39134
rect 64248 38866 64568 38898
rect 74488 39454 74808 39486
rect 74488 39218 74530 39454
rect 74766 39218 74808 39454
rect 74488 39134 74808 39218
rect 74488 38898 74530 39134
rect 74766 38898 74808 39134
rect 74488 38866 74808 38898
rect 84728 39454 85048 39486
rect 84728 39218 84770 39454
rect 85006 39218 85048 39454
rect 84728 39134 85048 39218
rect 84728 38898 84770 39134
rect 85006 38898 85048 39134
rect 84728 38866 85048 38898
rect 94968 39454 95288 39486
rect 94968 39218 95010 39454
rect 95246 39218 95288 39454
rect 94968 39134 95288 39218
rect 94968 38898 95010 39134
rect 95246 38898 95288 39134
rect 94968 38866 95288 38898
rect 105208 39454 105528 39486
rect 105208 39218 105250 39454
rect 105486 39218 105528 39454
rect 105208 39134 105528 39218
rect 105208 38898 105250 39134
rect 105486 38898 105528 39134
rect 105208 38866 105528 38898
rect 115448 39454 115768 39486
rect 115448 39218 115490 39454
rect 115726 39218 115768 39454
rect 115448 39134 115768 39218
rect 115448 38898 115490 39134
rect 115726 38898 115768 39134
rect 115448 38866 115768 38898
rect 125688 39454 126008 39486
rect 125688 39218 125730 39454
rect 125966 39218 126008 39454
rect 125688 39134 126008 39218
rect 125688 38898 125730 39134
rect 125966 38898 126008 39134
rect 125688 38866 126008 38898
rect 135928 39454 136248 39486
rect 135928 39218 135970 39454
rect 136206 39218 136248 39454
rect 135928 39134 136248 39218
rect 135928 38898 135970 39134
rect 136206 38898 136248 39134
rect 135928 38866 136248 38898
rect 146168 39454 146488 39486
rect 146168 39218 146210 39454
rect 146446 39218 146488 39454
rect 146168 39134 146488 39218
rect 146168 38898 146210 39134
rect 146446 38898 146488 39134
rect 146168 38866 146488 38898
rect 156408 39454 156728 39486
rect 156408 39218 156450 39454
rect 156686 39218 156728 39454
rect 156408 39134 156728 39218
rect 156408 38898 156450 39134
rect 156686 38898 156728 39134
rect 156408 38866 156728 38898
rect 166648 39454 166968 39486
rect 166648 39218 166690 39454
rect 166926 39218 166968 39454
rect 166648 39134 166968 39218
rect 166648 38898 166690 39134
rect 166926 38898 166968 39134
rect 166648 38866 166968 38898
rect 176888 39454 177208 39486
rect 176888 39218 176930 39454
rect 177166 39218 177208 39454
rect 176888 39134 177208 39218
rect 176888 38898 176930 39134
rect 177166 38898 177208 39134
rect 176888 38866 177208 38898
rect 187128 39454 187448 39486
rect 187128 39218 187170 39454
rect 187406 39218 187448 39454
rect 187128 39134 187448 39218
rect 187128 38898 187170 39134
rect 187406 38898 187448 39134
rect 187128 38866 187448 38898
rect 197368 39454 197688 39486
rect 197368 39218 197410 39454
rect 197646 39218 197688 39454
rect 197368 39134 197688 39218
rect 197368 38898 197410 39134
rect 197646 38898 197688 39134
rect 197368 38866 197688 38898
rect 207608 39454 207928 39486
rect 207608 39218 207650 39454
rect 207886 39218 207928 39454
rect 207608 39134 207928 39218
rect 207608 38898 207650 39134
rect 207886 38898 207928 39134
rect 207608 38866 207928 38898
rect 217848 39454 218168 39486
rect 217848 39218 217890 39454
rect 218126 39218 218168 39454
rect 217848 39134 218168 39218
rect 217848 38898 217890 39134
rect 218126 38898 218168 39134
rect 217848 38866 218168 38898
rect 228088 39454 228408 39486
rect 228088 39218 228130 39454
rect 228366 39218 228408 39454
rect 228088 39134 228408 39218
rect 228088 38898 228130 39134
rect 228366 38898 228408 39134
rect 228088 38866 228408 38898
rect 238328 39454 238648 39486
rect 238328 39218 238370 39454
rect 238606 39218 238648 39454
rect 238328 39134 238648 39218
rect 238328 38898 238370 39134
rect 238606 38898 238648 39134
rect 238328 38866 238648 38898
rect 248568 39454 248888 39486
rect 248568 39218 248610 39454
rect 248846 39218 248888 39454
rect 248568 39134 248888 39218
rect 248568 38898 248610 39134
rect 248846 38898 248888 39134
rect 248568 38866 248888 38898
rect 258808 39454 259128 39486
rect 258808 39218 258850 39454
rect 259086 39218 259128 39454
rect 258808 39134 259128 39218
rect 258808 38898 258850 39134
rect 259086 38898 259128 39134
rect 258808 38866 259128 38898
rect 269048 39454 269368 39486
rect 269048 39218 269090 39454
rect 269326 39218 269368 39454
rect 269048 39134 269368 39218
rect 269048 38898 269090 39134
rect 269326 38898 269368 39134
rect 269048 38866 269368 38898
rect 279288 39454 279608 39486
rect 279288 39218 279330 39454
rect 279566 39218 279608 39454
rect 279288 39134 279608 39218
rect 279288 38898 279330 39134
rect 279566 38898 279608 39134
rect 279288 38866 279608 38898
rect 289528 39454 289848 39486
rect 289528 39218 289570 39454
rect 289806 39218 289848 39454
rect 289528 39134 289848 39218
rect 289528 38898 289570 39134
rect 289806 38898 289848 39134
rect 289528 38866 289848 38898
rect 299768 39454 300088 39486
rect 299768 39218 299810 39454
rect 300046 39218 300088 39454
rect 299768 39134 300088 39218
rect 299768 38898 299810 39134
rect 300046 38898 300088 39134
rect 299768 38866 300088 38898
rect 310008 39454 310328 39486
rect 310008 39218 310050 39454
rect 310286 39218 310328 39454
rect 310008 39134 310328 39218
rect 310008 38898 310050 39134
rect 310286 38898 310328 39134
rect 310008 38866 310328 38898
rect 320248 39454 320568 39486
rect 320248 39218 320290 39454
rect 320526 39218 320568 39454
rect 320248 39134 320568 39218
rect 320248 38898 320290 39134
rect 320526 38898 320568 39134
rect 320248 38866 320568 38898
rect 330488 39454 330808 39486
rect 330488 39218 330530 39454
rect 330766 39218 330808 39454
rect 330488 39134 330808 39218
rect 330488 38898 330530 39134
rect 330766 38898 330808 39134
rect 330488 38866 330808 38898
rect 340728 39454 341048 39486
rect 340728 39218 340770 39454
rect 341006 39218 341048 39454
rect 340728 39134 341048 39218
rect 340728 38898 340770 39134
rect 341006 38898 341048 39134
rect 340728 38866 341048 38898
rect 350968 39454 351288 39486
rect 350968 39218 351010 39454
rect 351246 39218 351288 39454
rect 350968 39134 351288 39218
rect 350968 38898 351010 39134
rect 351246 38898 351288 39134
rect 350968 38866 351288 38898
rect 361208 39454 361528 39486
rect 361208 39218 361250 39454
rect 361486 39218 361528 39454
rect 361208 39134 361528 39218
rect 361208 38898 361250 39134
rect 361486 38898 361528 39134
rect 361208 38866 361528 38898
rect 371448 39454 371768 39486
rect 371448 39218 371490 39454
rect 371726 39218 371768 39454
rect 371448 39134 371768 39218
rect 371448 38898 371490 39134
rect 371726 38898 371768 39134
rect 371448 38866 371768 38898
rect 381688 39454 382008 39486
rect 381688 39218 381730 39454
rect 381966 39218 382008 39454
rect 381688 39134 382008 39218
rect 381688 38898 381730 39134
rect 381966 38898 382008 39134
rect 381688 38866 382008 38898
rect 391928 39454 392248 39486
rect 391928 39218 391970 39454
rect 392206 39218 392248 39454
rect 391928 39134 392248 39218
rect 391928 38898 391970 39134
rect 392206 38898 392248 39134
rect 391928 38866 392248 38898
rect 402168 39454 402488 39486
rect 402168 39218 402210 39454
rect 402446 39218 402488 39454
rect 402168 39134 402488 39218
rect 402168 38898 402210 39134
rect 402446 38898 402488 39134
rect 402168 38866 402488 38898
rect 412408 39454 412728 39486
rect 412408 39218 412450 39454
rect 412686 39218 412728 39454
rect 412408 39134 412728 39218
rect 412408 38898 412450 39134
rect 412686 38898 412728 39134
rect 412408 38866 412728 38898
rect 422648 39454 422968 39486
rect 422648 39218 422690 39454
rect 422926 39218 422968 39454
rect 422648 39134 422968 39218
rect 422648 38898 422690 39134
rect 422926 38898 422968 39134
rect 422648 38866 422968 38898
rect 432888 39454 433208 39486
rect 432888 39218 432930 39454
rect 433166 39218 433208 39454
rect 432888 39134 433208 39218
rect 432888 38898 432930 39134
rect 433166 38898 433208 39134
rect 432888 38866 433208 38898
rect 443128 39454 443448 39486
rect 443128 39218 443170 39454
rect 443406 39218 443448 39454
rect 443128 39134 443448 39218
rect 443128 38898 443170 39134
rect 443406 38898 443448 39134
rect 443128 38866 443448 38898
rect 453368 39454 453688 39486
rect 453368 39218 453410 39454
rect 453646 39218 453688 39454
rect 453368 39134 453688 39218
rect 453368 38898 453410 39134
rect 453646 38898 453688 39134
rect 453368 38866 453688 38898
rect 463608 39454 463928 39486
rect 463608 39218 463650 39454
rect 463886 39218 463928 39454
rect 463608 39134 463928 39218
rect 463608 38898 463650 39134
rect 463886 38898 463928 39134
rect 463608 38866 463928 38898
rect 473848 39454 474168 39486
rect 473848 39218 473890 39454
rect 474126 39218 474168 39454
rect 473848 39134 474168 39218
rect 473848 38898 473890 39134
rect 474126 38898 474168 39134
rect 473848 38866 474168 38898
rect 484088 39454 484408 39486
rect 484088 39218 484130 39454
rect 484366 39218 484408 39454
rect 484088 39134 484408 39218
rect 484088 38898 484130 39134
rect 484366 38898 484408 39134
rect 484088 38866 484408 38898
rect 494328 39454 494648 39486
rect 494328 39218 494370 39454
rect 494606 39218 494648 39454
rect 494328 39134 494648 39218
rect 494328 38898 494370 39134
rect 494606 38898 494648 39134
rect 494328 38866 494648 38898
rect 504568 39454 504888 39486
rect 504568 39218 504610 39454
rect 504846 39218 504888 39454
rect 504568 39134 504888 39218
rect 504568 38898 504610 39134
rect 504846 38898 504888 39134
rect 504568 38866 504888 38898
rect 514808 39454 515128 39486
rect 514808 39218 514850 39454
rect 515086 39218 515128 39454
rect 514808 39134 515128 39218
rect 514808 38898 514850 39134
rect 515086 38898 515128 39134
rect 514808 38866 515128 38898
rect 525048 39454 525368 39486
rect 525048 39218 525090 39454
rect 525326 39218 525368 39454
rect 525048 39134 525368 39218
rect 525048 38898 525090 39134
rect 525326 38898 525368 39134
rect 525048 38866 525368 38898
rect 535288 39454 535608 39486
rect 535288 39218 535330 39454
rect 535566 39218 535608 39454
rect 535288 39134 535608 39218
rect 535288 38898 535330 39134
rect 535566 38898 535608 39134
rect 535288 38866 535608 38898
rect 28408 21454 28728 21486
rect 28408 21218 28450 21454
rect 28686 21218 28728 21454
rect 28408 21134 28728 21218
rect 28408 20898 28450 21134
rect 28686 20898 28728 21134
rect 28408 20866 28728 20898
rect 38648 21454 38968 21486
rect 38648 21218 38690 21454
rect 38926 21218 38968 21454
rect 38648 21134 38968 21218
rect 38648 20898 38690 21134
rect 38926 20898 38968 21134
rect 38648 20866 38968 20898
rect 48888 21454 49208 21486
rect 48888 21218 48930 21454
rect 49166 21218 49208 21454
rect 48888 21134 49208 21218
rect 48888 20898 48930 21134
rect 49166 20898 49208 21134
rect 48888 20866 49208 20898
rect 59128 21454 59448 21486
rect 59128 21218 59170 21454
rect 59406 21218 59448 21454
rect 59128 21134 59448 21218
rect 59128 20898 59170 21134
rect 59406 20898 59448 21134
rect 59128 20866 59448 20898
rect 69368 21454 69688 21486
rect 69368 21218 69410 21454
rect 69646 21218 69688 21454
rect 69368 21134 69688 21218
rect 69368 20898 69410 21134
rect 69646 20898 69688 21134
rect 69368 20866 69688 20898
rect 79608 21454 79928 21486
rect 79608 21218 79650 21454
rect 79886 21218 79928 21454
rect 79608 21134 79928 21218
rect 79608 20898 79650 21134
rect 79886 20898 79928 21134
rect 79608 20866 79928 20898
rect 89848 21454 90168 21486
rect 89848 21218 89890 21454
rect 90126 21218 90168 21454
rect 89848 21134 90168 21218
rect 89848 20898 89890 21134
rect 90126 20898 90168 21134
rect 89848 20866 90168 20898
rect 100088 21454 100408 21486
rect 100088 21218 100130 21454
rect 100366 21218 100408 21454
rect 100088 21134 100408 21218
rect 100088 20898 100130 21134
rect 100366 20898 100408 21134
rect 100088 20866 100408 20898
rect 110328 21454 110648 21486
rect 110328 21218 110370 21454
rect 110606 21218 110648 21454
rect 110328 21134 110648 21218
rect 110328 20898 110370 21134
rect 110606 20898 110648 21134
rect 110328 20866 110648 20898
rect 120568 21454 120888 21486
rect 120568 21218 120610 21454
rect 120846 21218 120888 21454
rect 120568 21134 120888 21218
rect 120568 20898 120610 21134
rect 120846 20898 120888 21134
rect 120568 20866 120888 20898
rect 130808 21454 131128 21486
rect 130808 21218 130850 21454
rect 131086 21218 131128 21454
rect 130808 21134 131128 21218
rect 130808 20898 130850 21134
rect 131086 20898 131128 21134
rect 130808 20866 131128 20898
rect 141048 21454 141368 21486
rect 141048 21218 141090 21454
rect 141326 21218 141368 21454
rect 141048 21134 141368 21218
rect 141048 20898 141090 21134
rect 141326 20898 141368 21134
rect 141048 20866 141368 20898
rect 151288 21454 151608 21486
rect 151288 21218 151330 21454
rect 151566 21218 151608 21454
rect 151288 21134 151608 21218
rect 151288 20898 151330 21134
rect 151566 20898 151608 21134
rect 151288 20866 151608 20898
rect 161528 21454 161848 21486
rect 161528 21218 161570 21454
rect 161806 21218 161848 21454
rect 161528 21134 161848 21218
rect 161528 20898 161570 21134
rect 161806 20898 161848 21134
rect 161528 20866 161848 20898
rect 171768 21454 172088 21486
rect 171768 21218 171810 21454
rect 172046 21218 172088 21454
rect 171768 21134 172088 21218
rect 171768 20898 171810 21134
rect 172046 20898 172088 21134
rect 171768 20866 172088 20898
rect 182008 21454 182328 21486
rect 182008 21218 182050 21454
rect 182286 21218 182328 21454
rect 182008 21134 182328 21218
rect 182008 20898 182050 21134
rect 182286 20898 182328 21134
rect 182008 20866 182328 20898
rect 192248 21454 192568 21486
rect 192248 21218 192290 21454
rect 192526 21218 192568 21454
rect 192248 21134 192568 21218
rect 192248 20898 192290 21134
rect 192526 20898 192568 21134
rect 192248 20866 192568 20898
rect 202488 21454 202808 21486
rect 202488 21218 202530 21454
rect 202766 21218 202808 21454
rect 202488 21134 202808 21218
rect 202488 20898 202530 21134
rect 202766 20898 202808 21134
rect 202488 20866 202808 20898
rect 212728 21454 213048 21486
rect 212728 21218 212770 21454
rect 213006 21218 213048 21454
rect 212728 21134 213048 21218
rect 212728 20898 212770 21134
rect 213006 20898 213048 21134
rect 212728 20866 213048 20898
rect 222968 21454 223288 21486
rect 222968 21218 223010 21454
rect 223246 21218 223288 21454
rect 222968 21134 223288 21218
rect 222968 20898 223010 21134
rect 223246 20898 223288 21134
rect 222968 20866 223288 20898
rect 233208 21454 233528 21486
rect 233208 21218 233250 21454
rect 233486 21218 233528 21454
rect 233208 21134 233528 21218
rect 233208 20898 233250 21134
rect 233486 20898 233528 21134
rect 233208 20866 233528 20898
rect 243448 21454 243768 21486
rect 243448 21218 243490 21454
rect 243726 21218 243768 21454
rect 243448 21134 243768 21218
rect 243448 20898 243490 21134
rect 243726 20898 243768 21134
rect 243448 20866 243768 20898
rect 253688 21454 254008 21486
rect 253688 21218 253730 21454
rect 253966 21218 254008 21454
rect 253688 21134 254008 21218
rect 253688 20898 253730 21134
rect 253966 20898 254008 21134
rect 253688 20866 254008 20898
rect 263928 21454 264248 21486
rect 263928 21218 263970 21454
rect 264206 21218 264248 21454
rect 263928 21134 264248 21218
rect 263928 20898 263970 21134
rect 264206 20898 264248 21134
rect 263928 20866 264248 20898
rect 274168 21454 274488 21486
rect 274168 21218 274210 21454
rect 274446 21218 274488 21454
rect 274168 21134 274488 21218
rect 274168 20898 274210 21134
rect 274446 20898 274488 21134
rect 274168 20866 274488 20898
rect 284408 21454 284728 21486
rect 284408 21218 284450 21454
rect 284686 21218 284728 21454
rect 284408 21134 284728 21218
rect 284408 20898 284450 21134
rect 284686 20898 284728 21134
rect 284408 20866 284728 20898
rect 294648 21454 294968 21486
rect 294648 21218 294690 21454
rect 294926 21218 294968 21454
rect 294648 21134 294968 21218
rect 294648 20898 294690 21134
rect 294926 20898 294968 21134
rect 294648 20866 294968 20898
rect 304888 21454 305208 21486
rect 304888 21218 304930 21454
rect 305166 21218 305208 21454
rect 304888 21134 305208 21218
rect 304888 20898 304930 21134
rect 305166 20898 305208 21134
rect 304888 20866 305208 20898
rect 315128 21454 315448 21486
rect 315128 21218 315170 21454
rect 315406 21218 315448 21454
rect 315128 21134 315448 21218
rect 315128 20898 315170 21134
rect 315406 20898 315448 21134
rect 315128 20866 315448 20898
rect 325368 21454 325688 21486
rect 325368 21218 325410 21454
rect 325646 21218 325688 21454
rect 325368 21134 325688 21218
rect 325368 20898 325410 21134
rect 325646 20898 325688 21134
rect 325368 20866 325688 20898
rect 335608 21454 335928 21486
rect 335608 21218 335650 21454
rect 335886 21218 335928 21454
rect 335608 21134 335928 21218
rect 335608 20898 335650 21134
rect 335886 20898 335928 21134
rect 335608 20866 335928 20898
rect 345848 21454 346168 21486
rect 345848 21218 345890 21454
rect 346126 21218 346168 21454
rect 345848 21134 346168 21218
rect 345848 20898 345890 21134
rect 346126 20898 346168 21134
rect 345848 20866 346168 20898
rect 356088 21454 356408 21486
rect 356088 21218 356130 21454
rect 356366 21218 356408 21454
rect 356088 21134 356408 21218
rect 356088 20898 356130 21134
rect 356366 20898 356408 21134
rect 356088 20866 356408 20898
rect 366328 21454 366648 21486
rect 366328 21218 366370 21454
rect 366606 21218 366648 21454
rect 366328 21134 366648 21218
rect 366328 20898 366370 21134
rect 366606 20898 366648 21134
rect 366328 20866 366648 20898
rect 376568 21454 376888 21486
rect 376568 21218 376610 21454
rect 376846 21218 376888 21454
rect 376568 21134 376888 21218
rect 376568 20898 376610 21134
rect 376846 20898 376888 21134
rect 376568 20866 376888 20898
rect 386808 21454 387128 21486
rect 386808 21218 386850 21454
rect 387086 21218 387128 21454
rect 386808 21134 387128 21218
rect 386808 20898 386850 21134
rect 387086 20898 387128 21134
rect 386808 20866 387128 20898
rect 397048 21454 397368 21486
rect 397048 21218 397090 21454
rect 397326 21218 397368 21454
rect 397048 21134 397368 21218
rect 397048 20898 397090 21134
rect 397326 20898 397368 21134
rect 397048 20866 397368 20898
rect 407288 21454 407608 21486
rect 407288 21218 407330 21454
rect 407566 21218 407608 21454
rect 407288 21134 407608 21218
rect 407288 20898 407330 21134
rect 407566 20898 407608 21134
rect 407288 20866 407608 20898
rect 417528 21454 417848 21486
rect 417528 21218 417570 21454
rect 417806 21218 417848 21454
rect 417528 21134 417848 21218
rect 417528 20898 417570 21134
rect 417806 20898 417848 21134
rect 417528 20866 417848 20898
rect 427768 21454 428088 21486
rect 427768 21218 427810 21454
rect 428046 21218 428088 21454
rect 427768 21134 428088 21218
rect 427768 20898 427810 21134
rect 428046 20898 428088 21134
rect 427768 20866 428088 20898
rect 438008 21454 438328 21486
rect 438008 21218 438050 21454
rect 438286 21218 438328 21454
rect 438008 21134 438328 21218
rect 438008 20898 438050 21134
rect 438286 20898 438328 21134
rect 438008 20866 438328 20898
rect 448248 21454 448568 21486
rect 448248 21218 448290 21454
rect 448526 21218 448568 21454
rect 448248 21134 448568 21218
rect 448248 20898 448290 21134
rect 448526 20898 448568 21134
rect 448248 20866 448568 20898
rect 458488 21454 458808 21486
rect 458488 21218 458530 21454
rect 458766 21218 458808 21454
rect 458488 21134 458808 21218
rect 458488 20898 458530 21134
rect 458766 20898 458808 21134
rect 458488 20866 458808 20898
rect 468728 21454 469048 21486
rect 468728 21218 468770 21454
rect 469006 21218 469048 21454
rect 468728 21134 469048 21218
rect 468728 20898 468770 21134
rect 469006 20898 469048 21134
rect 468728 20866 469048 20898
rect 478968 21454 479288 21486
rect 478968 21218 479010 21454
rect 479246 21218 479288 21454
rect 478968 21134 479288 21218
rect 478968 20898 479010 21134
rect 479246 20898 479288 21134
rect 478968 20866 479288 20898
rect 489208 21454 489528 21486
rect 489208 21218 489250 21454
rect 489486 21218 489528 21454
rect 489208 21134 489528 21218
rect 489208 20898 489250 21134
rect 489486 20898 489528 21134
rect 489208 20866 489528 20898
rect 499448 21454 499768 21486
rect 499448 21218 499490 21454
rect 499726 21218 499768 21454
rect 499448 21134 499768 21218
rect 499448 20898 499490 21134
rect 499726 20898 499768 21134
rect 499448 20866 499768 20898
rect 509688 21454 510008 21486
rect 509688 21218 509730 21454
rect 509966 21218 510008 21454
rect 509688 21134 510008 21218
rect 509688 20898 509730 21134
rect 509966 20898 510008 21134
rect 509688 20866 510008 20898
rect 519928 21454 520248 21486
rect 519928 21218 519970 21454
rect 520206 21218 520248 21454
rect 519928 21134 520248 21218
rect 519928 20898 519970 21134
rect 520206 20898 520248 21134
rect 519928 20866 520248 20898
rect 530168 21454 530488 21486
rect 530168 21218 530210 21454
rect 530446 21218 530488 21454
rect 530168 21134 530488 21218
rect 530168 20898 530210 21134
rect 530446 20898 530488 21134
rect 530168 20866 530488 20898
rect 15754 6938 15786 7174
rect 16022 6938 16106 7174
rect 16342 6938 16374 7174
rect 15754 6854 16374 6938
rect 15754 6618 15786 6854
rect 16022 6618 16106 6854
rect 16342 6618 16374 6854
rect 15754 -2266 16374 6618
rect 17154 -1306 17774 13000
rect 17154 -1542 17186 -1306
rect 17422 -1542 17506 -1306
rect 17742 -1542 17774 -1306
rect 17154 -1626 17774 -1542
rect 17154 -1862 17186 -1626
rect 17422 -1862 17506 -1626
rect 17742 -1862 17774 -1626
rect 17154 -1894 17774 -1862
rect 15754 -2502 15786 -2266
rect 16022 -2502 16106 -2266
rect 16342 -2502 16374 -2266
rect 15754 -2586 16374 -2502
rect 15754 -2822 15786 -2586
rect 16022 -2822 16106 -2586
rect 16342 -2822 16374 -2586
rect 15754 -3814 16374 -2822
rect 14354 -5382 14386 -5146
rect 14622 -5382 14706 -5146
rect 14942 -5382 14974 -5146
rect 14354 -5466 14974 -5382
rect 14354 -5702 14386 -5466
rect 14622 -5702 14706 -5466
rect 14942 -5702 14974 -5466
rect 14354 -5734 14974 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 18074 -7066 18694 13000
rect 19474 10894 20094 13000
rect 19474 10658 19506 10894
rect 19742 10658 19826 10894
rect 20062 10658 20094 10894
rect 19474 10574 20094 10658
rect 19474 10338 19506 10574
rect 19742 10338 19826 10574
rect 20062 10338 20094 10574
rect 19474 -4186 20094 10338
rect 20874 -3226 21494 13000
rect 22274 3454 22894 13000
rect 22274 3218 22306 3454
rect 22542 3218 22626 3454
rect 22862 3218 22894 3454
rect 22274 3134 22894 3218
rect 22274 2898 22306 3134
rect 22542 2898 22626 3134
rect 22862 2898 22894 3134
rect 22274 -346 22894 2898
rect 22274 -582 22306 -346
rect 22542 -582 22626 -346
rect 22862 -582 22894 -346
rect 22274 -666 22894 -582
rect 22274 -902 22306 -666
rect 22542 -902 22626 -666
rect 22862 -902 22894 -666
rect 22274 -1894 22894 -902
rect 20874 -3462 20906 -3226
rect 21142 -3462 21226 -3226
rect 21462 -3462 21494 -3226
rect 20874 -3546 21494 -3462
rect 20874 -3782 20906 -3546
rect 21142 -3782 21226 -3546
rect 21462 -3782 21494 -3546
rect 20874 -3814 21494 -3782
rect 19474 -4422 19506 -4186
rect 19742 -4422 19826 -4186
rect 20062 -4422 20094 -4186
rect 19474 -4506 20094 -4422
rect 19474 -4742 19506 -4506
rect 19742 -4742 19826 -4506
rect 20062 -4742 20094 -4506
rect 19474 -5734 20094 -4742
rect 18074 -7302 18106 -7066
rect 18342 -7302 18426 -7066
rect 18662 -7302 18694 -7066
rect 18074 -7386 18694 -7302
rect 18074 -7622 18106 -7386
rect 18342 -7622 18426 -7386
rect 18662 -7622 18694 -7386
rect 18074 -7654 18694 -7622
rect 23194 -6106 23814 13000
rect 24594 -5146 25214 13000
rect 25994 7174 26614 13000
rect 25994 6938 26026 7174
rect 26262 6938 26346 7174
rect 26582 6938 26614 7174
rect 25994 6854 26614 6938
rect 25994 6618 26026 6854
rect 26262 6618 26346 6854
rect 26582 6618 26614 6854
rect 25994 -2266 26614 6618
rect 27394 -1306 28014 13000
rect 27394 -1542 27426 -1306
rect 27662 -1542 27746 -1306
rect 27982 -1542 28014 -1306
rect 27394 -1626 28014 -1542
rect 27394 -1862 27426 -1626
rect 27662 -1862 27746 -1626
rect 27982 -1862 28014 -1626
rect 27394 -1894 28014 -1862
rect 25994 -2502 26026 -2266
rect 26262 -2502 26346 -2266
rect 26582 -2502 26614 -2266
rect 25994 -2586 26614 -2502
rect 25994 -2822 26026 -2586
rect 26262 -2822 26346 -2586
rect 26582 -2822 26614 -2586
rect 25994 -3814 26614 -2822
rect 24594 -5382 24626 -5146
rect 24862 -5382 24946 -5146
rect 25182 -5382 25214 -5146
rect 24594 -5466 25214 -5382
rect 24594 -5702 24626 -5466
rect 24862 -5702 24946 -5466
rect 25182 -5702 25214 -5466
rect 24594 -5734 25214 -5702
rect 23194 -6342 23226 -6106
rect 23462 -6342 23546 -6106
rect 23782 -6342 23814 -6106
rect 23194 -6426 23814 -6342
rect 23194 -6662 23226 -6426
rect 23462 -6662 23546 -6426
rect 23782 -6662 23814 -6426
rect 23194 -7654 23814 -6662
rect 28314 -7066 28934 13000
rect 29714 10894 30334 13000
rect 29714 10658 29746 10894
rect 29982 10658 30066 10894
rect 30302 10658 30334 10894
rect 29714 10574 30334 10658
rect 29714 10338 29746 10574
rect 29982 10338 30066 10574
rect 30302 10338 30334 10574
rect 29714 -4186 30334 10338
rect 31114 -3226 31734 13000
rect 32514 3454 33134 13000
rect 32514 3218 32546 3454
rect 32782 3218 32866 3454
rect 33102 3218 33134 3454
rect 32514 3134 33134 3218
rect 32514 2898 32546 3134
rect 32782 2898 32866 3134
rect 33102 2898 33134 3134
rect 32514 -346 33134 2898
rect 32514 -582 32546 -346
rect 32782 -582 32866 -346
rect 33102 -582 33134 -346
rect 32514 -666 33134 -582
rect 32514 -902 32546 -666
rect 32782 -902 32866 -666
rect 33102 -902 33134 -666
rect 32514 -1894 33134 -902
rect 31114 -3462 31146 -3226
rect 31382 -3462 31466 -3226
rect 31702 -3462 31734 -3226
rect 31114 -3546 31734 -3462
rect 31114 -3782 31146 -3546
rect 31382 -3782 31466 -3546
rect 31702 -3782 31734 -3546
rect 31114 -3814 31734 -3782
rect 29714 -4422 29746 -4186
rect 29982 -4422 30066 -4186
rect 30302 -4422 30334 -4186
rect 29714 -4506 30334 -4422
rect 29714 -4742 29746 -4506
rect 29982 -4742 30066 -4506
rect 30302 -4742 30334 -4506
rect 29714 -5734 30334 -4742
rect 28314 -7302 28346 -7066
rect 28582 -7302 28666 -7066
rect 28902 -7302 28934 -7066
rect 28314 -7386 28934 -7302
rect 28314 -7622 28346 -7386
rect 28582 -7622 28666 -7386
rect 28902 -7622 28934 -7386
rect 28314 -7654 28934 -7622
rect 33434 -6106 34054 13000
rect 34834 -5146 35454 13000
rect 36234 7174 36854 13000
rect 36234 6938 36266 7174
rect 36502 6938 36586 7174
rect 36822 6938 36854 7174
rect 36234 6854 36854 6938
rect 36234 6618 36266 6854
rect 36502 6618 36586 6854
rect 36822 6618 36854 6854
rect 36234 -2266 36854 6618
rect 37634 -1306 38254 13000
rect 37634 -1542 37666 -1306
rect 37902 -1542 37986 -1306
rect 38222 -1542 38254 -1306
rect 37634 -1626 38254 -1542
rect 37634 -1862 37666 -1626
rect 37902 -1862 37986 -1626
rect 38222 -1862 38254 -1626
rect 37634 -1894 38254 -1862
rect 36234 -2502 36266 -2266
rect 36502 -2502 36586 -2266
rect 36822 -2502 36854 -2266
rect 36234 -2586 36854 -2502
rect 36234 -2822 36266 -2586
rect 36502 -2822 36586 -2586
rect 36822 -2822 36854 -2586
rect 36234 -3814 36854 -2822
rect 34834 -5382 34866 -5146
rect 35102 -5382 35186 -5146
rect 35422 -5382 35454 -5146
rect 34834 -5466 35454 -5382
rect 34834 -5702 34866 -5466
rect 35102 -5702 35186 -5466
rect 35422 -5702 35454 -5466
rect 34834 -5734 35454 -5702
rect 33434 -6342 33466 -6106
rect 33702 -6342 33786 -6106
rect 34022 -6342 34054 -6106
rect 33434 -6426 34054 -6342
rect 33434 -6662 33466 -6426
rect 33702 -6662 33786 -6426
rect 34022 -6662 34054 -6426
rect 33434 -7654 34054 -6662
rect 38554 -7066 39174 13000
rect 39954 10894 40574 13000
rect 39954 10658 39986 10894
rect 40222 10658 40306 10894
rect 40542 10658 40574 10894
rect 39954 10574 40574 10658
rect 39954 10338 39986 10574
rect 40222 10338 40306 10574
rect 40542 10338 40574 10574
rect 39954 -4186 40574 10338
rect 41354 -3226 41974 13000
rect 42754 3454 43374 13000
rect 42754 3218 42786 3454
rect 43022 3218 43106 3454
rect 43342 3218 43374 3454
rect 42754 3134 43374 3218
rect 42754 2898 42786 3134
rect 43022 2898 43106 3134
rect 43342 2898 43374 3134
rect 42754 -346 43374 2898
rect 42754 -582 42786 -346
rect 43022 -582 43106 -346
rect 43342 -582 43374 -346
rect 42754 -666 43374 -582
rect 42754 -902 42786 -666
rect 43022 -902 43106 -666
rect 43342 -902 43374 -666
rect 42754 -1894 43374 -902
rect 41354 -3462 41386 -3226
rect 41622 -3462 41706 -3226
rect 41942 -3462 41974 -3226
rect 41354 -3546 41974 -3462
rect 41354 -3782 41386 -3546
rect 41622 -3782 41706 -3546
rect 41942 -3782 41974 -3546
rect 41354 -3814 41974 -3782
rect 39954 -4422 39986 -4186
rect 40222 -4422 40306 -4186
rect 40542 -4422 40574 -4186
rect 39954 -4506 40574 -4422
rect 39954 -4742 39986 -4506
rect 40222 -4742 40306 -4506
rect 40542 -4742 40574 -4506
rect 39954 -5734 40574 -4742
rect 38554 -7302 38586 -7066
rect 38822 -7302 38906 -7066
rect 39142 -7302 39174 -7066
rect 38554 -7386 39174 -7302
rect 38554 -7622 38586 -7386
rect 38822 -7622 38906 -7386
rect 39142 -7622 39174 -7386
rect 38554 -7654 39174 -7622
rect 43674 -6106 44294 13000
rect 45074 -5146 45694 13000
rect 46474 7174 47094 13000
rect 46474 6938 46506 7174
rect 46742 6938 46826 7174
rect 47062 6938 47094 7174
rect 46474 6854 47094 6938
rect 46474 6618 46506 6854
rect 46742 6618 46826 6854
rect 47062 6618 47094 6854
rect 46474 -2266 47094 6618
rect 47874 -1306 48494 13000
rect 47874 -1542 47906 -1306
rect 48142 -1542 48226 -1306
rect 48462 -1542 48494 -1306
rect 47874 -1626 48494 -1542
rect 47874 -1862 47906 -1626
rect 48142 -1862 48226 -1626
rect 48462 -1862 48494 -1626
rect 47874 -1894 48494 -1862
rect 46474 -2502 46506 -2266
rect 46742 -2502 46826 -2266
rect 47062 -2502 47094 -2266
rect 46474 -2586 47094 -2502
rect 46474 -2822 46506 -2586
rect 46742 -2822 46826 -2586
rect 47062 -2822 47094 -2586
rect 46474 -3814 47094 -2822
rect 45074 -5382 45106 -5146
rect 45342 -5382 45426 -5146
rect 45662 -5382 45694 -5146
rect 45074 -5466 45694 -5382
rect 45074 -5702 45106 -5466
rect 45342 -5702 45426 -5466
rect 45662 -5702 45694 -5466
rect 45074 -5734 45694 -5702
rect 43674 -6342 43706 -6106
rect 43942 -6342 44026 -6106
rect 44262 -6342 44294 -6106
rect 43674 -6426 44294 -6342
rect 43674 -6662 43706 -6426
rect 43942 -6662 44026 -6426
rect 44262 -6662 44294 -6426
rect 43674 -7654 44294 -6662
rect 48794 -7066 49414 13000
rect 50194 10894 50814 13000
rect 50194 10658 50226 10894
rect 50462 10658 50546 10894
rect 50782 10658 50814 10894
rect 50194 10574 50814 10658
rect 50194 10338 50226 10574
rect 50462 10338 50546 10574
rect 50782 10338 50814 10574
rect 50194 -4186 50814 10338
rect 51594 -3226 52214 13000
rect 52994 3454 53614 13000
rect 52994 3218 53026 3454
rect 53262 3218 53346 3454
rect 53582 3218 53614 3454
rect 52994 3134 53614 3218
rect 52994 2898 53026 3134
rect 53262 2898 53346 3134
rect 53582 2898 53614 3134
rect 52994 -346 53614 2898
rect 52994 -582 53026 -346
rect 53262 -582 53346 -346
rect 53582 -582 53614 -346
rect 52994 -666 53614 -582
rect 52994 -902 53026 -666
rect 53262 -902 53346 -666
rect 53582 -902 53614 -666
rect 52994 -1894 53614 -902
rect 51594 -3462 51626 -3226
rect 51862 -3462 51946 -3226
rect 52182 -3462 52214 -3226
rect 51594 -3546 52214 -3462
rect 51594 -3782 51626 -3546
rect 51862 -3782 51946 -3546
rect 52182 -3782 52214 -3546
rect 51594 -3814 52214 -3782
rect 50194 -4422 50226 -4186
rect 50462 -4422 50546 -4186
rect 50782 -4422 50814 -4186
rect 50194 -4506 50814 -4422
rect 50194 -4742 50226 -4506
rect 50462 -4742 50546 -4506
rect 50782 -4742 50814 -4506
rect 50194 -5734 50814 -4742
rect 48794 -7302 48826 -7066
rect 49062 -7302 49146 -7066
rect 49382 -7302 49414 -7066
rect 48794 -7386 49414 -7302
rect 48794 -7622 48826 -7386
rect 49062 -7622 49146 -7386
rect 49382 -7622 49414 -7386
rect 48794 -7654 49414 -7622
rect 53914 -6106 54534 13000
rect 55314 -5146 55934 13000
rect 56714 7174 57334 13000
rect 56714 6938 56746 7174
rect 56982 6938 57066 7174
rect 57302 6938 57334 7174
rect 56714 6854 57334 6938
rect 56714 6618 56746 6854
rect 56982 6618 57066 6854
rect 57302 6618 57334 6854
rect 56714 -2266 57334 6618
rect 58114 -1306 58734 13000
rect 58114 -1542 58146 -1306
rect 58382 -1542 58466 -1306
rect 58702 -1542 58734 -1306
rect 58114 -1626 58734 -1542
rect 58114 -1862 58146 -1626
rect 58382 -1862 58466 -1626
rect 58702 -1862 58734 -1626
rect 58114 -1894 58734 -1862
rect 56714 -2502 56746 -2266
rect 56982 -2502 57066 -2266
rect 57302 -2502 57334 -2266
rect 56714 -2586 57334 -2502
rect 56714 -2822 56746 -2586
rect 56982 -2822 57066 -2586
rect 57302 -2822 57334 -2586
rect 56714 -3814 57334 -2822
rect 55314 -5382 55346 -5146
rect 55582 -5382 55666 -5146
rect 55902 -5382 55934 -5146
rect 55314 -5466 55934 -5382
rect 55314 -5702 55346 -5466
rect 55582 -5702 55666 -5466
rect 55902 -5702 55934 -5466
rect 55314 -5734 55934 -5702
rect 53914 -6342 53946 -6106
rect 54182 -6342 54266 -6106
rect 54502 -6342 54534 -6106
rect 53914 -6426 54534 -6342
rect 53914 -6662 53946 -6426
rect 54182 -6662 54266 -6426
rect 54502 -6662 54534 -6426
rect 53914 -7654 54534 -6662
rect 59034 -7066 59654 13000
rect 60434 10894 61054 13000
rect 60434 10658 60466 10894
rect 60702 10658 60786 10894
rect 61022 10658 61054 10894
rect 60434 10574 61054 10658
rect 60434 10338 60466 10574
rect 60702 10338 60786 10574
rect 61022 10338 61054 10574
rect 60434 -4186 61054 10338
rect 61834 -3226 62454 13000
rect 63234 3454 63854 13000
rect 63234 3218 63266 3454
rect 63502 3218 63586 3454
rect 63822 3218 63854 3454
rect 63234 3134 63854 3218
rect 63234 2898 63266 3134
rect 63502 2898 63586 3134
rect 63822 2898 63854 3134
rect 63234 -346 63854 2898
rect 63234 -582 63266 -346
rect 63502 -582 63586 -346
rect 63822 -582 63854 -346
rect 63234 -666 63854 -582
rect 63234 -902 63266 -666
rect 63502 -902 63586 -666
rect 63822 -902 63854 -666
rect 63234 -1894 63854 -902
rect 61834 -3462 61866 -3226
rect 62102 -3462 62186 -3226
rect 62422 -3462 62454 -3226
rect 61834 -3546 62454 -3462
rect 61834 -3782 61866 -3546
rect 62102 -3782 62186 -3546
rect 62422 -3782 62454 -3546
rect 61834 -3814 62454 -3782
rect 60434 -4422 60466 -4186
rect 60702 -4422 60786 -4186
rect 61022 -4422 61054 -4186
rect 60434 -4506 61054 -4422
rect 60434 -4742 60466 -4506
rect 60702 -4742 60786 -4506
rect 61022 -4742 61054 -4506
rect 60434 -5734 61054 -4742
rect 59034 -7302 59066 -7066
rect 59302 -7302 59386 -7066
rect 59622 -7302 59654 -7066
rect 59034 -7386 59654 -7302
rect 59034 -7622 59066 -7386
rect 59302 -7622 59386 -7386
rect 59622 -7622 59654 -7386
rect 59034 -7654 59654 -7622
rect 64154 -6106 64774 13000
rect 65554 -5146 66174 13000
rect 66954 7174 67574 13000
rect 66954 6938 66986 7174
rect 67222 6938 67306 7174
rect 67542 6938 67574 7174
rect 66954 6854 67574 6938
rect 66954 6618 66986 6854
rect 67222 6618 67306 6854
rect 67542 6618 67574 6854
rect 66954 -2266 67574 6618
rect 68354 -1306 68974 13000
rect 68354 -1542 68386 -1306
rect 68622 -1542 68706 -1306
rect 68942 -1542 68974 -1306
rect 68354 -1626 68974 -1542
rect 68354 -1862 68386 -1626
rect 68622 -1862 68706 -1626
rect 68942 -1862 68974 -1626
rect 68354 -1894 68974 -1862
rect 66954 -2502 66986 -2266
rect 67222 -2502 67306 -2266
rect 67542 -2502 67574 -2266
rect 66954 -2586 67574 -2502
rect 66954 -2822 66986 -2586
rect 67222 -2822 67306 -2586
rect 67542 -2822 67574 -2586
rect 66954 -3814 67574 -2822
rect 65554 -5382 65586 -5146
rect 65822 -5382 65906 -5146
rect 66142 -5382 66174 -5146
rect 65554 -5466 66174 -5382
rect 65554 -5702 65586 -5466
rect 65822 -5702 65906 -5466
rect 66142 -5702 66174 -5466
rect 65554 -5734 66174 -5702
rect 64154 -6342 64186 -6106
rect 64422 -6342 64506 -6106
rect 64742 -6342 64774 -6106
rect 64154 -6426 64774 -6342
rect 64154 -6662 64186 -6426
rect 64422 -6662 64506 -6426
rect 64742 -6662 64774 -6426
rect 64154 -7654 64774 -6662
rect 69274 -7066 69894 13000
rect 70674 10894 71294 13000
rect 70674 10658 70706 10894
rect 70942 10658 71026 10894
rect 71262 10658 71294 10894
rect 70674 10574 71294 10658
rect 70674 10338 70706 10574
rect 70942 10338 71026 10574
rect 71262 10338 71294 10574
rect 70674 -4186 71294 10338
rect 72074 -3226 72694 13000
rect 73474 3454 74094 13000
rect 73474 3218 73506 3454
rect 73742 3218 73826 3454
rect 74062 3218 74094 3454
rect 73474 3134 74094 3218
rect 73474 2898 73506 3134
rect 73742 2898 73826 3134
rect 74062 2898 74094 3134
rect 73474 -346 74094 2898
rect 73474 -582 73506 -346
rect 73742 -582 73826 -346
rect 74062 -582 74094 -346
rect 73474 -666 74094 -582
rect 73474 -902 73506 -666
rect 73742 -902 73826 -666
rect 74062 -902 74094 -666
rect 73474 -1894 74094 -902
rect 72074 -3462 72106 -3226
rect 72342 -3462 72426 -3226
rect 72662 -3462 72694 -3226
rect 72074 -3546 72694 -3462
rect 72074 -3782 72106 -3546
rect 72342 -3782 72426 -3546
rect 72662 -3782 72694 -3546
rect 72074 -3814 72694 -3782
rect 70674 -4422 70706 -4186
rect 70942 -4422 71026 -4186
rect 71262 -4422 71294 -4186
rect 70674 -4506 71294 -4422
rect 70674 -4742 70706 -4506
rect 70942 -4742 71026 -4506
rect 71262 -4742 71294 -4506
rect 70674 -5734 71294 -4742
rect 69274 -7302 69306 -7066
rect 69542 -7302 69626 -7066
rect 69862 -7302 69894 -7066
rect 69274 -7386 69894 -7302
rect 69274 -7622 69306 -7386
rect 69542 -7622 69626 -7386
rect 69862 -7622 69894 -7386
rect 69274 -7654 69894 -7622
rect 74394 -6106 75014 13000
rect 75794 -5146 76414 13000
rect 77194 7174 77814 13000
rect 77194 6938 77226 7174
rect 77462 6938 77546 7174
rect 77782 6938 77814 7174
rect 77194 6854 77814 6938
rect 77194 6618 77226 6854
rect 77462 6618 77546 6854
rect 77782 6618 77814 6854
rect 77194 -2266 77814 6618
rect 78594 -1306 79214 13000
rect 78594 -1542 78626 -1306
rect 78862 -1542 78946 -1306
rect 79182 -1542 79214 -1306
rect 78594 -1626 79214 -1542
rect 78594 -1862 78626 -1626
rect 78862 -1862 78946 -1626
rect 79182 -1862 79214 -1626
rect 78594 -1894 79214 -1862
rect 77194 -2502 77226 -2266
rect 77462 -2502 77546 -2266
rect 77782 -2502 77814 -2266
rect 77194 -2586 77814 -2502
rect 77194 -2822 77226 -2586
rect 77462 -2822 77546 -2586
rect 77782 -2822 77814 -2586
rect 77194 -3814 77814 -2822
rect 75794 -5382 75826 -5146
rect 76062 -5382 76146 -5146
rect 76382 -5382 76414 -5146
rect 75794 -5466 76414 -5382
rect 75794 -5702 75826 -5466
rect 76062 -5702 76146 -5466
rect 76382 -5702 76414 -5466
rect 75794 -5734 76414 -5702
rect 74394 -6342 74426 -6106
rect 74662 -6342 74746 -6106
rect 74982 -6342 75014 -6106
rect 74394 -6426 75014 -6342
rect 74394 -6662 74426 -6426
rect 74662 -6662 74746 -6426
rect 74982 -6662 75014 -6426
rect 74394 -7654 75014 -6662
rect 79514 -7066 80134 13000
rect 80914 10894 81534 13000
rect 80914 10658 80946 10894
rect 81182 10658 81266 10894
rect 81502 10658 81534 10894
rect 80914 10574 81534 10658
rect 80914 10338 80946 10574
rect 81182 10338 81266 10574
rect 81502 10338 81534 10574
rect 80914 -4186 81534 10338
rect 82314 -3226 82934 13000
rect 83714 3454 84334 13000
rect 83714 3218 83746 3454
rect 83982 3218 84066 3454
rect 84302 3218 84334 3454
rect 83714 3134 84334 3218
rect 83714 2898 83746 3134
rect 83982 2898 84066 3134
rect 84302 2898 84334 3134
rect 83714 -346 84334 2898
rect 83714 -582 83746 -346
rect 83982 -582 84066 -346
rect 84302 -582 84334 -346
rect 83714 -666 84334 -582
rect 83714 -902 83746 -666
rect 83982 -902 84066 -666
rect 84302 -902 84334 -666
rect 83714 -1894 84334 -902
rect 82314 -3462 82346 -3226
rect 82582 -3462 82666 -3226
rect 82902 -3462 82934 -3226
rect 82314 -3546 82934 -3462
rect 82314 -3782 82346 -3546
rect 82582 -3782 82666 -3546
rect 82902 -3782 82934 -3546
rect 82314 -3814 82934 -3782
rect 80914 -4422 80946 -4186
rect 81182 -4422 81266 -4186
rect 81502 -4422 81534 -4186
rect 80914 -4506 81534 -4422
rect 80914 -4742 80946 -4506
rect 81182 -4742 81266 -4506
rect 81502 -4742 81534 -4506
rect 80914 -5734 81534 -4742
rect 79514 -7302 79546 -7066
rect 79782 -7302 79866 -7066
rect 80102 -7302 80134 -7066
rect 79514 -7386 80134 -7302
rect 79514 -7622 79546 -7386
rect 79782 -7622 79866 -7386
rect 80102 -7622 80134 -7386
rect 79514 -7654 80134 -7622
rect 84634 -6106 85254 13000
rect 86034 -5146 86654 13000
rect 87434 7174 88054 13000
rect 87434 6938 87466 7174
rect 87702 6938 87786 7174
rect 88022 6938 88054 7174
rect 87434 6854 88054 6938
rect 87434 6618 87466 6854
rect 87702 6618 87786 6854
rect 88022 6618 88054 6854
rect 87434 -2266 88054 6618
rect 88834 -1306 89454 13000
rect 88834 -1542 88866 -1306
rect 89102 -1542 89186 -1306
rect 89422 -1542 89454 -1306
rect 88834 -1626 89454 -1542
rect 88834 -1862 88866 -1626
rect 89102 -1862 89186 -1626
rect 89422 -1862 89454 -1626
rect 88834 -1894 89454 -1862
rect 87434 -2502 87466 -2266
rect 87702 -2502 87786 -2266
rect 88022 -2502 88054 -2266
rect 87434 -2586 88054 -2502
rect 87434 -2822 87466 -2586
rect 87702 -2822 87786 -2586
rect 88022 -2822 88054 -2586
rect 87434 -3814 88054 -2822
rect 86034 -5382 86066 -5146
rect 86302 -5382 86386 -5146
rect 86622 -5382 86654 -5146
rect 86034 -5466 86654 -5382
rect 86034 -5702 86066 -5466
rect 86302 -5702 86386 -5466
rect 86622 -5702 86654 -5466
rect 86034 -5734 86654 -5702
rect 84634 -6342 84666 -6106
rect 84902 -6342 84986 -6106
rect 85222 -6342 85254 -6106
rect 84634 -6426 85254 -6342
rect 84634 -6662 84666 -6426
rect 84902 -6662 84986 -6426
rect 85222 -6662 85254 -6426
rect 84634 -7654 85254 -6662
rect 89754 -7066 90374 13000
rect 91154 10894 91774 13000
rect 91154 10658 91186 10894
rect 91422 10658 91506 10894
rect 91742 10658 91774 10894
rect 91154 10574 91774 10658
rect 91154 10338 91186 10574
rect 91422 10338 91506 10574
rect 91742 10338 91774 10574
rect 91154 -4186 91774 10338
rect 92554 -3226 93174 13000
rect 93954 3454 94574 13000
rect 93954 3218 93986 3454
rect 94222 3218 94306 3454
rect 94542 3218 94574 3454
rect 93954 3134 94574 3218
rect 93954 2898 93986 3134
rect 94222 2898 94306 3134
rect 94542 2898 94574 3134
rect 93954 -346 94574 2898
rect 93954 -582 93986 -346
rect 94222 -582 94306 -346
rect 94542 -582 94574 -346
rect 93954 -666 94574 -582
rect 93954 -902 93986 -666
rect 94222 -902 94306 -666
rect 94542 -902 94574 -666
rect 93954 -1894 94574 -902
rect 92554 -3462 92586 -3226
rect 92822 -3462 92906 -3226
rect 93142 -3462 93174 -3226
rect 92554 -3546 93174 -3462
rect 92554 -3782 92586 -3546
rect 92822 -3782 92906 -3546
rect 93142 -3782 93174 -3546
rect 92554 -3814 93174 -3782
rect 91154 -4422 91186 -4186
rect 91422 -4422 91506 -4186
rect 91742 -4422 91774 -4186
rect 91154 -4506 91774 -4422
rect 91154 -4742 91186 -4506
rect 91422 -4742 91506 -4506
rect 91742 -4742 91774 -4506
rect 91154 -5734 91774 -4742
rect 89754 -7302 89786 -7066
rect 90022 -7302 90106 -7066
rect 90342 -7302 90374 -7066
rect 89754 -7386 90374 -7302
rect 89754 -7622 89786 -7386
rect 90022 -7622 90106 -7386
rect 90342 -7622 90374 -7386
rect 89754 -7654 90374 -7622
rect 94874 -6106 95494 13000
rect 96274 -5146 96894 13000
rect 97674 7174 98294 13000
rect 97674 6938 97706 7174
rect 97942 6938 98026 7174
rect 98262 6938 98294 7174
rect 97674 6854 98294 6938
rect 97674 6618 97706 6854
rect 97942 6618 98026 6854
rect 98262 6618 98294 6854
rect 97674 -2266 98294 6618
rect 99074 -1306 99694 13000
rect 99074 -1542 99106 -1306
rect 99342 -1542 99426 -1306
rect 99662 -1542 99694 -1306
rect 99074 -1626 99694 -1542
rect 99074 -1862 99106 -1626
rect 99342 -1862 99426 -1626
rect 99662 -1862 99694 -1626
rect 99074 -1894 99694 -1862
rect 97674 -2502 97706 -2266
rect 97942 -2502 98026 -2266
rect 98262 -2502 98294 -2266
rect 97674 -2586 98294 -2502
rect 97674 -2822 97706 -2586
rect 97942 -2822 98026 -2586
rect 98262 -2822 98294 -2586
rect 97674 -3814 98294 -2822
rect 96274 -5382 96306 -5146
rect 96542 -5382 96626 -5146
rect 96862 -5382 96894 -5146
rect 96274 -5466 96894 -5382
rect 96274 -5702 96306 -5466
rect 96542 -5702 96626 -5466
rect 96862 -5702 96894 -5466
rect 96274 -5734 96894 -5702
rect 94874 -6342 94906 -6106
rect 95142 -6342 95226 -6106
rect 95462 -6342 95494 -6106
rect 94874 -6426 95494 -6342
rect 94874 -6662 94906 -6426
rect 95142 -6662 95226 -6426
rect 95462 -6662 95494 -6426
rect 94874 -7654 95494 -6662
rect 99994 -7066 100614 13000
rect 101394 10894 102014 13000
rect 101394 10658 101426 10894
rect 101662 10658 101746 10894
rect 101982 10658 102014 10894
rect 101394 10574 102014 10658
rect 101394 10338 101426 10574
rect 101662 10338 101746 10574
rect 101982 10338 102014 10574
rect 101394 -4186 102014 10338
rect 102794 -3226 103414 13000
rect 104194 3454 104814 13000
rect 104194 3218 104226 3454
rect 104462 3218 104546 3454
rect 104782 3218 104814 3454
rect 104194 3134 104814 3218
rect 104194 2898 104226 3134
rect 104462 2898 104546 3134
rect 104782 2898 104814 3134
rect 104194 -346 104814 2898
rect 104194 -582 104226 -346
rect 104462 -582 104546 -346
rect 104782 -582 104814 -346
rect 104194 -666 104814 -582
rect 104194 -902 104226 -666
rect 104462 -902 104546 -666
rect 104782 -902 104814 -666
rect 104194 -1894 104814 -902
rect 102794 -3462 102826 -3226
rect 103062 -3462 103146 -3226
rect 103382 -3462 103414 -3226
rect 102794 -3546 103414 -3462
rect 102794 -3782 102826 -3546
rect 103062 -3782 103146 -3546
rect 103382 -3782 103414 -3546
rect 102794 -3814 103414 -3782
rect 101394 -4422 101426 -4186
rect 101662 -4422 101746 -4186
rect 101982 -4422 102014 -4186
rect 101394 -4506 102014 -4422
rect 101394 -4742 101426 -4506
rect 101662 -4742 101746 -4506
rect 101982 -4742 102014 -4506
rect 101394 -5734 102014 -4742
rect 99994 -7302 100026 -7066
rect 100262 -7302 100346 -7066
rect 100582 -7302 100614 -7066
rect 99994 -7386 100614 -7302
rect 99994 -7622 100026 -7386
rect 100262 -7622 100346 -7386
rect 100582 -7622 100614 -7386
rect 99994 -7654 100614 -7622
rect 105114 -6106 105734 13000
rect 106514 -5146 107134 13000
rect 107914 7174 108534 13000
rect 107914 6938 107946 7174
rect 108182 6938 108266 7174
rect 108502 6938 108534 7174
rect 107914 6854 108534 6938
rect 107914 6618 107946 6854
rect 108182 6618 108266 6854
rect 108502 6618 108534 6854
rect 107914 -2266 108534 6618
rect 109314 -1306 109934 13000
rect 109314 -1542 109346 -1306
rect 109582 -1542 109666 -1306
rect 109902 -1542 109934 -1306
rect 109314 -1626 109934 -1542
rect 109314 -1862 109346 -1626
rect 109582 -1862 109666 -1626
rect 109902 -1862 109934 -1626
rect 109314 -1894 109934 -1862
rect 107914 -2502 107946 -2266
rect 108182 -2502 108266 -2266
rect 108502 -2502 108534 -2266
rect 107914 -2586 108534 -2502
rect 107914 -2822 107946 -2586
rect 108182 -2822 108266 -2586
rect 108502 -2822 108534 -2586
rect 107914 -3814 108534 -2822
rect 106514 -5382 106546 -5146
rect 106782 -5382 106866 -5146
rect 107102 -5382 107134 -5146
rect 106514 -5466 107134 -5382
rect 106514 -5702 106546 -5466
rect 106782 -5702 106866 -5466
rect 107102 -5702 107134 -5466
rect 106514 -5734 107134 -5702
rect 105114 -6342 105146 -6106
rect 105382 -6342 105466 -6106
rect 105702 -6342 105734 -6106
rect 105114 -6426 105734 -6342
rect 105114 -6662 105146 -6426
rect 105382 -6662 105466 -6426
rect 105702 -6662 105734 -6426
rect 105114 -7654 105734 -6662
rect 110234 -7066 110854 13000
rect 111634 10894 112254 13000
rect 111634 10658 111666 10894
rect 111902 10658 111986 10894
rect 112222 10658 112254 10894
rect 111634 10574 112254 10658
rect 111634 10338 111666 10574
rect 111902 10338 111986 10574
rect 112222 10338 112254 10574
rect 111634 -4186 112254 10338
rect 113034 -3226 113654 13000
rect 114434 3454 115054 13000
rect 114434 3218 114466 3454
rect 114702 3218 114786 3454
rect 115022 3218 115054 3454
rect 114434 3134 115054 3218
rect 114434 2898 114466 3134
rect 114702 2898 114786 3134
rect 115022 2898 115054 3134
rect 114434 -346 115054 2898
rect 114434 -582 114466 -346
rect 114702 -582 114786 -346
rect 115022 -582 115054 -346
rect 114434 -666 115054 -582
rect 114434 -902 114466 -666
rect 114702 -902 114786 -666
rect 115022 -902 115054 -666
rect 114434 -1894 115054 -902
rect 113034 -3462 113066 -3226
rect 113302 -3462 113386 -3226
rect 113622 -3462 113654 -3226
rect 113034 -3546 113654 -3462
rect 113034 -3782 113066 -3546
rect 113302 -3782 113386 -3546
rect 113622 -3782 113654 -3546
rect 113034 -3814 113654 -3782
rect 111634 -4422 111666 -4186
rect 111902 -4422 111986 -4186
rect 112222 -4422 112254 -4186
rect 111634 -4506 112254 -4422
rect 111634 -4742 111666 -4506
rect 111902 -4742 111986 -4506
rect 112222 -4742 112254 -4506
rect 111634 -5734 112254 -4742
rect 110234 -7302 110266 -7066
rect 110502 -7302 110586 -7066
rect 110822 -7302 110854 -7066
rect 110234 -7386 110854 -7302
rect 110234 -7622 110266 -7386
rect 110502 -7622 110586 -7386
rect 110822 -7622 110854 -7386
rect 110234 -7654 110854 -7622
rect 115354 -6106 115974 13000
rect 116754 -5146 117374 13000
rect 118154 7174 118774 13000
rect 118154 6938 118186 7174
rect 118422 6938 118506 7174
rect 118742 6938 118774 7174
rect 118154 6854 118774 6938
rect 118154 6618 118186 6854
rect 118422 6618 118506 6854
rect 118742 6618 118774 6854
rect 118154 -2266 118774 6618
rect 119554 -1306 120174 13000
rect 119554 -1542 119586 -1306
rect 119822 -1542 119906 -1306
rect 120142 -1542 120174 -1306
rect 119554 -1626 120174 -1542
rect 119554 -1862 119586 -1626
rect 119822 -1862 119906 -1626
rect 120142 -1862 120174 -1626
rect 119554 -1894 120174 -1862
rect 118154 -2502 118186 -2266
rect 118422 -2502 118506 -2266
rect 118742 -2502 118774 -2266
rect 118154 -2586 118774 -2502
rect 118154 -2822 118186 -2586
rect 118422 -2822 118506 -2586
rect 118742 -2822 118774 -2586
rect 118154 -3814 118774 -2822
rect 116754 -5382 116786 -5146
rect 117022 -5382 117106 -5146
rect 117342 -5382 117374 -5146
rect 116754 -5466 117374 -5382
rect 116754 -5702 116786 -5466
rect 117022 -5702 117106 -5466
rect 117342 -5702 117374 -5466
rect 116754 -5734 117374 -5702
rect 115354 -6342 115386 -6106
rect 115622 -6342 115706 -6106
rect 115942 -6342 115974 -6106
rect 115354 -6426 115974 -6342
rect 115354 -6662 115386 -6426
rect 115622 -6662 115706 -6426
rect 115942 -6662 115974 -6426
rect 115354 -7654 115974 -6662
rect 120474 -7066 121094 13000
rect 121874 10894 122494 13000
rect 121874 10658 121906 10894
rect 122142 10658 122226 10894
rect 122462 10658 122494 10894
rect 121874 10574 122494 10658
rect 121874 10338 121906 10574
rect 122142 10338 122226 10574
rect 122462 10338 122494 10574
rect 121874 -4186 122494 10338
rect 123274 -3226 123894 13000
rect 124674 3454 125294 13000
rect 124674 3218 124706 3454
rect 124942 3218 125026 3454
rect 125262 3218 125294 3454
rect 124674 3134 125294 3218
rect 124674 2898 124706 3134
rect 124942 2898 125026 3134
rect 125262 2898 125294 3134
rect 124674 -346 125294 2898
rect 124674 -582 124706 -346
rect 124942 -582 125026 -346
rect 125262 -582 125294 -346
rect 124674 -666 125294 -582
rect 124674 -902 124706 -666
rect 124942 -902 125026 -666
rect 125262 -902 125294 -666
rect 124674 -1894 125294 -902
rect 123274 -3462 123306 -3226
rect 123542 -3462 123626 -3226
rect 123862 -3462 123894 -3226
rect 123274 -3546 123894 -3462
rect 123274 -3782 123306 -3546
rect 123542 -3782 123626 -3546
rect 123862 -3782 123894 -3546
rect 123274 -3814 123894 -3782
rect 121874 -4422 121906 -4186
rect 122142 -4422 122226 -4186
rect 122462 -4422 122494 -4186
rect 121874 -4506 122494 -4422
rect 121874 -4742 121906 -4506
rect 122142 -4742 122226 -4506
rect 122462 -4742 122494 -4506
rect 121874 -5734 122494 -4742
rect 120474 -7302 120506 -7066
rect 120742 -7302 120826 -7066
rect 121062 -7302 121094 -7066
rect 120474 -7386 121094 -7302
rect 120474 -7622 120506 -7386
rect 120742 -7622 120826 -7386
rect 121062 -7622 121094 -7386
rect 120474 -7654 121094 -7622
rect 125594 -6106 126214 13000
rect 126994 -5146 127614 13000
rect 128394 7174 129014 13000
rect 128394 6938 128426 7174
rect 128662 6938 128746 7174
rect 128982 6938 129014 7174
rect 128394 6854 129014 6938
rect 128394 6618 128426 6854
rect 128662 6618 128746 6854
rect 128982 6618 129014 6854
rect 128394 -2266 129014 6618
rect 129794 -1306 130414 13000
rect 129794 -1542 129826 -1306
rect 130062 -1542 130146 -1306
rect 130382 -1542 130414 -1306
rect 129794 -1626 130414 -1542
rect 129794 -1862 129826 -1626
rect 130062 -1862 130146 -1626
rect 130382 -1862 130414 -1626
rect 129794 -1894 130414 -1862
rect 128394 -2502 128426 -2266
rect 128662 -2502 128746 -2266
rect 128982 -2502 129014 -2266
rect 128394 -2586 129014 -2502
rect 128394 -2822 128426 -2586
rect 128662 -2822 128746 -2586
rect 128982 -2822 129014 -2586
rect 128394 -3814 129014 -2822
rect 126994 -5382 127026 -5146
rect 127262 -5382 127346 -5146
rect 127582 -5382 127614 -5146
rect 126994 -5466 127614 -5382
rect 126994 -5702 127026 -5466
rect 127262 -5702 127346 -5466
rect 127582 -5702 127614 -5466
rect 126994 -5734 127614 -5702
rect 125594 -6342 125626 -6106
rect 125862 -6342 125946 -6106
rect 126182 -6342 126214 -6106
rect 125594 -6426 126214 -6342
rect 125594 -6662 125626 -6426
rect 125862 -6662 125946 -6426
rect 126182 -6662 126214 -6426
rect 125594 -7654 126214 -6662
rect 130714 -7066 131334 13000
rect 132114 10894 132734 13000
rect 132114 10658 132146 10894
rect 132382 10658 132466 10894
rect 132702 10658 132734 10894
rect 132114 10574 132734 10658
rect 132114 10338 132146 10574
rect 132382 10338 132466 10574
rect 132702 10338 132734 10574
rect 132114 -4186 132734 10338
rect 133514 -3226 134134 13000
rect 134914 3454 135534 13000
rect 134914 3218 134946 3454
rect 135182 3218 135266 3454
rect 135502 3218 135534 3454
rect 134914 3134 135534 3218
rect 134914 2898 134946 3134
rect 135182 2898 135266 3134
rect 135502 2898 135534 3134
rect 134914 -346 135534 2898
rect 134914 -582 134946 -346
rect 135182 -582 135266 -346
rect 135502 -582 135534 -346
rect 134914 -666 135534 -582
rect 134914 -902 134946 -666
rect 135182 -902 135266 -666
rect 135502 -902 135534 -666
rect 134914 -1894 135534 -902
rect 133514 -3462 133546 -3226
rect 133782 -3462 133866 -3226
rect 134102 -3462 134134 -3226
rect 133514 -3546 134134 -3462
rect 133514 -3782 133546 -3546
rect 133782 -3782 133866 -3546
rect 134102 -3782 134134 -3546
rect 133514 -3814 134134 -3782
rect 132114 -4422 132146 -4186
rect 132382 -4422 132466 -4186
rect 132702 -4422 132734 -4186
rect 132114 -4506 132734 -4422
rect 132114 -4742 132146 -4506
rect 132382 -4742 132466 -4506
rect 132702 -4742 132734 -4506
rect 132114 -5734 132734 -4742
rect 130714 -7302 130746 -7066
rect 130982 -7302 131066 -7066
rect 131302 -7302 131334 -7066
rect 130714 -7386 131334 -7302
rect 130714 -7622 130746 -7386
rect 130982 -7622 131066 -7386
rect 131302 -7622 131334 -7386
rect 130714 -7654 131334 -7622
rect 135834 -6106 136454 13000
rect 137234 -5146 137854 13000
rect 138634 7174 139254 13000
rect 138634 6938 138666 7174
rect 138902 6938 138986 7174
rect 139222 6938 139254 7174
rect 138634 6854 139254 6938
rect 138634 6618 138666 6854
rect 138902 6618 138986 6854
rect 139222 6618 139254 6854
rect 138634 -2266 139254 6618
rect 140034 -1306 140654 13000
rect 140034 -1542 140066 -1306
rect 140302 -1542 140386 -1306
rect 140622 -1542 140654 -1306
rect 140034 -1626 140654 -1542
rect 140034 -1862 140066 -1626
rect 140302 -1862 140386 -1626
rect 140622 -1862 140654 -1626
rect 140034 -1894 140654 -1862
rect 138634 -2502 138666 -2266
rect 138902 -2502 138986 -2266
rect 139222 -2502 139254 -2266
rect 138634 -2586 139254 -2502
rect 138634 -2822 138666 -2586
rect 138902 -2822 138986 -2586
rect 139222 -2822 139254 -2586
rect 138634 -3814 139254 -2822
rect 137234 -5382 137266 -5146
rect 137502 -5382 137586 -5146
rect 137822 -5382 137854 -5146
rect 137234 -5466 137854 -5382
rect 137234 -5702 137266 -5466
rect 137502 -5702 137586 -5466
rect 137822 -5702 137854 -5466
rect 137234 -5734 137854 -5702
rect 135834 -6342 135866 -6106
rect 136102 -6342 136186 -6106
rect 136422 -6342 136454 -6106
rect 135834 -6426 136454 -6342
rect 135834 -6662 135866 -6426
rect 136102 -6662 136186 -6426
rect 136422 -6662 136454 -6426
rect 135834 -7654 136454 -6662
rect 140954 -7066 141574 13000
rect 142354 10894 142974 13000
rect 142354 10658 142386 10894
rect 142622 10658 142706 10894
rect 142942 10658 142974 10894
rect 142354 10574 142974 10658
rect 142354 10338 142386 10574
rect 142622 10338 142706 10574
rect 142942 10338 142974 10574
rect 142354 -4186 142974 10338
rect 143754 -3226 144374 13000
rect 145154 3454 145774 13000
rect 145154 3218 145186 3454
rect 145422 3218 145506 3454
rect 145742 3218 145774 3454
rect 145154 3134 145774 3218
rect 145154 2898 145186 3134
rect 145422 2898 145506 3134
rect 145742 2898 145774 3134
rect 145154 -346 145774 2898
rect 145154 -582 145186 -346
rect 145422 -582 145506 -346
rect 145742 -582 145774 -346
rect 145154 -666 145774 -582
rect 145154 -902 145186 -666
rect 145422 -902 145506 -666
rect 145742 -902 145774 -666
rect 145154 -1894 145774 -902
rect 143754 -3462 143786 -3226
rect 144022 -3462 144106 -3226
rect 144342 -3462 144374 -3226
rect 143754 -3546 144374 -3462
rect 143754 -3782 143786 -3546
rect 144022 -3782 144106 -3546
rect 144342 -3782 144374 -3546
rect 143754 -3814 144374 -3782
rect 142354 -4422 142386 -4186
rect 142622 -4422 142706 -4186
rect 142942 -4422 142974 -4186
rect 142354 -4506 142974 -4422
rect 142354 -4742 142386 -4506
rect 142622 -4742 142706 -4506
rect 142942 -4742 142974 -4506
rect 142354 -5734 142974 -4742
rect 140954 -7302 140986 -7066
rect 141222 -7302 141306 -7066
rect 141542 -7302 141574 -7066
rect 140954 -7386 141574 -7302
rect 140954 -7622 140986 -7386
rect 141222 -7622 141306 -7386
rect 141542 -7622 141574 -7386
rect 140954 -7654 141574 -7622
rect 146074 -6106 146694 13000
rect 147474 -5146 148094 13000
rect 148874 7174 149494 13000
rect 148874 6938 148906 7174
rect 149142 6938 149226 7174
rect 149462 6938 149494 7174
rect 148874 6854 149494 6938
rect 148874 6618 148906 6854
rect 149142 6618 149226 6854
rect 149462 6618 149494 6854
rect 148874 -2266 149494 6618
rect 150274 -1306 150894 13000
rect 150274 -1542 150306 -1306
rect 150542 -1542 150626 -1306
rect 150862 -1542 150894 -1306
rect 150274 -1626 150894 -1542
rect 150274 -1862 150306 -1626
rect 150542 -1862 150626 -1626
rect 150862 -1862 150894 -1626
rect 150274 -1894 150894 -1862
rect 148874 -2502 148906 -2266
rect 149142 -2502 149226 -2266
rect 149462 -2502 149494 -2266
rect 148874 -2586 149494 -2502
rect 148874 -2822 148906 -2586
rect 149142 -2822 149226 -2586
rect 149462 -2822 149494 -2586
rect 148874 -3814 149494 -2822
rect 147474 -5382 147506 -5146
rect 147742 -5382 147826 -5146
rect 148062 -5382 148094 -5146
rect 147474 -5466 148094 -5382
rect 147474 -5702 147506 -5466
rect 147742 -5702 147826 -5466
rect 148062 -5702 148094 -5466
rect 147474 -5734 148094 -5702
rect 146074 -6342 146106 -6106
rect 146342 -6342 146426 -6106
rect 146662 -6342 146694 -6106
rect 146074 -6426 146694 -6342
rect 146074 -6662 146106 -6426
rect 146342 -6662 146426 -6426
rect 146662 -6662 146694 -6426
rect 146074 -7654 146694 -6662
rect 151194 -7066 151814 13000
rect 152594 10894 153214 13000
rect 152594 10658 152626 10894
rect 152862 10658 152946 10894
rect 153182 10658 153214 10894
rect 152594 10574 153214 10658
rect 152594 10338 152626 10574
rect 152862 10338 152946 10574
rect 153182 10338 153214 10574
rect 152594 -4186 153214 10338
rect 153994 -3226 154614 13000
rect 155394 3454 156014 13000
rect 155394 3218 155426 3454
rect 155662 3218 155746 3454
rect 155982 3218 156014 3454
rect 155394 3134 156014 3218
rect 155394 2898 155426 3134
rect 155662 2898 155746 3134
rect 155982 2898 156014 3134
rect 155394 -346 156014 2898
rect 155394 -582 155426 -346
rect 155662 -582 155746 -346
rect 155982 -582 156014 -346
rect 155394 -666 156014 -582
rect 155394 -902 155426 -666
rect 155662 -902 155746 -666
rect 155982 -902 156014 -666
rect 155394 -1894 156014 -902
rect 153994 -3462 154026 -3226
rect 154262 -3462 154346 -3226
rect 154582 -3462 154614 -3226
rect 153994 -3546 154614 -3462
rect 153994 -3782 154026 -3546
rect 154262 -3782 154346 -3546
rect 154582 -3782 154614 -3546
rect 153994 -3814 154614 -3782
rect 152594 -4422 152626 -4186
rect 152862 -4422 152946 -4186
rect 153182 -4422 153214 -4186
rect 152594 -4506 153214 -4422
rect 152594 -4742 152626 -4506
rect 152862 -4742 152946 -4506
rect 153182 -4742 153214 -4506
rect 152594 -5734 153214 -4742
rect 151194 -7302 151226 -7066
rect 151462 -7302 151546 -7066
rect 151782 -7302 151814 -7066
rect 151194 -7386 151814 -7302
rect 151194 -7622 151226 -7386
rect 151462 -7622 151546 -7386
rect 151782 -7622 151814 -7386
rect 151194 -7654 151814 -7622
rect 156314 -6106 156934 13000
rect 157714 -5146 158334 13000
rect 159114 7174 159734 13000
rect 159114 6938 159146 7174
rect 159382 6938 159466 7174
rect 159702 6938 159734 7174
rect 159114 6854 159734 6938
rect 159114 6618 159146 6854
rect 159382 6618 159466 6854
rect 159702 6618 159734 6854
rect 159114 -2266 159734 6618
rect 160514 -1306 161134 13000
rect 160514 -1542 160546 -1306
rect 160782 -1542 160866 -1306
rect 161102 -1542 161134 -1306
rect 160514 -1626 161134 -1542
rect 160514 -1862 160546 -1626
rect 160782 -1862 160866 -1626
rect 161102 -1862 161134 -1626
rect 160514 -1894 161134 -1862
rect 159114 -2502 159146 -2266
rect 159382 -2502 159466 -2266
rect 159702 -2502 159734 -2266
rect 159114 -2586 159734 -2502
rect 159114 -2822 159146 -2586
rect 159382 -2822 159466 -2586
rect 159702 -2822 159734 -2586
rect 159114 -3814 159734 -2822
rect 157714 -5382 157746 -5146
rect 157982 -5382 158066 -5146
rect 158302 -5382 158334 -5146
rect 157714 -5466 158334 -5382
rect 157714 -5702 157746 -5466
rect 157982 -5702 158066 -5466
rect 158302 -5702 158334 -5466
rect 157714 -5734 158334 -5702
rect 156314 -6342 156346 -6106
rect 156582 -6342 156666 -6106
rect 156902 -6342 156934 -6106
rect 156314 -6426 156934 -6342
rect 156314 -6662 156346 -6426
rect 156582 -6662 156666 -6426
rect 156902 -6662 156934 -6426
rect 156314 -7654 156934 -6662
rect 161434 -7066 162054 13000
rect 162834 10894 163454 13000
rect 162834 10658 162866 10894
rect 163102 10658 163186 10894
rect 163422 10658 163454 10894
rect 162834 10574 163454 10658
rect 162834 10338 162866 10574
rect 163102 10338 163186 10574
rect 163422 10338 163454 10574
rect 162834 -4186 163454 10338
rect 164234 -3226 164854 13000
rect 165634 3454 166254 13000
rect 165634 3218 165666 3454
rect 165902 3218 165986 3454
rect 166222 3218 166254 3454
rect 165634 3134 166254 3218
rect 165634 2898 165666 3134
rect 165902 2898 165986 3134
rect 166222 2898 166254 3134
rect 165634 -346 166254 2898
rect 165634 -582 165666 -346
rect 165902 -582 165986 -346
rect 166222 -582 166254 -346
rect 165634 -666 166254 -582
rect 165634 -902 165666 -666
rect 165902 -902 165986 -666
rect 166222 -902 166254 -666
rect 165634 -1894 166254 -902
rect 164234 -3462 164266 -3226
rect 164502 -3462 164586 -3226
rect 164822 -3462 164854 -3226
rect 164234 -3546 164854 -3462
rect 164234 -3782 164266 -3546
rect 164502 -3782 164586 -3546
rect 164822 -3782 164854 -3546
rect 164234 -3814 164854 -3782
rect 162834 -4422 162866 -4186
rect 163102 -4422 163186 -4186
rect 163422 -4422 163454 -4186
rect 162834 -4506 163454 -4422
rect 162834 -4742 162866 -4506
rect 163102 -4742 163186 -4506
rect 163422 -4742 163454 -4506
rect 162834 -5734 163454 -4742
rect 161434 -7302 161466 -7066
rect 161702 -7302 161786 -7066
rect 162022 -7302 162054 -7066
rect 161434 -7386 162054 -7302
rect 161434 -7622 161466 -7386
rect 161702 -7622 161786 -7386
rect 162022 -7622 162054 -7386
rect 161434 -7654 162054 -7622
rect 166554 -6106 167174 13000
rect 167954 -5146 168574 13000
rect 169354 7174 169974 13000
rect 169354 6938 169386 7174
rect 169622 6938 169706 7174
rect 169942 6938 169974 7174
rect 169354 6854 169974 6938
rect 169354 6618 169386 6854
rect 169622 6618 169706 6854
rect 169942 6618 169974 6854
rect 169354 -2266 169974 6618
rect 170754 -1306 171374 13000
rect 170754 -1542 170786 -1306
rect 171022 -1542 171106 -1306
rect 171342 -1542 171374 -1306
rect 170754 -1626 171374 -1542
rect 170754 -1862 170786 -1626
rect 171022 -1862 171106 -1626
rect 171342 -1862 171374 -1626
rect 170754 -1894 171374 -1862
rect 169354 -2502 169386 -2266
rect 169622 -2502 169706 -2266
rect 169942 -2502 169974 -2266
rect 169354 -2586 169974 -2502
rect 169354 -2822 169386 -2586
rect 169622 -2822 169706 -2586
rect 169942 -2822 169974 -2586
rect 169354 -3814 169974 -2822
rect 167954 -5382 167986 -5146
rect 168222 -5382 168306 -5146
rect 168542 -5382 168574 -5146
rect 167954 -5466 168574 -5382
rect 167954 -5702 167986 -5466
rect 168222 -5702 168306 -5466
rect 168542 -5702 168574 -5466
rect 167954 -5734 168574 -5702
rect 166554 -6342 166586 -6106
rect 166822 -6342 166906 -6106
rect 167142 -6342 167174 -6106
rect 166554 -6426 167174 -6342
rect 166554 -6662 166586 -6426
rect 166822 -6662 166906 -6426
rect 167142 -6662 167174 -6426
rect 166554 -7654 167174 -6662
rect 171674 -7066 172294 13000
rect 173074 10894 173694 13000
rect 173074 10658 173106 10894
rect 173342 10658 173426 10894
rect 173662 10658 173694 10894
rect 173074 10574 173694 10658
rect 173074 10338 173106 10574
rect 173342 10338 173426 10574
rect 173662 10338 173694 10574
rect 173074 -4186 173694 10338
rect 174474 -3226 175094 13000
rect 175874 3454 176494 13000
rect 175874 3218 175906 3454
rect 176142 3218 176226 3454
rect 176462 3218 176494 3454
rect 175874 3134 176494 3218
rect 175874 2898 175906 3134
rect 176142 2898 176226 3134
rect 176462 2898 176494 3134
rect 175874 -346 176494 2898
rect 175874 -582 175906 -346
rect 176142 -582 176226 -346
rect 176462 -582 176494 -346
rect 175874 -666 176494 -582
rect 175874 -902 175906 -666
rect 176142 -902 176226 -666
rect 176462 -902 176494 -666
rect 175874 -1894 176494 -902
rect 174474 -3462 174506 -3226
rect 174742 -3462 174826 -3226
rect 175062 -3462 175094 -3226
rect 174474 -3546 175094 -3462
rect 174474 -3782 174506 -3546
rect 174742 -3782 174826 -3546
rect 175062 -3782 175094 -3546
rect 174474 -3814 175094 -3782
rect 173074 -4422 173106 -4186
rect 173342 -4422 173426 -4186
rect 173662 -4422 173694 -4186
rect 173074 -4506 173694 -4422
rect 173074 -4742 173106 -4506
rect 173342 -4742 173426 -4506
rect 173662 -4742 173694 -4506
rect 173074 -5734 173694 -4742
rect 171674 -7302 171706 -7066
rect 171942 -7302 172026 -7066
rect 172262 -7302 172294 -7066
rect 171674 -7386 172294 -7302
rect 171674 -7622 171706 -7386
rect 171942 -7622 172026 -7386
rect 172262 -7622 172294 -7386
rect 171674 -7654 172294 -7622
rect 176794 -6106 177414 13000
rect 178194 -5146 178814 13000
rect 179594 7174 180214 13000
rect 179594 6938 179626 7174
rect 179862 6938 179946 7174
rect 180182 6938 180214 7174
rect 179594 6854 180214 6938
rect 179594 6618 179626 6854
rect 179862 6618 179946 6854
rect 180182 6618 180214 6854
rect 179594 -2266 180214 6618
rect 180994 -1306 181614 13000
rect 180994 -1542 181026 -1306
rect 181262 -1542 181346 -1306
rect 181582 -1542 181614 -1306
rect 180994 -1626 181614 -1542
rect 180994 -1862 181026 -1626
rect 181262 -1862 181346 -1626
rect 181582 -1862 181614 -1626
rect 180994 -1894 181614 -1862
rect 179594 -2502 179626 -2266
rect 179862 -2502 179946 -2266
rect 180182 -2502 180214 -2266
rect 179594 -2586 180214 -2502
rect 179594 -2822 179626 -2586
rect 179862 -2822 179946 -2586
rect 180182 -2822 180214 -2586
rect 179594 -3814 180214 -2822
rect 178194 -5382 178226 -5146
rect 178462 -5382 178546 -5146
rect 178782 -5382 178814 -5146
rect 178194 -5466 178814 -5382
rect 178194 -5702 178226 -5466
rect 178462 -5702 178546 -5466
rect 178782 -5702 178814 -5466
rect 178194 -5734 178814 -5702
rect 176794 -6342 176826 -6106
rect 177062 -6342 177146 -6106
rect 177382 -6342 177414 -6106
rect 176794 -6426 177414 -6342
rect 176794 -6662 176826 -6426
rect 177062 -6662 177146 -6426
rect 177382 -6662 177414 -6426
rect 176794 -7654 177414 -6662
rect 181914 -7066 182534 13000
rect 183314 10894 183934 13000
rect 183314 10658 183346 10894
rect 183582 10658 183666 10894
rect 183902 10658 183934 10894
rect 183314 10574 183934 10658
rect 183314 10338 183346 10574
rect 183582 10338 183666 10574
rect 183902 10338 183934 10574
rect 183314 -4186 183934 10338
rect 184714 -3226 185334 13000
rect 186114 3454 186734 13000
rect 186114 3218 186146 3454
rect 186382 3218 186466 3454
rect 186702 3218 186734 3454
rect 186114 3134 186734 3218
rect 186114 2898 186146 3134
rect 186382 2898 186466 3134
rect 186702 2898 186734 3134
rect 186114 -346 186734 2898
rect 186114 -582 186146 -346
rect 186382 -582 186466 -346
rect 186702 -582 186734 -346
rect 186114 -666 186734 -582
rect 186114 -902 186146 -666
rect 186382 -902 186466 -666
rect 186702 -902 186734 -666
rect 186114 -1894 186734 -902
rect 184714 -3462 184746 -3226
rect 184982 -3462 185066 -3226
rect 185302 -3462 185334 -3226
rect 184714 -3546 185334 -3462
rect 184714 -3782 184746 -3546
rect 184982 -3782 185066 -3546
rect 185302 -3782 185334 -3546
rect 184714 -3814 185334 -3782
rect 183314 -4422 183346 -4186
rect 183582 -4422 183666 -4186
rect 183902 -4422 183934 -4186
rect 183314 -4506 183934 -4422
rect 183314 -4742 183346 -4506
rect 183582 -4742 183666 -4506
rect 183902 -4742 183934 -4506
rect 183314 -5734 183934 -4742
rect 181914 -7302 181946 -7066
rect 182182 -7302 182266 -7066
rect 182502 -7302 182534 -7066
rect 181914 -7386 182534 -7302
rect 181914 -7622 181946 -7386
rect 182182 -7622 182266 -7386
rect 182502 -7622 182534 -7386
rect 181914 -7654 182534 -7622
rect 187034 -6106 187654 13000
rect 188434 -5146 189054 13000
rect 189834 7174 190454 13000
rect 189834 6938 189866 7174
rect 190102 6938 190186 7174
rect 190422 6938 190454 7174
rect 189834 6854 190454 6938
rect 189834 6618 189866 6854
rect 190102 6618 190186 6854
rect 190422 6618 190454 6854
rect 189834 -2266 190454 6618
rect 191234 -1306 191854 13000
rect 191234 -1542 191266 -1306
rect 191502 -1542 191586 -1306
rect 191822 -1542 191854 -1306
rect 191234 -1626 191854 -1542
rect 191234 -1862 191266 -1626
rect 191502 -1862 191586 -1626
rect 191822 -1862 191854 -1626
rect 191234 -1894 191854 -1862
rect 189834 -2502 189866 -2266
rect 190102 -2502 190186 -2266
rect 190422 -2502 190454 -2266
rect 189834 -2586 190454 -2502
rect 189834 -2822 189866 -2586
rect 190102 -2822 190186 -2586
rect 190422 -2822 190454 -2586
rect 189834 -3814 190454 -2822
rect 188434 -5382 188466 -5146
rect 188702 -5382 188786 -5146
rect 189022 -5382 189054 -5146
rect 188434 -5466 189054 -5382
rect 188434 -5702 188466 -5466
rect 188702 -5702 188786 -5466
rect 189022 -5702 189054 -5466
rect 188434 -5734 189054 -5702
rect 187034 -6342 187066 -6106
rect 187302 -6342 187386 -6106
rect 187622 -6342 187654 -6106
rect 187034 -6426 187654 -6342
rect 187034 -6662 187066 -6426
rect 187302 -6662 187386 -6426
rect 187622 -6662 187654 -6426
rect 187034 -7654 187654 -6662
rect 192154 -7066 192774 13000
rect 193554 10894 194174 13000
rect 193554 10658 193586 10894
rect 193822 10658 193906 10894
rect 194142 10658 194174 10894
rect 193554 10574 194174 10658
rect 193554 10338 193586 10574
rect 193822 10338 193906 10574
rect 194142 10338 194174 10574
rect 193554 -4186 194174 10338
rect 194954 -3226 195574 13000
rect 196354 3454 196974 13000
rect 196354 3218 196386 3454
rect 196622 3218 196706 3454
rect 196942 3218 196974 3454
rect 196354 3134 196974 3218
rect 196354 2898 196386 3134
rect 196622 2898 196706 3134
rect 196942 2898 196974 3134
rect 196354 -346 196974 2898
rect 196354 -582 196386 -346
rect 196622 -582 196706 -346
rect 196942 -582 196974 -346
rect 196354 -666 196974 -582
rect 196354 -902 196386 -666
rect 196622 -902 196706 -666
rect 196942 -902 196974 -666
rect 196354 -1894 196974 -902
rect 194954 -3462 194986 -3226
rect 195222 -3462 195306 -3226
rect 195542 -3462 195574 -3226
rect 194954 -3546 195574 -3462
rect 194954 -3782 194986 -3546
rect 195222 -3782 195306 -3546
rect 195542 -3782 195574 -3546
rect 194954 -3814 195574 -3782
rect 193554 -4422 193586 -4186
rect 193822 -4422 193906 -4186
rect 194142 -4422 194174 -4186
rect 193554 -4506 194174 -4422
rect 193554 -4742 193586 -4506
rect 193822 -4742 193906 -4506
rect 194142 -4742 194174 -4506
rect 193554 -5734 194174 -4742
rect 192154 -7302 192186 -7066
rect 192422 -7302 192506 -7066
rect 192742 -7302 192774 -7066
rect 192154 -7386 192774 -7302
rect 192154 -7622 192186 -7386
rect 192422 -7622 192506 -7386
rect 192742 -7622 192774 -7386
rect 192154 -7654 192774 -7622
rect 197274 -6106 197894 13000
rect 198674 -5146 199294 13000
rect 200074 7174 200694 13000
rect 200074 6938 200106 7174
rect 200342 6938 200426 7174
rect 200662 6938 200694 7174
rect 200074 6854 200694 6938
rect 200074 6618 200106 6854
rect 200342 6618 200426 6854
rect 200662 6618 200694 6854
rect 200074 -2266 200694 6618
rect 201474 -1306 202094 13000
rect 201474 -1542 201506 -1306
rect 201742 -1542 201826 -1306
rect 202062 -1542 202094 -1306
rect 201474 -1626 202094 -1542
rect 201474 -1862 201506 -1626
rect 201742 -1862 201826 -1626
rect 202062 -1862 202094 -1626
rect 201474 -1894 202094 -1862
rect 200074 -2502 200106 -2266
rect 200342 -2502 200426 -2266
rect 200662 -2502 200694 -2266
rect 200074 -2586 200694 -2502
rect 200074 -2822 200106 -2586
rect 200342 -2822 200426 -2586
rect 200662 -2822 200694 -2586
rect 200074 -3814 200694 -2822
rect 198674 -5382 198706 -5146
rect 198942 -5382 199026 -5146
rect 199262 -5382 199294 -5146
rect 198674 -5466 199294 -5382
rect 198674 -5702 198706 -5466
rect 198942 -5702 199026 -5466
rect 199262 -5702 199294 -5466
rect 198674 -5734 199294 -5702
rect 197274 -6342 197306 -6106
rect 197542 -6342 197626 -6106
rect 197862 -6342 197894 -6106
rect 197274 -6426 197894 -6342
rect 197274 -6662 197306 -6426
rect 197542 -6662 197626 -6426
rect 197862 -6662 197894 -6426
rect 197274 -7654 197894 -6662
rect 202394 -7066 203014 13000
rect 203794 10894 204414 13000
rect 203794 10658 203826 10894
rect 204062 10658 204146 10894
rect 204382 10658 204414 10894
rect 203794 10574 204414 10658
rect 203794 10338 203826 10574
rect 204062 10338 204146 10574
rect 204382 10338 204414 10574
rect 203794 -4186 204414 10338
rect 205194 -3226 205814 13000
rect 206594 3454 207214 13000
rect 206594 3218 206626 3454
rect 206862 3218 206946 3454
rect 207182 3218 207214 3454
rect 206594 3134 207214 3218
rect 206594 2898 206626 3134
rect 206862 2898 206946 3134
rect 207182 2898 207214 3134
rect 206594 -346 207214 2898
rect 206594 -582 206626 -346
rect 206862 -582 206946 -346
rect 207182 -582 207214 -346
rect 206594 -666 207214 -582
rect 206594 -902 206626 -666
rect 206862 -902 206946 -666
rect 207182 -902 207214 -666
rect 206594 -1894 207214 -902
rect 205194 -3462 205226 -3226
rect 205462 -3462 205546 -3226
rect 205782 -3462 205814 -3226
rect 205194 -3546 205814 -3462
rect 205194 -3782 205226 -3546
rect 205462 -3782 205546 -3546
rect 205782 -3782 205814 -3546
rect 205194 -3814 205814 -3782
rect 203794 -4422 203826 -4186
rect 204062 -4422 204146 -4186
rect 204382 -4422 204414 -4186
rect 203794 -4506 204414 -4422
rect 203794 -4742 203826 -4506
rect 204062 -4742 204146 -4506
rect 204382 -4742 204414 -4506
rect 203794 -5734 204414 -4742
rect 202394 -7302 202426 -7066
rect 202662 -7302 202746 -7066
rect 202982 -7302 203014 -7066
rect 202394 -7386 203014 -7302
rect 202394 -7622 202426 -7386
rect 202662 -7622 202746 -7386
rect 202982 -7622 203014 -7386
rect 202394 -7654 203014 -7622
rect 207514 -6106 208134 13000
rect 208914 -5146 209534 13000
rect 210314 7174 210934 13000
rect 210314 6938 210346 7174
rect 210582 6938 210666 7174
rect 210902 6938 210934 7174
rect 210314 6854 210934 6938
rect 210314 6618 210346 6854
rect 210582 6618 210666 6854
rect 210902 6618 210934 6854
rect 210314 -2266 210934 6618
rect 211714 -1306 212334 13000
rect 211714 -1542 211746 -1306
rect 211982 -1542 212066 -1306
rect 212302 -1542 212334 -1306
rect 211714 -1626 212334 -1542
rect 211714 -1862 211746 -1626
rect 211982 -1862 212066 -1626
rect 212302 -1862 212334 -1626
rect 211714 -1894 212334 -1862
rect 210314 -2502 210346 -2266
rect 210582 -2502 210666 -2266
rect 210902 -2502 210934 -2266
rect 210314 -2586 210934 -2502
rect 210314 -2822 210346 -2586
rect 210582 -2822 210666 -2586
rect 210902 -2822 210934 -2586
rect 210314 -3814 210934 -2822
rect 208914 -5382 208946 -5146
rect 209182 -5382 209266 -5146
rect 209502 -5382 209534 -5146
rect 208914 -5466 209534 -5382
rect 208914 -5702 208946 -5466
rect 209182 -5702 209266 -5466
rect 209502 -5702 209534 -5466
rect 208914 -5734 209534 -5702
rect 207514 -6342 207546 -6106
rect 207782 -6342 207866 -6106
rect 208102 -6342 208134 -6106
rect 207514 -6426 208134 -6342
rect 207514 -6662 207546 -6426
rect 207782 -6662 207866 -6426
rect 208102 -6662 208134 -6426
rect 207514 -7654 208134 -6662
rect 212634 -7066 213254 13000
rect 214034 10894 214654 13000
rect 214034 10658 214066 10894
rect 214302 10658 214386 10894
rect 214622 10658 214654 10894
rect 214034 10574 214654 10658
rect 214034 10338 214066 10574
rect 214302 10338 214386 10574
rect 214622 10338 214654 10574
rect 214034 -4186 214654 10338
rect 215434 -3226 216054 13000
rect 216834 3454 217454 13000
rect 216834 3218 216866 3454
rect 217102 3218 217186 3454
rect 217422 3218 217454 3454
rect 216834 3134 217454 3218
rect 216834 2898 216866 3134
rect 217102 2898 217186 3134
rect 217422 2898 217454 3134
rect 216834 -346 217454 2898
rect 216834 -582 216866 -346
rect 217102 -582 217186 -346
rect 217422 -582 217454 -346
rect 216834 -666 217454 -582
rect 216834 -902 216866 -666
rect 217102 -902 217186 -666
rect 217422 -902 217454 -666
rect 216834 -1894 217454 -902
rect 215434 -3462 215466 -3226
rect 215702 -3462 215786 -3226
rect 216022 -3462 216054 -3226
rect 215434 -3546 216054 -3462
rect 215434 -3782 215466 -3546
rect 215702 -3782 215786 -3546
rect 216022 -3782 216054 -3546
rect 215434 -3814 216054 -3782
rect 214034 -4422 214066 -4186
rect 214302 -4422 214386 -4186
rect 214622 -4422 214654 -4186
rect 214034 -4506 214654 -4422
rect 214034 -4742 214066 -4506
rect 214302 -4742 214386 -4506
rect 214622 -4742 214654 -4506
rect 214034 -5734 214654 -4742
rect 212634 -7302 212666 -7066
rect 212902 -7302 212986 -7066
rect 213222 -7302 213254 -7066
rect 212634 -7386 213254 -7302
rect 212634 -7622 212666 -7386
rect 212902 -7622 212986 -7386
rect 213222 -7622 213254 -7386
rect 212634 -7654 213254 -7622
rect 217754 -6106 218374 13000
rect 219154 -5146 219774 13000
rect 220554 7174 221174 13000
rect 220554 6938 220586 7174
rect 220822 6938 220906 7174
rect 221142 6938 221174 7174
rect 220554 6854 221174 6938
rect 220554 6618 220586 6854
rect 220822 6618 220906 6854
rect 221142 6618 221174 6854
rect 220554 -2266 221174 6618
rect 221954 -1306 222574 13000
rect 221954 -1542 221986 -1306
rect 222222 -1542 222306 -1306
rect 222542 -1542 222574 -1306
rect 221954 -1626 222574 -1542
rect 221954 -1862 221986 -1626
rect 222222 -1862 222306 -1626
rect 222542 -1862 222574 -1626
rect 221954 -1894 222574 -1862
rect 220554 -2502 220586 -2266
rect 220822 -2502 220906 -2266
rect 221142 -2502 221174 -2266
rect 220554 -2586 221174 -2502
rect 220554 -2822 220586 -2586
rect 220822 -2822 220906 -2586
rect 221142 -2822 221174 -2586
rect 220554 -3814 221174 -2822
rect 219154 -5382 219186 -5146
rect 219422 -5382 219506 -5146
rect 219742 -5382 219774 -5146
rect 219154 -5466 219774 -5382
rect 219154 -5702 219186 -5466
rect 219422 -5702 219506 -5466
rect 219742 -5702 219774 -5466
rect 219154 -5734 219774 -5702
rect 217754 -6342 217786 -6106
rect 218022 -6342 218106 -6106
rect 218342 -6342 218374 -6106
rect 217754 -6426 218374 -6342
rect 217754 -6662 217786 -6426
rect 218022 -6662 218106 -6426
rect 218342 -6662 218374 -6426
rect 217754 -7654 218374 -6662
rect 222874 -7066 223494 13000
rect 224274 10894 224894 13000
rect 224274 10658 224306 10894
rect 224542 10658 224626 10894
rect 224862 10658 224894 10894
rect 224274 10574 224894 10658
rect 224274 10338 224306 10574
rect 224542 10338 224626 10574
rect 224862 10338 224894 10574
rect 224274 -4186 224894 10338
rect 225674 -3226 226294 13000
rect 227074 3454 227694 13000
rect 227074 3218 227106 3454
rect 227342 3218 227426 3454
rect 227662 3218 227694 3454
rect 227074 3134 227694 3218
rect 227074 2898 227106 3134
rect 227342 2898 227426 3134
rect 227662 2898 227694 3134
rect 227074 -346 227694 2898
rect 227074 -582 227106 -346
rect 227342 -582 227426 -346
rect 227662 -582 227694 -346
rect 227074 -666 227694 -582
rect 227074 -902 227106 -666
rect 227342 -902 227426 -666
rect 227662 -902 227694 -666
rect 227074 -1894 227694 -902
rect 225674 -3462 225706 -3226
rect 225942 -3462 226026 -3226
rect 226262 -3462 226294 -3226
rect 225674 -3546 226294 -3462
rect 225674 -3782 225706 -3546
rect 225942 -3782 226026 -3546
rect 226262 -3782 226294 -3546
rect 225674 -3814 226294 -3782
rect 224274 -4422 224306 -4186
rect 224542 -4422 224626 -4186
rect 224862 -4422 224894 -4186
rect 224274 -4506 224894 -4422
rect 224274 -4742 224306 -4506
rect 224542 -4742 224626 -4506
rect 224862 -4742 224894 -4506
rect 224274 -5734 224894 -4742
rect 222874 -7302 222906 -7066
rect 223142 -7302 223226 -7066
rect 223462 -7302 223494 -7066
rect 222874 -7386 223494 -7302
rect 222874 -7622 222906 -7386
rect 223142 -7622 223226 -7386
rect 223462 -7622 223494 -7386
rect 222874 -7654 223494 -7622
rect 227994 -6106 228614 13000
rect 229394 -5146 230014 13000
rect 230794 7174 231414 13000
rect 230794 6938 230826 7174
rect 231062 6938 231146 7174
rect 231382 6938 231414 7174
rect 230794 6854 231414 6938
rect 230794 6618 230826 6854
rect 231062 6618 231146 6854
rect 231382 6618 231414 6854
rect 230794 -2266 231414 6618
rect 232194 -1306 232814 13000
rect 232194 -1542 232226 -1306
rect 232462 -1542 232546 -1306
rect 232782 -1542 232814 -1306
rect 232194 -1626 232814 -1542
rect 232194 -1862 232226 -1626
rect 232462 -1862 232546 -1626
rect 232782 -1862 232814 -1626
rect 232194 -1894 232814 -1862
rect 230794 -2502 230826 -2266
rect 231062 -2502 231146 -2266
rect 231382 -2502 231414 -2266
rect 230794 -2586 231414 -2502
rect 230794 -2822 230826 -2586
rect 231062 -2822 231146 -2586
rect 231382 -2822 231414 -2586
rect 230794 -3814 231414 -2822
rect 229394 -5382 229426 -5146
rect 229662 -5382 229746 -5146
rect 229982 -5382 230014 -5146
rect 229394 -5466 230014 -5382
rect 229394 -5702 229426 -5466
rect 229662 -5702 229746 -5466
rect 229982 -5702 230014 -5466
rect 229394 -5734 230014 -5702
rect 227994 -6342 228026 -6106
rect 228262 -6342 228346 -6106
rect 228582 -6342 228614 -6106
rect 227994 -6426 228614 -6342
rect 227994 -6662 228026 -6426
rect 228262 -6662 228346 -6426
rect 228582 -6662 228614 -6426
rect 227994 -7654 228614 -6662
rect 233114 -7066 233734 13000
rect 234514 10894 235134 13000
rect 234514 10658 234546 10894
rect 234782 10658 234866 10894
rect 235102 10658 235134 10894
rect 234514 10574 235134 10658
rect 234514 10338 234546 10574
rect 234782 10338 234866 10574
rect 235102 10338 235134 10574
rect 234514 -4186 235134 10338
rect 235914 -3226 236534 13000
rect 237314 3454 237934 13000
rect 237314 3218 237346 3454
rect 237582 3218 237666 3454
rect 237902 3218 237934 3454
rect 237314 3134 237934 3218
rect 237314 2898 237346 3134
rect 237582 2898 237666 3134
rect 237902 2898 237934 3134
rect 237314 -346 237934 2898
rect 237314 -582 237346 -346
rect 237582 -582 237666 -346
rect 237902 -582 237934 -346
rect 237314 -666 237934 -582
rect 237314 -902 237346 -666
rect 237582 -902 237666 -666
rect 237902 -902 237934 -666
rect 237314 -1894 237934 -902
rect 235914 -3462 235946 -3226
rect 236182 -3462 236266 -3226
rect 236502 -3462 236534 -3226
rect 235914 -3546 236534 -3462
rect 235914 -3782 235946 -3546
rect 236182 -3782 236266 -3546
rect 236502 -3782 236534 -3546
rect 235914 -3814 236534 -3782
rect 234514 -4422 234546 -4186
rect 234782 -4422 234866 -4186
rect 235102 -4422 235134 -4186
rect 234514 -4506 235134 -4422
rect 234514 -4742 234546 -4506
rect 234782 -4742 234866 -4506
rect 235102 -4742 235134 -4506
rect 234514 -5734 235134 -4742
rect 233114 -7302 233146 -7066
rect 233382 -7302 233466 -7066
rect 233702 -7302 233734 -7066
rect 233114 -7386 233734 -7302
rect 233114 -7622 233146 -7386
rect 233382 -7622 233466 -7386
rect 233702 -7622 233734 -7386
rect 233114 -7654 233734 -7622
rect 238234 -6106 238854 13000
rect 239634 -5146 240254 13000
rect 241034 7174 241654 13000
rect 241034 6938 241066 7174
rect 241302 6938 241386 7174
rect 241622 6938 241654 7174
rect 241034 6854 241654 6938
rect 241034 6618 241066 6854
rect 241302 6618 241386 6854
rect 241622 6618 241654 6854
rect 241034 -2266 241654 6618
rect 242434 -1306 243054 13000
rect 242434 -1542 242466 -1306
rect 242702 -1542 242786 -1306
rect 243022 -1542 243054 -1306
rect 242434 -1626 243054 -1542
rect 242434 -1862 242466 -1626
rect 242702 -1862 242786 -1626
rect 243022 -1862 243054 -1626
rect 242434 -1894 243054 -1862
rect 241034 -2502 241066 -2266
rect 241302 -2502 241386 -2266
rect 241622 -2502 241654 -2266
rect 241034 -2586 241654 -2502
rect 241034 -2822 241066 -2586
rect 241302 -2822 241386 -2586
rect 241622 -2822 241654 -2586
rect 241034 -3814 241654 -2822
rect 239634 -5382 239666 -5146
rect 239902 -5382 239986 -5146
rect 240222 -5382 240254 -5146
rect 239634 -5466 240254 -5382
rect 239634 -5702 239666 -5466
rect 239902 -5702 239986 -5466
rect 240222 -5702 240254 -5466
rect 239634 -5734 240254 -5702
rect 238234 -6342 238266 -6106
rect 238502 -6342 238586 -6106
rect 238822 -6342 238854 -6106
rect 238234 -6426 238854 -6342
rect 238234 -6662 238266 -6426
rect 238502 -6662 238586 -6426
rect 238822 -6662 238854 -6426
rect 238234 -7654 238854 -6662
rect 243354 -7066 243974 13000
rect 244754 10894 245374 13000
rect 244754 10658 244786 10894
rect 245022 10658 245106 10894
rect 245342 10658 245374 10894
rect 244754 10574 245374 10658
rect 244754 10338 244786 10574
rect 245022 10338 245106 10574
rect 245342 10338 245374 10574
rect 244754 -4186 245374 10338
rect 246154 -3226 246774 13000
rect 247554 3454 248174 13000
rect 247554 3218 247586 3454
rect 247822 3218 247906 3454
rect 248142 3218 248174 3454
rect 247554 3134 248174 3218
rect 247554 2898 247586 3134
rect 247822 2898 247906 3134
rect 248142 2898 248174 3134
rect 247554 -346 248174 2898
rect 247554 -582 247586 -346
rect 247822 -582 247906 -346
rect 248142 -582 248174 -346
rect 247554 -666 248174 -582
rect 247554 -902 247586 -666
rect 247822 -902 247906 -666
rect 248142 -902 248174 -666
rect 247554 -1894 248174 -902
rect 246154 -3462 246186 -3226
rect 246422 -3462 246506 -3226
rect 246742 -3462 246774 -3226
rect 246154 -3546 246774 -3462
rect 246154 -3782 246186 -3546
rect 246422 -3782 246506 -3546
rect 246742 -3782 246774 -3546
rect 246154 -3814 246774 -3782
rect 244754 -4422 244786 -4186
rect 245022 -4422 245106 -4186
rect 245342 -4422 245374 -4186
rect 244754 -4506 245374 -4422
rect 244754 -4742 244786 -4506
rect 245022 -4742 245106 -4506
rect 245342 -4742 245374 -4506
rect 244754 -5734 245374 -4742
rect 243354 -7302 243386 -7066
rect 243622 -7302 243706 -7066
rect 243942 -7302 243974 -7066
rect 243354 -7386 243974 -7302
rect 243354 -7622 243386 -7386
rect 243622 -7622 243706 -7386
rect 243942 -7622 243974 -7386
rect 243354 -7654 243974 -7622
rect 248474 -6106 249094 13000
rect 249874 -5146 250494 13000
rect 251274 7174 251894 13000
rect 251274 6938 251306 7174
rect 251542 6938 251626 7174
rect 251862 6938 251894 7174
rect 251274 6854 251894 6938
rect 251274 6618 251306 6854
rect 251542 6618 251626 6854
rect 251862 6618 251894 6854
rect 251274 -2266 251894 6618
rect 252674 -1306 253294 13000
rect 252674 -1542 252706 -1306
rect 252942 -1542 253026 -1306
rect 253262 -1542 253294 -1306
rect 252674 -1626 253294 -1542
rect 252674 -1862 252706 -1626
rect 252942 -1862 253026 -1626
rect 253262 -1862 253294 -1626
rect 252674 -1894 253294 -1862
rect 251274 -2502 251306 -2266
rect 251542 -2502 251626 -2266
rect 251862 -2502 251894 -2266
rect 251274 -2586 251894 -2502
rect 251274 -2822 251306 -2586
rect 251542 -2822 251626 -2586
rect 251862 -2822 251894 -2586
rect 251274 -3814 251894 -2822
rect 249874 -5382 249906 -5146
rect 250142 -5382 250226 -5146
rect 250462 -5382 250494 -5146
rect 249874 -5466 250494 -5382
rect 249874 -5702 249906 -5466
rect 250142 -5702 250226 -5466
rect 250462 -5702 250494 -5466
rect 249874 -5734 250494 -5702
rect 248474 -6342 248506 -6106
rect 248742 -6342 248826 -6106
rect 249062 -6342 249094 -6106
rect 248474 -6426 249094 -6342
rect 248474 -6662 248506 -6426
rect 248742 -6662 248826 -6426
rect 249062 -6662 249094 -6426
rect 248474 -7654 249094 -6662
rect 253594 -7066 254214 13000
rect 254994 10894 255614 13000
rect 254994 10658 255026 10894
rect 255262 10658 255346 10894
rect 255582 10658 255614 10894
rect 254994 10574 255614 10658
rect 254994 10338 255026 10574
rect 255262 10338 255346 10574
rect 255582 10338 255614 10574
rect 254994 -4186 255614 10338
rect 256394 -3226 257014 13000
rect 257794 3454 258414 13000
rect 257794 3218 257826 3454
rect 258062 3218 258146 3454
rect 258382 3218 258414 3454
rect 257794 3134 258414 3218
rect 257794 2898 257826 3134
rect 258062 2898 258146 3134
rect 258382 2898 258414 3134
rect 257794 -346 258414 2898
rect 257794 -582 257826 -346
rect 258062 -582 258146 -346
rect 258382 -582 258414 -346
rect 257794 -666 258414 -582
rect 257794 -902 257826 -666
rect 258062 -902 258146 -666
rect 258382 -902 258414 -666
rect 257794 -1894 258414 -902
rect 256394 -3462 256426 -3226
rect 256662 -3462 256746 -3226
rect 256982 -3462 257014 -3226
rect 256394 -3546 257014 -3462
rect 256394 -3782 256426 -3546
rect 256662 -3782 256746 -3546
rect 256982 -3782 257014 -3546
rect 256394 -3814 257014 -3782
rect 254994 -4422 255026 -4186
rect 255262 -4422 255346 -4186
rect 255582 -4422 255614 -4186
rect 254994 -4506 255614 -4422
rect 254994 -4742 255026 -4506
rect 255262 -4742 255346 -4506
rect 255582 -4742 255614 -4506
rect 254994 -5734 255614 -4742
rect 253594 -7302 253626 -7066
rect 253862 -7302 253946 -7066
rect 254182 -7302 254214 -7066
rect 253594 -7386 254214 -7302
rect 253594 -7622 253626 -7386
rect 253862 -7622 253946 -7386
rect 254182 -7622 254214 -7386
rect 253594 -7654 254214 -7622
rect 258714 -6106 259334 13000
rect 260114 -5146 260734 13000
rect 261514 7174 262134 13000
rect 261514 6938 261546 7174
rect 261782 6938 261866 7174
rect 262102 6938 262134 7174
rect 261514 6854 262134 6938
rect 261514 6618 261546 6854
rect 261782 6618 261866 6854
rect 262102 6618 262134 6854
rect 261514 -2266 262134 6618
rect 262914 -1306 263534 13000
rect 262914 -1542 262946 -1306
rect 263182 -1542 263266 -1306
rect 263502 -1542 263534 -1306
rect 262914 -1626 263534 -1542
rect 262914 -1862 262946 -1626
rect 263182 -1862 263266 -1626
rect 263502 -1862 263534 -1626
rect 262914 -1894 263534 -1862
rect 261514 -2502 261546 -2266
rect 261782 -2502 261866 -2266
rect 262102 -2502 262134 -2266
rect 261514 -2586 262134 -2502
rect 261514 -2822 261546 -2586
rect 261782 -2822 261866 -2586
rect 262102 -2822 262134 -2586
rect 261514 -3814 262134 -2822
rect 260114 -5382 260146 -5146
rect 260382 -5382 260466 -5146
rect 260702 -5382 260734 -5146
rect 260114 -5466 260734 -5382
rect 260114 -5702 260146 -5466
rect 260382 -5702 260466 -5466
rect 260702 -5702 260734 -5466
rect 260114 -5734 260734 -5702
rect 258714 -6342 258746 -6106
rect 258982 -6342 259066 -6106
rect 259302 -6342 259334 -6106
rect 258714 -6426 259334 -6342
rect 258714 -6662 258746 -6426
rect 258982 -6662 259066 -6426
rect 259302 -6662 259334 -6426
rect 258714 -7654 259334 -6662
rect 263834 -7066 264454 13000
rect 265234 10894 265854 13000
rect 265234 10658 265266 10894
rect 265502 10658 265586 10894
rect 265822 10658 265854 10894
rect 265234 10574 265854 10658
rect 265234 10338 265266 10574
rect 265502 10338 265586 10574
rect 265822 10338 265854 10574
rect 265234 -4186 265854 10338
rect 266634 -3226 267254 13000
rect 268034 3454 268654 13000
rect 268034 3218 268066 3454
rect 268302 3218 268386 3454
rect 268622 3218 268654 3454
rect 268034 3134 268654 3218
rect 268034 2898 268066 3134
rect 268302 2898 268386 3134
rect 268622 2898 268654 3134
rect 268034 -346 268654 2898
rect 268034 -582 268066 -346
rect 268302 -582 268386 -346
rect 268622 -582 268654 -346
rect 268034 -666 268654 -582
rect 268034 -902 268066 -666
rect 268302 -902 268386 -666
rect 268622 -902 268654 -666
rect 268034 -1894 268654 -902
rect 266634 -3462 266666 -3226
rect 266902 -3462 266986 -3226
rect 267222 -3462 267254 -3226
rect 266634 -3546 267254 -3462
rect 266634 -3782 266666 -3546
rect 266902 -3782 266986 -3546
rect 267222 -3782 267254 -3546
rect 266634 -3814 267254 -3782
rect 265234 -4422 265266 -4186
rect 265502 -4422 265586 -4186
rect 265822 -4422 265854 -4186
rect 265234 -4506 265854 -4422
rect 265234 -4742 265266 -4506
rect 265502 -4742 265586 -4506
rect 265822 -4742 265854 -4506
rect 265234 -5734 265854 -4742
rect 263834 -7302 263866 -7066
rect 264102 -7302 264186 -7066
rect 264422 -7302 264454 -7066
rect 263834 -7386 264454 -7302
rect 263834 -7622 263866 -7386
rect 264102 -7622 264186 -7386
rect 264422 -7622 264454 -7386
rect 263834 -7654 264454 -7622
rect 268954 -6106 269574 13000
rect 270354 -5146 270974 13000
rect 271754 7174 272374 13000
rect 271754 6938 271786 7174
rect 272022 6938 272106 7174
rect 272342 6938 272374 7174
rect 271754 6854 272374 6938
rect 271754 6618 271786 6854
rect 272022 6618 272106 6854
rect 272342 6618 272374 6854
rect 271754 -2266 272374 6618
rect 273154 -1306 273774 13000
rect 273154 -1542 273186 -1306
rect 273422 -1542 273506 -1306
rect 273742 -1542 273774 -1306
rect 273154 -1626 273774 -1542
rect 273154 -1862 273186 -1626
rect 273422 -1862 273506 -1626
rect 273742 -1862 273774 -1626
rect 273154 -1894 273774 -1862
rect 271754 -2502 271786 -2266
rect 272022 -2502 272106 -2266
rect 272342 -2502 272374 -2266
rect 271754 -2586 272374 -2502
rect 271754 -2822 271786 -2586
rect 272022 -2822 272106 -2586
rect 272342 -2822 272374 -2586
rect 271754 -3814 272374 -2822
rect 270354 -5382 270386 -5146
rect 270622 -5382 270706 -5146
rect 270942 -5382 270974 -5146
rect 270354 -5466 270974 -5382
rect 270354 -5702 270386 -5466
rect 270622 -5702 270706 -5466
rect 270942 -5702 270974 -5466
rect 270354 -5734 270974 -5702
rect 268954 -6342 268986 -6106
rect 269222 -6342 269306 -6106
rect 269542 -6342 269574 -6106
rect 268954 -6426 269574 -6342
rect 268954 -6662 268986 -6426
rect 269222 -6662 269306 -6426
rect 269542 -6662 269574 -6426
rect 268954 -7654 269574 -6662
rect 274074 -7066 274694 13000
rect 275474 10894 276094 13000
rect 275474 10658 275506 10894
rect 275742 10658 275826 10894
rect 276062 10658 276094 10894
rect 275474 10574 276094 10658
rect 275474 10338 275506 10574
rect 275742 10338 275826 10574
rect 276062 10338 276094 10574
rect 275474 -4186 276094 10338
rect 276874 -3226 277494 13000
rect 278274 3454 278894 13000
rect 278274 3218 278306 3454
rect 278542 3218 278626 3454
rect 278862 3218 278894 3454
rect 278274 3134 278894 3218
rect 278274 2898 278306 3134
rect 278542 2898 278626 3134
rect 278862 2898 278894 3134
rect 278274 -346 278894 2898
rect 278274 -582 278306 -346
rect 278542 -582 278626 -346
rect 278862 -582 278894 -346
rect 278274 -666 278894 -582
rect 278274 -902 278306 -666
rect 278542 -902 278626 -666
rect 278862 -902 278894 -666
rect 278274 -1894 278894 -902
rect 276874 -3462 276906 -3226
rect 277142 -3462 277226 -3226
rect 277462 -3462 277494 -3226
rect 276874 -3546 277494 -3462
rect 276874 -3782 276906 -3546
rect 277142 -3782 277226 -3546
rect 277462 -3782 277494 -3546
rect 276874 -3814 277494 -3782
rect 275474 -4422 275506 -4186
rect 275742 -4422 275826 -4186
rect 276062 -4422 276094 -4186
rect 275474 -4506 276094 -4422
rect 275474 -4742 275506 -4506
rect 275742 -4742 275826 -4506
rect 276062 -4742 276094 -4506
rect 275474 -5734 276094 -4742
rect 274074 -7302 274106 -7066
rect 274342 -7302 274426 -7066
rect 274662 -7302 274694 -7066
rect 274074 -7386 274694 -7302
rect 274074 -7622 274106 -7386
rect 274342 -7622 274426 -7386
rect 274662 -7622 274694 -7386
rect 274074 -7654 274694 -7622
rect 279194 -6106 279814 13000
rect 280594 -5146 281214 13000
rect 281994 7174 282614 13000
rect 281994 6938 282026 7174
rect 282262 6938 282346 7174
rect 282582 6938 282614 7174
rect 281994 6854 282614 6938
rect 281994 6618 282026 6854
rect 282262 6618 282346 6854
rect 282582 6618 282614 6854
rect 281994 -2266 282614 6618
rect 283394 -1306 284014 13000
rect 283394 -1542 283426 -1306
rect 283662 -1542 283746 -1306
rect 283982 -1542 284014 -1306
rect 283394 -1626 284014 -1542
rect 283394 -1862 283426 -1626
rect 283662 -1862 283746 -1626
rect 283982 -1862 284014 -1626
rect 283394 -1894 284014 -1862
rect 281994 -2502 282026 -2266
rect 282262 -2502 282346 -2266
rect 282582 -2502 282614 -2266
rect 281994 -2586 282614 -2502
rect 281994 -2822 282026 -2586
rect 282262 -2822 282346 -2586
rect 282582 -2822 282614 -2586
rect 281994 -3814 282614 -2822
rect 280594 -5382 280626 -5146
rect 280862 -5382 280946 -5146
rect 281182 -5382 281214 -5146
rect 280594 -5466 281214 -5382
rect 280594 -5702 280626 -5466
rect 280862 -5702 280946 -5466
rect 281182 -5702 281214 -5466
rect 280594 -5734 281214 -5702
rect 279194 -6342 279226 -6106
rect 279462 -6342 279546 -6106
rect 279782 -6342 279814 -6106
rect 279194 -6426 279814 -6342
rect 279194 -6662 279226 -6426
rect 279462 -6662 279546 -6426
rect 279782 -6662 279814 -6426
rect 279194 -7654 279814 -6662
rect 284314 -7066 284934 13000
rect 285714 10894 286334 13000
rect 285714 10658 285746 10894
rect 285982 10658 286066 10894
rect 286302 10658 286334 10894
rect 285714 10574 286334 10658
rect 285714 10338 285746 10574
rect 285982 10338 286066 10574
rect 286302 10338 286334 10574
rect 285714 -4186 286334 10338
rect 287114 -3226 287734 13000
rect 288514 3454 289134 13000
rect 288514 3218 288546 3454
rect 288782 3218 288866 3454
rect 289102 3218 289134 3454
rect 288514 3134 289134 3218
rect 288514 2898 288546 3134
rect 288782 2898 288866 3134
rect 289102 2898 289134 3134
rect 288514 -346 289134 2898
rect 288514 -582 288546 -346
rect 288782 -582 288866 -346
rect 289102 -582 289134 -346
rect 288514 -666 289134 -582
rect 288514 -902 288546 -666
rect 288782 -902 288866 -666
rect 289102 -902 289134 -666
rect 288514 -1894 289134 -902
rect 287114 -3462 287146 -3226
rect 287382 -3462 287466 -3226
rect 287702 -3462 287734 -3226
rect 287114 -3546 287734 -3462
rect 287114 -3782 287146 -3546
rect 287382 -3782 287466 -3546
rect 287702 -3782 287734 -3546
rect 287114 -3814 287734 -3782
rect 285714 -4422 285746 -4186
rect 285982 -4422 286066 -4186
rect 286302 -4422 286334 -4186
rect 285714 -4506 286334 -4422
rect 285714 -4742 285746 -4506
rect 285982 -4742 286066 -4506
rect 286302 -4742 286334 -4506
rect 285714 -5734 286334 -4742
rect 284314 -7302 284346 -7066
rect 284582 -7302 284666 -7066
rect 284902 -7302 284934 -7066
rect 284314 -7386 284934 -7302
rect 284314 -7622 284346 -7386
rect 284582 -7622 284666 -7386
rect 284902 -7622 284934 -7386
rect 284314 -7654 284934 -7622
rect 289434 -6106 290054 13000
rect 290834 -5146 291454 13000
rect 292234 7174 292854 13000
rect 292234 6938 292266 7174
rect 292502 6938 292586 7174
rect 292822 6938 292854 7174
rect 292234 6854 292854 6938
rect 292234 6618 292266 6854
rect 292502 6618 292586 6854
rect 292822 6618 292854 6854
rect 292234 -2266 292854 6618
rect 293634 -1306 294254 13000
rect 293634 -1542 293666 -1306
rect 293902 -1542 293986 -1306
rect 294222 -1542 294254 -1306
rect 293634 -1626 294254 -1542
rect 293634 -1862 293666 -1626
rect 293902 -1862 293986 -1626
rect 294222 -1862 294254 -1626
rect 293634 -1894 294254 -1862
rect 292234 -2502 292266 -2266
rect 292502 -2502 292586 -2266
rect 292822 -2502 292854 -2266
rect 292234 -2586 292854 -2502
rect 292234 -2822 292266 -2586
rect 292502 -2822 292586 -2586
rect 292822 -2822 292854 -2586
rect 292234 -3814 292854 -2822
rect 290834 -5382 290866 -5146
rect 291102 -5382 291186 -5146
rect 291422 -5382 291454 -5146
rect 290834 -5466 291454 -5382
rect 290834 -5702 290866 -5466
rect 291102 -5702 291186 -5466
rect 291422 -5702 291454 -5466
rect 290834 -5734 291454 -5702
rect 289434 -6342 289466 -6106
rect 289702 -6342 289786 -6106
rect 290022 -6342 290054 -6106
rect 289434 -6426 290054 -6342
rect 289434 -6662 289466 -6426
rect 289702 -6662 289786 -6426
rect 290022 -6662 290054 -6426
rect 289434 -7654 290054 -6662
rect 294554 -7066 295174 13000
rect 295954 10894 296574 13000
rect 295954 10658 295986 10894
rect 296222 10658 296306 10894
rect 296542 10658 296574 10894
rect 295954 10574 296574 10658
rect 295954 10338 295986 10574
rect 296222 10338 296306 10574
rect 296542 10338 296574 10574
rect 295954 -4186 296574 10338
rect 297354 -3226 297974 13000
rect 298754 3454 299374 13000
rect 298754 3218 298786 3454
rect 299022 3218 299106 3454
rect 299342 3218 299374 3454
rect 298754 3134 299374 3218
rect 298754 2898 298786 3134
rect 299022 2898 299106 3134
rect 299342 2898 299374 3134
rect 298754 -346 299374 2898
rect 298754 -582 298786 -346
rect 299022 -582 299106 -346
rect 299342 -582 299374 -346
rect 298754 -666 299374 -582
rect 298754 -902 298786 -666
rect 299022 -902 299106 -666
rect 299342 -902 299374 -666
rect 298754 -1894 299374 -902
rect 297354 -3462 297386 -3226
rect 297622 -3462 297706 -3226
rect 297942 -3462 297974 -3226
rect 297354 -3546 297974 -3462
rect 297354 -3782 297386 -3546
rect 297622 -3782 297706 -3546
rect 297942 -3782 297974 -3546
rect 297354 -3814 297974 -3782
rect 295954 -4422 295986 -4186
rect 296222 -4422 296306 -4186
rect 296542 -4422 296574 -4186
rect 295954 -4506 296574 -4422
rect 295954 -4742 295986 -4506
rect 296222 -4742 296306 -4506
rect 296542 -4742 296574 -4506
rect 295954 -5734 296574 -4742
rect 294554 -7302 294586 -7066
rect 294822 -7302 294906 -7066
rect 295142 -7302 295174 -7066
rect 294554 -7386 295174 -7302
rect 294554 -7622 294586 -7386
rect 294822 -7622 294906 -7386
rect 295142 -7622 295174 -7386
rect 294554 -7654 295174 -7622
rect 299674 -6106 300294 13000
rect 301074 -5146 301694 13000
rect 302474 7174 303094 13000
rect 302474 6938 302506 7174
rect 302742 6938 302826 7174
rect 303062 6938 303094 7174
rect 302474 6854 303094 6938
rect 302474 6618 302506 6854
rect 302742 6618 302826 6854
rect 303062 6618 303094 6854
rect 302474 -2266 303094 6618
rect 303874 -1306 304494 13000
rect 303874 -1542 303906 -1306
rect 304142 -1542 304226 -1306
rect 304462 -1542 304494 -1306
rect 303874 -1626 304494 -1542
rect 303874 -1862 303906 -1626
rect 304142 -1862 304226 -1626
rect 304462 -1862 304494 -1626
rect 303874 -1894 304494 -1862
rect 302474 -2502 302506 -2266
rect 302742 -2502 302826 -2266
rect 303062 -2502 303094 -2266
rect 302474 -2586 303094 -2502
rect 302474 -2822 302506 -2586
rect 302742 -2822 302826 -2586
rect 303062 -2822 303094 -2586
rect 302474 -3814 303094 -2822
rect 301074 -5382 301106 -5146
rect 301342 -5382 301426 -5146
rect 301662 -5382 301694 -5146
rect 301074 -5466 301694 -5382
rect 301074 -5702 301106 -5466
rect 301342 -5702 301426 -5466
rect 301662 -5702 301694 -5466
rect 301074 -5734 301694 -5702
rect 299674 -6342 299706 -6106
rect 299942 -6342 300026 -6106
rect 300262 -6342 300294 -6106
rect 299674 -6426 300294 -6342
rect 299674 -6662 299706 -6426
rect 299942 -6662 300026 -6426
rect 300262 -6662 300294 -6426
rect 299674 -7654 300294 -6662
rect 304794 -7066 305414 13000
rect 306194 10894 306814 13000
rect 306194 10658 306226 10894
rect 306462 10658 306546 10894
rect 306782 10658 306814 10894
rect 306194 10574 306814 10658
rect 306194 10338 306226 10574
rect 306462 10338 306546 10574
rect 306782 10338 306814 10574
rect 306194 -4186 306814 10338
rect 307594 -3226 308214 13000
rect 308994 3454 309614 13000
rect 308994 3218 309026 3454
rect 309262 3218 309346 3454
rect 309582 3218 309614 3454
rect 308994 3134 309614 3218
rect 308994 2898 309026 3134
rect 309262 2898 309346 3134
rect 309582 2898 309614 3134
rect 308994 -346 309614 2898
rect 308994 -582 309026 -346
rect 309262 -582 309346 -346
rect 309582 -582 309614 -346
rect 308994 -666 309614 -582
rect 308994 -902 309026 -666
rect 309262 -902 309346 -666
rect 309582 -902 309614 -666
rect 308994 -1894 309614 -902
rect 307594 -3462 307626 -3226
rect 307862 -3462 307946 -3226
rect 308182 -3462 308214 -3226
rect 307594 -3546 308214 -3462
rect 307594 -3782 307626 -3546
rect 307862 -3782 307946 -3546
rect 308182 -3782 308214 -3546
rect 307594 -3814 308214 -3782
rect 306194 -4422 306226 -4186
rect 306462 -4422 306546 -4186
rect 306782 -4422 306814 -4186
rect 306194 -4506 306814 -4422
rect 306194 -4742 306226 -4506
rect 306462 -4742 306546 -4506
rect 306782 -4742 306814 -4506
rect 306194 -5734 306814 -4742
rect 304794 -7302 304826 -7066
rect 305062 -7302 305146 -7066
rect 305382 -7302 305414 -7066
rect 304794 -7386 305414 -7302
rect 304794 -7622 304826 -7386
rect 305062 -7622 305146 -7386
rect 305382 -7622 305414 -7386
rect 304794 -7654 305414 -7622
rect 309914 -6106 310534 13000
rect 311314 -5146 311934 13000
rect 312714 7174 313334 13000
rect 312714 6938 312746 7174
rect 312982 6938 313066 7174
rect 313302 6938 313334 7174
rect 312714 6854 313334 6938
rect 312714 6618 312746 6854
rect 312982 6618 313066 6854
rect 313302 6618 313334 6854
rect 312714 -2266 313334 6618
rect 314114 -1306 314734 13000
rect 314114 -1542 314146 -1306
rect 314382 -1542 314466 -1306
rect 314702 -1542 314734 -1306
rect 314114 -1626 314734 -1542
rect 314114 -1862 314146 -1626
rect 314382 -1862 314466 -1626
rect 314702 -1862 314734 -1626
rect 314114 -1894 314734 -1862
rect 312714 -2502 312746 -2266
rect 312982 -2502 313066 -2266
rect 313302 -2502 313334 -2266
rect 312714 -2586 313334 -2502
rect 312714 -2822 312746 -2586
rect 312982 -2822 313066 -2586
rect 313302 -2822 313334 -2586
rect 312714 -3814 313334 -2822
rect 311314 -5382 311346 -5146
rect 311582 -5382 311666 -5146
rect 311902 -5382 311934 -5146
rect 311314 -5466 311934 -5382
rect 311314 -5702 311346 -5466
rect 311582 -5702 311666 -5466
rect 311902 -5702 311934 -5466
rect 311314 -5734 311934 -5702
rect 309914 -6342 309946 -6106
rect 310182 -6342 310266 -6106
rect 310502 -6342 310534 -6106
rect 309914 -6426 310534 -6342
rect 309914 -6662 309946 -6426
rect 310182 -6662 310266 -6426
rect 310502 -6662 310534 -6426
rect 309914 -7654 310534 -6662
rect 315034 -7066 315654 13000
rect 316434 10894 317054 13000
rect 316434 10658 316466 10894
rect 316702 10658 316786 10894
rect 317022 10658 317054 10894
rect 316434 10574 317054 10658
rect 316434 10338 316466 10574
rect 316702 10338 316786 10574
rect 317022 10338 317054 10574
rect 316434 -4186 317054 10338
rect 317834 -3226 318454 13000
rect 319234 3454 319854 13000
rect 319234 3218 319266 3454
rect 319502 3218 319586 3454
rect 319822 3218 319854 3454
rect 319234 3134 319854 3218
rect 319234 2898 319266 3134
rect 319502 2898 319586 3134
rect 319822 2898 319854 3134
rect 319234 -346 319854 2898
rect 319234 -582 319266 -346
rect 319502 -582 319586 -346
rect 319822 -582 319854 -346
rect 319234 -666 319854 -582
rect 319234 -902 319266 -666
rect 319502 -902 319586 -666
rect 319822 -902 319854 -666
rect 319234 -1894 319854 -902
rect 317834 -3462 317866 -3226
rect 318102 -3462 318186 -3226
rect 318422 -3462 318454 -3226
rect 317834 -3546 318454 -3462
rect 317834 -3782 317866 -3546
rect 318102 -3782 318186 -3546
rect 318422 -3782 318454 -3546
rect 317834 -3814 318454 -3782
rect 316434 -4422 316466 -4186
rect 316702 -4422 316786 -4186
rect 317022 -4422 317054 -4186
rect 316434 -4506 317054 -4422
rect 316434 -4742 316466 -4506
rect 316702 -4742 316786 -4506
rect 317022 -4742 317054 -4506
rect 316434 -5734 317054 -4742
rect 315034 -7302 315066 -7066
rect 315302 -7302 315386 -7066
rect 315622 -7302 315654 -7066
rect 315034 -7386 315654 -7302
rect 315034 -7622 315066 -7386
rect 315302 -7622 315386 -7386
rect 315622 -7622 315654 -7386
rect 315034 -7654 315654 -7622
rect 320154 -6106 320774 13000
rect 321554 -5146 322174 13000
rect 322954 7174 323574 13000
rect 322954 6938 322986 7174
rect 323222 6938 323306 7174
rect 323542 6938 323574 7174
rect 322954 6854 323574 6938
rect 322954 6618 322986 6854
rect 323222 6618 323306 6854
rect 323542 6618 323574 6854
rect 322954 -2266 323574 6618
rect 324354 -1306 324974 13000
rect 324354 -1542 324386 -1306
rect 324622 -1542 324706 -1306
rect 324942 -1542 324974 -1306
rect 324354 -1626 324974 -1542
rect 324354 -1862 324386 -1626
rect 324622 -1862 324706 -1626
rect 324942 -1862 324974 -1626
rect 324354 -1894 324974 -1862
rect 322954 -2502 322986 -2266
rect 323222 -2502 323306 -2266
rect 323542 -2502 323574 -2266
rect 322954 -2586 323574 -2502
rect 322954 -2822 322986 -2586
rect 323222 -2822 323306 -2586
rect 323542 -2822 323574 -2586
rect 322954 -3814 323574 -2822
rect 321554 -5382 321586 -5146
rect 321822 -5382 321906 -5146
rect 322142 -5382 322174 -5146
rect 321554 -5466 322174 -5382
rect 321554 -5702 321586 -5466
rect 321822 -5702 321906 -5466
rect 322142 -5702 322174 -5466
rect 321554 -5734 322174 -5702
rect 320154 -6342 320186 -6106
rect 320422 -6342 320506 -6106
rect 320742 -6342 320774 -6106
rect 320154 -6426 320774 -6342
rect 320154 -6662 320186 -6426
rect 320422 -6662 320506 -6426
rect 320742 -6662 320774 -6426
rect 320154 -7654 320774 -6662
rect 325274 -7066 325894 13000
rect 326674 10894 327294 13000
rect 326674 10658 326706 10894
rect 326942 10658 327026 10894
rect 327262 10658 327294 10894
rect 326674 10574 327294 10658
rect 326674 10338 326706 10574
rect 326942 10338 327026 10574
rect 327262 10338 327294 10574
rect 326674 -4186 327294 10338
rect 328074 -3226 328694 13000
rect 329474 3454 330094 13000
rect 329474 3218 329506 3454
rect 329742 3218 329826 3454
rect 330062 3218 330094 3454
rect 329474 3134 330094 3218
rect 329474 2898 329506 3134
rect 329742 2898 329826 3134
rect 330062 2898 330094 3134
rect 329474 -346 330094 2898
rect 329474 -582 329506 -346
rect 329742 -582 329826 -346
rect 330062 -582 330094 -346
rect 329474 -666 330094 -582
rect 329474 -902 329506 -666
rect 329742 -902 329826 -666
rect 330062 -902 330094 -666
rect 329474 -1894 330094 -902
rect 328074 -3462 328106 -3226
rect 328342 -3462 328426 -3226
rect 328662 -3462 328694 -3226
rect 328074 -3546 328694 -3462
rect 328074 -3782 328106 -3546
rect 328342 -3782 328426 -3546
rect 328662 -3782 328694 -3546
rect 328074 -3814 328694 -3782
rect 326674 -4422 326706 -4186
rect 326942 -4422 327026 -4186
rect 327262 -4422 327294 -4186
rect 326674 -4506 327294 -4422
rect 326674 -4742 326706 -4506
rect 326942 -4742 327026 -4506
rect 327262 -4742 327294 -4506
rect 326674 -5734 327294 -4742
rect 325274 -7302 325306 -7066
rect 325542 -7302 325626 -7066
rect 325862 -7302 325894 -7066
rect 325274 -7386 325894 -7302
rect 325274 -7622 325306 -7386
rect 325542 -7622 325626 -7386
rect 325862 -7622 325894 -7386
rect 325274 -7654 325894 -7622
rect 330394 -6106 331014 13000
rect 331794 -5146 332414 13000
rect 333194 7174 333814 13000
rect 333194 6938 333226 7174
rect 333462 6938 333546 7174
rect 333782 6938 333814 7174
rect 333194 6854 333814 6938
rect 333194 6618 333226 6854
rect 333462 6618 333546 6854
rect 333782 6618 333814 6854
rect 333194 -2266 333814 6618
rect 334594 -1306 335214 13000
rect 334594 -1542 334626 -1306
rect 334862 -1542 334946 -1306
rect 335182 -1542 335214 -1306
rect 334594 -1626 335214 -1542
rect 334594 -1862 334626 -1626
rect 334862 -1862 334946 -1626
rect 335182 -1862 335214 -1626
rect 334594 -1894 335214 -1862
rect 333194 -2502 333226 -2266
rect 333462 -2502 333546 -2266
rect 333782 -2502 333814 -2266
rect 333194 -2586 333814 -2502
rect 333194 -2822 333226 -2586
rect 333462 -2822 333546 -2586
rect 333782 -2822 333814 -2586
rect 333194 -3814 333814 -2822
rect 331794 -5382 331826 -5146
rect 332062 -5382 332146 -5146
rect 332382 -5382 332414 -5146
rect 331794 -5466 332414 -5382
rect 331794 -5702 331826 -5466
rect 332062 -5702 332146 -5466
rect 332382 -5702 332414 -5466
rect 331794 -5734 332414 -5702
rect 330394 -6342 330426 -6106
rect 330662 -6342 330746 -6106
rect 330982 -6342 331014 -6106
rect 330394 -6426 331014 -6342
rect 330394 -6662 330426 -6426
rect 330662 -6662 330746 -6426
rect 330982 -6662 331014 -6426
rect 330394 -7654 331014 -6662
rect 335514 -7066 336134 13000
rect 336914 10894 337534 13000
rect 336914 10658 336946 10894
rect 337182 10658 337266 10894
rect 337502 10658 337534 10894
rect 336914 10574 337534 10658
rect 336914 10338 336946 10574
rect 337182 10338 337266 10574
rect 337502 10338 337534 10574
rect 336914 -4186 337534 10338
rect 338314 -3226 338934 13000
rect 339714 3454 340334 13000
rect 339714 3218 339746 3454
rect 339982 3218 340066 3454
rect 340302 3218 340334 3454
rect 339714 3134 340334 3218
rect 339714 2898 339746 3134
rect 339982 2898 340066 3134
rect 340302 2898 340334 3134
rect 339714 -346 340334 2898
rect 339714 -582 339746 -346
rect 339982 -582 340066 -346
rect 340302 -582 340334 -346
rect 339714 -666 340334 -582
rect 339714 -902 339746 -666
rect 339982 -902 340066 -666
rect 340302 -902 340334 -666
rect 339714 -1894 340334 -902
rect 338314 -3462 338346 -3226
rect 338582 -3462 338666 -3226
rect 338902 -3462 338934 -3226
rect 338314 -3546 338934 -3462
rect 338314 -3782 338346 -3546
rect 338582 -3782 338666 -3546
rect 338902 -3782 338934 -3546
rect 338314 -3814 338934 -3782
rect 336914 -4422 336946 -4186
rect 337182 -4422 337266 -4186
rect 337502 -4422 337534 -4186
rect 336914 -4506 337534 -4422
rect 336914 -4742 336946 -4506
rect 337182 -4742 337266 -4506
rect 337502 -4742 337534 -4506
rect 336914 -5734 337534 -4742
rect 335514 -7302 335546 -7066
rect 335782 -7302 335866 -7066
rect 336102 -7302 336134 -7066
rect 335514 -7386 336134 -7302
rect 335514 -7622 335546 -7386
rect 335782 -7622 335866 -7386
rect 336102 -7622 336134 -7386
rect 335514 -7654 336134 -7622
rect 340634 -6106 341254 13000
rect 342034 -5146 342654 13000
rect 343434 7174 344054 13000
rect 343434 6938 343466 7174
rect 343702 6938 343786 7174
rect 344022 6938 344054 7174
rect 343434 6854 344054 6938
rect 343434 6618 343466 6854
rect 343702 6618 343786 6854
rect 344022 6618 344054 6854
rect 343434 -2266 344054 6618
rect 344834 -1306 345454 13000
rect 344834 -1542 344866 -1306
rect 345102 -1542 345186 -1306
rect 345422 -1542 345454 -1306
rect 344834 -1626 345454 -1542
rect 344834 -1862 344866 -1626
rect 345102 -1862 345186 -1626
rect 345422 -1862 345454 -1626
rect 344834 -1894 345454 -1862
rect 343434 -2502 343466 -2266
rect 343702 -2502 343786 -2266
rect 344022 -2502 344054 -2266
rect 343434 -2586 344054 -2502
rect 343434 -2822 343466 -2586
rect 343702 -2822 343786 -2586
rect 344022 -2822 344054 -2586
rect 343434 -3814 344054 -2822
rect 342034 -5382 342066 -5146
rect 342302 -5382 342386 -5146
rect 342622 -5382 342654 -5146
rect 342034 -5466 342654 -5382
rect 342034 -5702 342066 -5466
rect 342302 -5702 342386 -5466
rect 342622 -5702 342654 -5466
rect 342034 -5734 342654 -5702
rect 340634 -6342 340666 -6106
rect 340902 -6342 340986 -6106
rect 341222 -6342 341254 -6106
rect 340634 -6426 341254 -6342
rect 340634 -6662 340666 -6426
rect 340902 -6662 340986 -6426
rect 341222 -6662 341254 -6426
rect 340634 -7654 341254 -6662
rect 345754 -7066 346374 13000
rect 347154 10894 347774 13000
rect 347154 10658 347186 10894
rect 347422 10658 347506 10894
rect 347742 10658 347774 10894
rect 347154 10574 347774 10658
rect 347154 10338 347186 10574
rect 347422 10338 347506 10574
rect 347742 10338 347774 10574
rect 347154 -4186 347774 10338
rect 348554 -3226 349174 13000
rect 349954 3454 350574 13000
rect 349954 3218 349986 3454
rect 350222 3218 350306 3454
rect 350542 3218 350574 3454
rect 349954 3134 350574 3218
rect 349954 2898 349986 3134
rect 350222 2898 350306 3134
rect 350542 2898 350574 3134
rect 349954 -346 350574 2898
rect 349954 -582 349986 -346
rect 350222 -582 350306 -346
rect 350542 -582 350574 -346
rect 349954 -666 350574 -582
rect 349954 -902 349986 -666
rect 350222 -902 350306 -666
rect 350542 -902 350574 -666
rect 349954 -1894 350574 -902
rect 348554 -3462 348586 -3226
rect 348822 -3462 348906 -3226
rect 349142 -3462 349174 -3226
rect 348554 -3546 349174 -3462
rect 348554 -3782 348586 -3546
rect 348822 -3782 348906 -3546
rect 349142 -3782 349174 -3546
rect 348554 -3814 349174 -3782
rect 347154 -4422 347186 -4186
rect 347422 -4422 347506 -4186
rect 347742 -4422 347774 -4186
rect 347154 -4506 347774 -4422
rect 347154 -4742 347186 -4506
rect 347422 -4742 347506 -4506
rect 347742 -4742 347774 -4506
rect 347154 -5734 347774 -4742
rect 345754 -7302 345786 -7066
rect 346022 -7302 346106 -7066
rect 346342 -7302 346374 -7066
rect 345754 -7386 346374 -7302
rect 345754 -7622 345786 -7386
rect 346022 -7622 346106 -7386
rect 346342 -7622 346374 -7386
rect 345754 -7654 346374 -7622
rect 350874 -6106 351494 13000
rect 352274 -5146 352894 13000
rect 353674 7174 354294 13000
rect 353674 6938 353706 7174
rect 353942 6938 354026 7174
rect 354262 6938 354294 7174
rect 353674 6854 354294 6938
rect 353674 6618 353706 6854
rect 353942 6618 354026 6854
rect 354262 6618 354294 6854
rect 353674 -2266 354294 6618
rect 355074 -1306 355694 13000
rect 355074 -1542 355106 -1306
rect 355342 -1542 355426 -1306
rect 355662 -1542 355694 -1306
rect 355074 -1626 355694 -1542
rect 355074 -1862 355106 -1626
rect 355342 -1862 355426 -1626
rect 355662 -1862 355694 -1626
rect 355074 -1894 355694 -1862
rect 353674 -2502 353706 -2266
rect 353942 -2502 354026 -2266
rect 354262 -2502 354294 -2266
rect 353674 -2586 354294 -2502
rect 353674 -2822 353706 -2586
rect 353942 -2822 354026 -2586
rect 354262 -2822 354294 -2586
rect 353674 -3814 354294 -2822
rect 352274 -5382 352306 -5146
rect 352542 -5382 352626 -5146
rect 352862 -5382 352894 -5146
rect 352274 -5466 352894 -5382
rect 352274 -5702 352306 -5466
rect 352542 -5702 352626 -5466
rect 352862 -5702 352894 -5466
rect 352274 -5734 352894 -5702
rect 350874 -6342 350906 -6106
rect 351142 -6342 351226 -6106
rect 351462 -6342 351494 -6106
rect 350874 -6426 351494 -6342
rect 350874 -6662 350906 -6426
rect 351142 -6662 351226 -6426
rect 351462 -6662 351494 -6426
rect 350874 -7654 351494 -6662
rect 355994 -7066 356614 13000
rect 357394 10894 358014 13000
rect 357394 10658 357426 10894
rect 357662 10658 357746 10894
rect 357982 10658 358014 10894
rect 357394 10574 358014 10658
rect 357394 10338 357426 10574
rect 357662 10338 357746 10574
rect 357982 10338 358014 10574
rect 357394 -4186 358014 10338
rect 358794 -3226 359414 13000
rect 360194 3454 360814 13000
rect 360194 3218 360226 3454
rect 360462 3218 360546 3454
rect 360782 3218 360814 3454
rect 360194 3134 360814 3218
rect 360194 2898 360226 3134
rect 360462 2898 360546 3134
rect 360782 2898 360814 3134
rect 360194 -346 360814 2898
rect 360194 -582 360226 -346
rect 360462 -582 360546 -346
rect 360782 -582 360814 -346
rect 360194 -666 360814 -582
rect 360194 -902 360226 -666
rect 360462 -902 360546 -666
rect 360782 -902 360814 -666
rect 360194 -1894 360814 -902
rect 358794 -3462 358826 -3226
rect 359062 -3462 359146 -3226
rect 359382 -3462 359414 -3226
rect 358794 -3546 359414 -3462
rect 358794 -3782 358826 -3546
rect 359062 -3782 359146 -3546
rect 359382 -3782 359414 -3546
rect 358794 -3814 359414 -3782
rect 357394 -4422 357426 -4186
rect 357662 -4422 357746 -4186
rect 357982 -4422 358014 -4186
rect 357394 -4506 358014 -4422
rect 357394 -4742 357426 -4506
rect 357662 -4742 357746 -4506
rect 357982 -4742 358014 -4506
rect 357394 -5734 358014 -4742
rect 355994 -7302 356026 -7066
rect 356262 -7302 356346 -7066
rect 356582 -7302 356614 -7066
rect 355994 -7386 356614 -7302
rect 355994 -7622 356026 -7386
rect 356262 -7622 356346 -7386
rect 356582 -7622 356614 -7386
rect 355994 -7654 356614 -7622
rect 361114 -6106 361734 13000
rect 362514 -5146 363134 13000
rect 363914 7174 364534 13000
rect 363914 6938 363946 7174
rect 364182 6938 364266 7174
rect 364502 6938 364534 7174
rect 363914 6854 364534 6938
rect 363914 6618 363946 6854
rect 364182 6618 364266 6854
rect 364502 6618 364534 6854
rect 363914 -2266 364534 6618
rect 365314 -1306 365934 13000
rect 365314 -1542 365346 -1306
rect 365582 -1542 365666 -1306
rect 365902 -1542 365934 -1306
rect 365314 -1626 365934 -1542
rect 365314 -1862 365346 -1626
rect 365582 -1862 365666 -1626
rect 365902 -1862 365934 -1626
rect 365314 -1894 365934 -1862
rect 363914 -2502 363946 -2266
rect 364182 -2502 364266 -2266
rect 364502 -2502 364534 -2266
rect 363914 -2586 364534 -2502
rect 363914 -2822 363946 -2586
rect 364182 -2822 364266 -2586
rect 364502 -2822 364534 -2586
rect 363914 -3814 364534 -2822
rect 362514 -5382 362546 -5146
rect 362782 -5382 362866 -5146
rect 363102 -5382 363134 -5146
rect 362514 -5466 363134 -5382
rect 362514 -5702 362546 -5466
rect 362782 -5702 362866 -5466
rect 363102 -5702 363134 -5466
rect 362514 -5734 363134 -5702
rect 361114 -6342 361146 -6106
rect 361382 -6342 361466 -6106
rect 361702 -6342 361734 -6106
rect 361114 -6426 361734 -6342
rect 361114 -6662 361146 -6426
rect 361382 -6662 361466 -6426
rect 361702 -6662 361734 -6426
rect 361114 -7654 361734 -6662
rect 366234 -7066 366854 13000
rect 367634 10894 368254 13000
rect 367634 10658 367666 10894
rect 367902 10658 367986 10894
rect 368222 10658 368254 10894
rect 367634 10574 368254 10658
rect 367634 10338 367666 10574
rect 367902 10338 367986 10574
rect 368222 10338 368254 10574
rect 367634 -4186 368254 10338
rect 369034 -3226 369654 13000
rect 370434 3454 371054 13000
rect 370434 3218 370466 3454
rect 370702 3218 370786 3454
rect 371022 3218 371054 3454
rect 370434 3134 371054 3218
rect 370434 2898 370466 3134
rect 370702 2898 370786 3134
rect 371022 2898 371054 3134
rect 370434 -346 371054 2898
rect 370434 -582 370466 -346
rect 370702 -582 370786 -346
rect 371022 -582 371054 -346
rect 370434 -666 371054 -582
rect 370434 -902 370466 -666
rect 370702 -902 370786 -666
rect 371022 -902 371054 -666
rect 370434 -1894 371054 -902
rect 369034 -3462 369066 -3226
rect 369302 -3462 369386 -3226
rect 369622 -3462 369654 -3226
rect 369034 -3546 369654 -3462
rect 369034 -3782 369066 -3546
rect 369302 -3782 369386 -3546
rect 369622 -3782 369654 -3546
rect 369034 -3814 369654 -3782
rect 367634 -4422 367666 -4186
rect 367902 -4422 367986 -4186
rect 368222 -4422 368254 -4186
rect 367634 -4506 368254 -4422
rect 367634 -4742 367666 -4506
rect 367902 -4742 367986 -4506
rect 368222 -4742 368254 -4506
rect 367634 -5734 368254 -4742
rect 366234 -7302 366266 -7066
rect 366502 -7302 366586 -7066
rect 366822 -7302 366854 -7066
rect 366234 -7386 366854 -7302
rect 366234 -7622 366266 -7386
rect 366502 -7622 366586 -7386
rect 366822 -7622 366854 -7386
rect 366234 -7654 366854 -7622
rect 371354 -6106 371974 13000
rect 372754 -5146 373374 13000
rect 374154 7174 374774 13000
rect 374154 6938 374186 7174
rect 374422 6938 374506 7174
rect 374742 6938 374774 7174
rect 374154 6854 374774 6938
rect 374154 6618 374186 6854
rect 374422 6618 374506 6854
rect 374742 6618 374774 6854
rect 374154 -2266 374774 6618
rect 375554 -1306 376174 13000
rect 375554 -1542 375586 -1306
rect 375822 -1542 375906 -1306
rect 376142 -1542 376174 -1306
rect 375554 -1626 376174 -1542
rect 375554 -1862 375586 -1626
rect 375822 -1862 375906 -1626
rect 376142 -1862 376174 -1626
rect 375554 -1894 376174 -1862
rect 374154 -2502 374186 -2266
rect 374422 -2502 374506 -2266
rect 374742 -2502 374774 -2266
rect 374154 -2586 374774 -2502
rect 374154 -2822 374186 -2586
rect 374422 -2822 374506 -2586
rect 374742 -2822 374774 -2586
rect 374154 -3814 374774 -2822
rect 372754 -5382 372786 -5146
rect 373022 -5382 373106 -5146
rect 373342 -5382 373374 -5146
rect 372754 -5466 373374 -5382
rect 372754 -5702 372786 -5466
rect 373022 -5702 373106 -5466
rect 373342 -5702 373374 -5466
rect 372754 -5734 373374 -5702
rect 371354 -6342 371386 -6106
rect 371622 -6342 371706 -6106
rect 371942 -6342 371974 -6106
rect 371354 -6426 371974 -6342
rect 371354 -6662 371386 -6426
rect 371622 -6662 371706 -6426
rect 371942 -6662 371974 -6426
rect 371354 -7654 371974 -6662
rect 376474 -7066 377094 13000
rect 377874 10894 378494 13000
rect 377874 10658 377906 10894
rect 378142 10658 378226 10894
rect 378462 10658 378494 10894
rect 377874 10574 378494 10658
rect 377874 10338 377906 10574
rect 378142 10338 378226 10574
rect 378462 10338 378494 10574
rect 377874 -4186 378494 10338
rect 379274 -3226 379894 13000
rect 380674 3454 381294 13000
rect 380674 3218 380706 3454
rect 380942 3218 381026 3454
rect 381262 3218 381294 3454
rect 380674 3134 381294 3218
rect 380674 2898 380706 3134
rect 380942 2898 381026 3134
rect 381262 2898 381294 3134
rect 380674 -346 381294 2898
rect 380674 -582 380706 -346
rect 380942 -582 381026 -346
rect 381262 -582 381294 -346
rect 380674 -666 381294 -582
rect 380674 -902 380706 -666
rect 380942 -902 381026 -666
rect 381262 -902 381294 -666
rect 380674 -1894 381294 -902
rect 379274 -3462 379306 -3226
rect 379542 -3462 379626 -3226
rect 379862 -3462 379894 -3226
rect 379274 -3546 379894 -3462
rect 379274 -3782 379306 -3546
rect 379542 -3782 379626 -3546
rect 379862 -3782 379894 -3546
rect 379274 -3814 379894 -3782
rect 377874 -4422 377906 -4186
rect 378142 -4422 378226 -4186
rect 378462 -4422 378494 -4186
rect 377874 -4506 378494 -4422
rect 377874 -4742 377906 -4506
rect 378142 -4742 378226 -4506
rect 378462 -4742 378494 -4506
rect 377874 -5734 378494 -4742
rect 376474 -7302 376506 -7066
rect 376742 -7302 376826 -7066
rect 377062 -7302 377094 -7066
rect 376474 -7386 377094 -7302
rect 376474 -7622 376506 -7386
rect 376742 -7622 376826 -7386
rect 377062 -7622 377094 -7386
rect 376474 -7654 377094 -7622
rect 381594 -6106 382214 13000
rect 382994 -5146 383614 13000
rect 384394 7174 385014 13000
rect 384394 6938 384426 7174
rect 384662 6938 384746 7174
rect 384982 6938 385014 7174
rect 384394 6854 385014 6938
rect 384394 6618 384426 6854
rect 384662 6618 384746 6854
rect 384982 6618 385014 6854
rect 384394 -2266 385014 6618
rect 385794 -1306 386414 13000
rect 385794 -1542 385826 -1306
rect 386062 -1542 386146 -1306
rect 386382 -1542 386414 -1306
rect 385794 -1626 386414 -1542
rect 385794 -1862 385826 -1626
rect 386062 -1862 386146 -1626
rect 386382 -1862 386414 -1626
rect 385794 -1894 386414 -1862
rect 384394 -2502 384426 -2266
rect 384662 -2502 384746 -2266
rect 384982 -2502 385014 -2266
rect 384394 -2586 385014 -2502
rect 384394 -2822 384426 -2586
rect 384662 -2822 384746 -2586
rect 384982 -2822 385014 -2586
rect 384394 -3814 385014 -2822
rect 382994 -5382 383026 -5146
rect 383262 -5382 383346 -5146
rect 383582 -5382 383614 -5146
rect 382994 -5466 383614 -5382
rect 382994 -5702 383026 -5466
rect 383262 -5702 383346 -5466
rect 383582 -5702 383614 -5466
rect 382994 -5734 383614 -5702
rect 381594 -6342 381626 -6106
rect 381862 -6342 381946 -6106
rect 382182 -6342 382214 -6106
rect 381594 -6426 382214 -6342
rect 381594 -6662 381626 -6426
rect 381862 -6662 381946 -6426
rect 382182 -6662 382214 -6426
rect 381594 -7654 382214 -6662
rect 386714 -7066 387334 13000
rect 388114 10894 388734 13000
rect 388114 10658 388146 10894
rect 388382 10658 388466 10894
rect 388702 10658 388734 10894
rect 388114 10574 388734 10658
rect 388114 10338 388146 10574
rect 388382 10338 388466 10574
rect 388702 10338 388734 10574
rect 388114 -4186 388734 10338
rect 389514 -3226 390134 13000
rect 390914 3454 391534 13000
rect 390914 3218 390946 3454
rect 391182 3218 391266 3454
rect 391502 3218 391534 3454
rect 390914 3134 391534 3218
rect 390914 2898 390946 3134
rect 391182 2898 391266 3134
rect 391502 2898 391534 3134
rect 390914 -346 391534 2898
rect 390914 -582 390946 -346
rect 391182 -582 391266 -346
rect 391502 -582 391534 -346
rect 390914 -666 391534 -582
rect 390914 -902 390946 -666
rect 391182 -902 391266 -666
rect 391502 -902 391534 -666
rect 390914 -1894 391534 -902
rect 389514 -3462 389546 -3226
rect 389782 -3462 389866 -3226
rect 390102 -3462 390134 -3226
rect 389514 -3546 390134 -3462
rect 389514 -3782 389546 -3546
rect 389782 -3782 389866 -3546
rect 390102 -3782 390134 -3546
rect 389514 -3814 390134 -3782
rect 388114 -4422 388146 -4186
rect 388382 -4422 388466 -4186
rect 388702 -4422 388734 -4186
rect 388114 -4506 388734 -4422
rect 388114 -4742 388146 -4506
rect 388382 -4742 388466 -4506
rect 388702 -4742 388734 -4506
rect 388114 -5734 388734 -4742
rect 386714 -7302 386746 -7066
rect 386982 -7302 387066 -7066
rect 387302 -7302 387334 -7066
rect 386714 -7386 387334 -7302
rect 386714 -7622 386746 -7386
rect 386982 -7622 387066 -7386
rect 387302 -7622 387334 -7386
rect 386714 -7654 387334 -7622
rect 391834 -6106 392454 13000
rect 393234 -5146 393854 13000
rect 394634 7174 395254 13000
rect 394634 6938 394666 7174
rect 394902 6938 394986 7174
rect 395222 6938 395254 7174
rect 394634 6854 395254 6938
rect 394634 6618 394666 6854
rect 394902 6618 394986 6854
rect 395222 6618 395254 6854
rect 394634 -2266 395254 6618
rect 396034 -1306 396654 13000
rect 396034 -1542 396066 -1306
rect 396302 -1542 396386 -1306
rect 396622 -1542 396654 -1306
rect 396034 -1626 396654 -1542
rect 396034 -1862 396066 -1626
rect 396302 -1862 396386 -1626
rect 396622 -1862 396654 -1626
rect 396034 -1894 396654 -1862
rect 394634 -2502 394666 -2266
rect 394902 -2502 394986 -2266
rect 395222 -2502 395254 -2266
rect 394634 -2586 395254 -2502
rect 394634 -2822 394666 -2586
rect 394902 -2822 394986 -2586
rect 395222 -2822 395254 -2586
rect 394634 -3814 395254 -2822
rect 393234 -5382 393266 -5146
rect 393502 -5382 393586 -5146
rect 393822 -5382 393854 -5146
rect 393234 -5466 393854 -5382
rect 393234 -5702 393266 -5466
rect 393502 -5702 393586 -5466
rect 393822 -5702 393854 -5466
rect 393234 -5734 393854 -5702
rect 391834 -6342 391866 -6106
rect 392102 -6342 392186 -6106
rect 392422 -6342 392454 -6106
rect 391834 -6426 392454 -6342
rect 391834 -6662 391866 -6426
rect 392102 -6662 392186 -6426
rect 392422 -6662 392454 -6426
rect 391834 -7654 392454 -6662
rect 396954 -7066 397574 13000
rect 398354 10894 398974 13000
rect 398354 10658 398386 10894
rect 398622 10658 398706 10894
rect 398942 10658 398974 10894
rect 398354 10574 398974 10658
rect 398354 10338 398386 10574
rect 398622 10338 398706 10574
rect 398942 10338 398974 10574
rect 398354 -4186 398974 10338
rect 399754 -3226 400374 13000
rect 401154 3454 401774 13000
rect 401154 3218 401186 3454
rect 401422 3218 401506 3454
rect 401742 3218 401774 3454
rect 401154 3134 401774 3218
rect 401154 2898 401186 3134
rect 401422 2898 401506 3134
rect 401742 2898 401774 3134
rect 401154 -346 401774 2898
rect 401154 -582 401186 -346
rect 401422 -582 401506 -346
rect 401742 -582 401774 -346
rect 401154 -666 401774 -582
rect 401154 -902 401186 -666
rect 401422 -902 401506 -666
rect 401742 -902 401774 -666
rect 401154 -1894 401774 -902
rect 399754 -3462 399786 -3226
rect 400022 -3462 400106 -3226
rect 400342 -3462 400374 -3226
rect 399754 -3546 400374 -3462
rect 399754 -3782 399786 -3546
rect 400022 -3782 400106 -3546
rect 400342 -3782 400374 -3546
rect 399754 -3814 400374 -3782
rect 398354 -4422 398386 -4186
rect 398622 -4422 398706 -4186
rect 398942 -4422 398974 -4186
rect 398354 -4506 398974 -4422
rect 398354 -4742 398386 -4506
rect 398622 -4742 398706 -4506
rect 398942 -4742 398974 -4506
rect 398354 -5734 398974 -4742
rect 396954 -7302 396986 -7066
rect 397222 -7302 397306 -7066
rect 397542 -7302 397574 -7066
rect 396954 -7386 397574 -7302
rect 396954 -7622 396986 -7386
rect 397222 -7622 397306 -7386
rect 397542 -7622 397574 -7386
rect 396954 -7654 397574 -7622
rect 402074 -6106 402694 13000
rect 403474 -5146 404094 13000
rect 404874 7174 405494 13000
rect 404874 6938 404906 7174
rect 405142 6938 405226 7174
rect 405462 6938 405494 7174
rect 404874 6854 405494 6938
rect 404874 6618 404906 6854
rect 405142 6618 405226 6854
rect 405462 6618 405494 6854
rect 404874 -2266 405494 6618
rect 406274 -1306 406894 13000
rect 406274 -1542 406306 -1306
rect 406542 -1542 406626 -1306
rect 406862 -1542 406894 -1306
rect 406274 -1626 406894 -1542
rect 406274 -1862 406306 -1626
rect 406542 -1862 406626 -1626
rect 406862 -1862 406894 -1626
rect 406274 -1894 406894 -1862
rect 404874 -2502 404906 -2266
rect 405142 -2502 405226 -2266
rect 405462 -2502 405494 -2266
rect 404874 -2586 405494 -2502
rect 404874 -2822 404906 -2586
rect 405142 -2822 405226 -2586
rect 405462 -2822 405494 -2586
rect 404874 -3814 405494 -2822
rect 403474 -5382 403506 -5146
rect 403742 -5382 403826 -5146
rect 404062 -5382 404094 -5146
rect 403474 -5466 404094 -5382
rect 403474 -5702 403506 -5466
rect 403742 -5702 403826 -5466
rect 404062 -5702 404094 -5466
rect 403474 -5734 404094 -5702
rect 402074 -6342 402106 -6106
rect 402342 -6342 402426 -6106
rect 402662 -6342 402694 -6106
rect 402074 -6426 402694 -6342
rect 402074 -6662 402106 -6426
rect 402342 -6662 402426 -6426
rect 402662 -6662 402694 -6426
rect 402074 -7654 402694 -6662
rect 407194 -7066 407814 13000
rect 408594 10894 409214 13000
rect 408594 10658 408626 10894
rect 408862 10658 408946 10894
rect 409182 10658 409214 10894
rect 408594 10574 409214 10658
rect 408594 10338 408626 10574
rect 408862 10338 408946 10574
rect 409182 10338 409214 10574
rect 408594 -4186 409214 10338
rect 409994 -3226 410614 13000
rect 411394 3454 412014 13000
rect 411394 3218 411426 3454
rect 411662 3218 411746 3454
rect 411982 3218 412014 3454
rect 411394 3134 412014 3218
rect 411394 2898 411426 3134
rect 411662 2898 411746 3134
rect 411982 2898 412014 3134
rect 411394 -346 412014 2898
rect 411394 -582 411426 -346
rect 411662 -582 411746 -346
rect 411982 -582 412014 -346
rect 411394 -666 412014 -582
rect 411394 -902 411426 -666
rect 411662 -902 411746 -666
rect 411982 -902 412014 -666
rect 411394 -1894 412014 -902
rect 409994 -3462 410026 -3226
rect 410262 -3462 410346 -3226
rect 410582 -3462 410614 -3226
rect 409994 -3546 410614 -3462
rect 409994 -3782 410026 -3546
rect 410262 -3782 410346 -3546
rect 410582 -3782 410614 -3546
rect 409994 -3814 410614 -3782
rect 408594 -4422 408626 -4186
rect 408862 -4422 408946 -4186
rect 409182 -4422 409214 -4186
rect 408594 -4506 409214 -4422
rect 408594 -4742 408626 -4506
rect 408862 -4742 408946 -4506
rect 409182 -4742 409214 -4506
rect 408594 -5734 409214 -4742
rect 407194 -7302 407226 -7066
rect 407462 -7302 407546 -7066
rect 407782 -7302 407814 -7066
rect 407194 -7386 407814 -7302
rect 407194 -7622 407226 -7386
rect 407462 -7622 407546 -7386
rect 407782 -7622 407814 -7386
rect 407194 -7654 407814 -7622
rect 412314 -6106 412934 13000
rect 413714 -5146 414334 13000
rect 415114 7174 415734 13000
rect 415114 6938 415146 7174
rect 415382 6938 415466 7174
rect 415702 6938 415734 7174
rect 415114 6854 415734 6938
rect 415114 6618 415146 6854
rect 415382 6618 415466 6854
rect 415702 6618 415734 6854
rect 415114 -2266 415734 6618
rect 416514 -1306 417134 13000
rect 416514 -1542 416546 -1306
rect 416782 -1542 416866 -1306
rect 417102 -1542 417134 -1306
rect 416514 -1626 417134 -1542
rect 416514 -1862 416546 -1626
rect 416782 -1862 416866 -1626
rect 417102 -1862 417134 -1626
rect 416514 -1894 417134 -1862
rect 415114 -2502 415146 -2266
rect 415382 -2502 415466 -2266
rect 415702 -2502 415734 -2266
rect 415114 -2586 415734 -2502
rect 415114 -2822 415146 -2586
rect 415382 -2822 415466 -2586
rect 415702 -2822 415734 -2586
rect 415114 -3814 415734 -2822
rect 413714 -5382 413746 -5146
rect 413982 -5382 414066 -5146
rect 414302 -5382 414334 -5146
rect 413714 -5466 414334 -5382
rect 413714 -5702 413746 -5466
rect 413982 -5702 414066 -5466
rect 414302 -5702 414334 -5466
rect 413714 -5734 414334 -5702
rect 412314 -6342 412346 -6106
rect 412582 -6342 412666 -6106
rect 412902 -6342 412934 -6106
rect 412314 -6426 412934 -6342
rect 412314 -6662 412346 -6426
rect 412582 -6662 412666 -6426
rect 412902 -6662 412934 -6426
rect 412314 -7654 412934 -6662
rect 417434 -7066 418054 13000
rect 418834 10894 419454 13000
rect 418834 10658 418866 10894
rect 419102 10658 419186 10894
rect 419422 10658 419454 10894
rect 418834 10574 419454 10658
rect 418834 10338 418866 10574
rect 419102 10338 419186 10574
rect 419422 10338 419454 10574
rect 418834 -4186 419454 10338
rect 420234 -3226 420854 13000
rect 421634 3454 422254 13000
rect 421634 3218 421666 3454
rect 421902 3218 421986 3454
rect 422222 3218 422254 3454
rect 421634 3134 422254 3218
rect 421634 2898 421666 3134
rect 421902 2898 421986 3134
rect 422222 2898 422254 3134
rect 421634 -346 422254 2898
rect 421634 -582 421666 -346
rect 421902 -582 421986 -346
rect 422222 -582 422254 -346
rect 421634 -666 422254 -582
rect 421634 -902 421666 -666
rect 421902 -902 421986 -666
rect 422222 -902 422254 -666
rect 421634 -1894 422254 -902
rect 420234 -3462 420266 -3226
rect 420502 -3462 420586 -3226
rect 420822 -3462 420854 -3226
rect 420234 -3546 420854 -3462
rect 420234 -3782 420266 -3546
rect 420502 -3782 420586 -3546
rect 420822 -3782 420854 -3546
rect 420234 -3814 420854 -3782
rect 418834 -4422 418866 -4186
rect 419102 -4422 419186 -4186
rect 419422 -4422 419454 -4186
rect 418834 -4506 419454 -4422
rect 418834 -4742 418866 -4506
rect 419102 -4742 419186 -4506
rect 419422 -4742 419454 -4506
rect 418834 -5734 419454 -4742
rect 417434 -7302 417466 -7066
rect 417702 -7302 417786 -7066
rect 418022 -7302 418054 -7066
rect 417434 -7386 418054 -7302
rect 417434 -7622 417466 -7386
rect 417702 -7622 417786 -7386
rect 418022 -7622 418054 -7386
rect 417434 -7654 418054 -7622
rect 422554 -6106 423174 13000
rect 423954 -5146 424574 13000
rect 425354 7174 425974 13000
rect 425354 6938 425386 7174
rect 425622 6938 425706 7174
rect 425942 6938 425974 7174
rect 425354 6854 425974 6938
rect 425354 6618 425386 6854
rect 425622 6618 425706 6854
rect 425942 6618 425974 6854
rect 425354 -2266 425974 6618
rect 426754 -1306 427374 13000
rect 426754 -1542 426786 -1306
rect 427022 -1542 427106 -1306
rect 427342 -1542 427374 -1306
rect 426754 -1626 427374 -1542
rect 426754 -1862 426786 -1626
rect 427022 -1862 427106 -1626
rect 427342 -1862 427374 -1626
rect 426754 -1894 427374 -1862
rect 425354 -2502 425386 -2266
rect 425622 -2502 425706 -2266
rect 425942 -2502 425974 -2266
rect 425354 -2586 425974 -2502
rect 425354 -2822 425386 -2586
rect 425622 -2822 425706 -2586
rect 425942 -2822 425974 -2586
rect 425354 -3814 425974 -2822
rect 423954 -5382 423986 -5146
rect 424222 -5382 424306 -5146
rect 424542 -5382 424574 -5146
rect 423954 -5466 424574 -5382
rect 423954 -5702 423986 -5466
rect 424222 -5702 424306 -5466
rect 424542 -5702 424574 -5466
rect 423954 -5734 424574 -5702
rect 422554 -6342 422586 -6106
rect 422822 -6342 422906 -6106
rect 423142 -6342 423174 -6106
rect 422554 -6426 423174 -6342
rect 422554 -6662 422586 -6426
rect 422822 -6662 422906 -6426
rect 423142 -6662 423174 -6426
rect 422554 -7654 423174 -6662
rect 427674 -7066 428294 13000
rect 429074 10894 429694 13000
rect 429074 10658 429106 10894
rect 429342 10658 429426 10894
rect 429662 10658 429694 10894
rect 429074 10574 429694 10658
rect 429074 10338 429106 10574
rect 429342 10338 429426 10574
rect 429662 10338 429694 10574
rect 429074 -4186 429694 10338
rect 430474 -3226 431094 13000
rect 431874 3454 432494 13000
rect 431874 3218 431906 3454
rect 432142 3218 432226 3454
rect 432462 3218 432494 3454
rect 431874 3134 432494 3218
rect 431874 2898 431906 3134
rect 432142 2898 432226 3134
rect 432462 2898 432494 3134
rect 431874 -346 432494 2898
rect 431874 -582 431906 -346
rect 432142 -582 432226 -346
rect 432462 -582 432494 -346
rect 431874 -666 432494 -582
rect 431874 -902 431906 -666
rect 432142 -902 432226 -666
rect 432462 -902 432494 -666
rect 431874 -1894 432494 -902
rect 430474 -3462 430506 -3226
rect 430742 -3462 430826 -3226
rect 431062 -3462 431094 -3226
rect 430474 -3546 431094 -3462
rect 430474 -3782 430506 -3546
rect 430742 -3782 430826 -3546
rect 431062 -3782 431094 -3546
rect 430474 -3814 431094 -3782
rect 429074 -4422 429106 -4186
rect 429342 -4422 429426 -4186
rect 429662 -4422 429694 -4186
rect 429074 -4506 429694 -4422
rect 429074 -4742 429106 -4506
rect 429342 -4742 429426 -4506
rect 429662 -4742 429694 -4506
rect 429074 -5734 429694 -4742
rect 427674 -7302 427706 -7066
rect 427942 -7302 428026 -7066
rect 428262 -7302 428294 -7066
rect 427674 -7386 428294 -7302
rect 427674 -7622 427706 -7386
rect 427942 -7622 428026 -7386
rect 428262 -7622 428294 -7386
rect 427674 -7654 428294 -7622
rect 432794 -6106 433414 13000
rect 434194 -5146 434814 13000
rect 435594 7174 436214 13000
rect 435594 6938 435626 7174
rect 435862 6938 435946 7174
rect 436182 6938 436214 7174
rect 435594 6854 436214 6938
rect 435594 6618 435626 6854
rect 435862 6618 435946 6854
rect 436182 6618 436214 6854
rect 435594 -2266 436214 6618
rect 436994 -1306 437614 13000
rect 436994 -1542 437026 -1306
rect 437262 -1542 437346 -1306
rect 437582 -1542 437614 -1306
rect 436994 -1626 437614 -1542
rect 436994 -1862 437026 -1626
rect 437262 -1862 437346 -1626
rect 437582 -1862 437614 -1626
rect 436994 -1894 437614 -1862
rect 435594 -2502 435626 -2266
rect 435862 -2502 435946 -2266
rect 436182 -2502 436214 -2266
rect 435594 -2586 436214 -2502
rect 435594 -2822 435626 -2586
rect 435862 -2822 435946 -2586
rect 436182 -2822 436214 -2586
rect 435594 -3814 436214 -2822
rect 434194 -5382 434226 -5146
rect 434462 -5382 434546 -5146
rect 434782 -5382 434814 -5146
rect 434194 -5466 434814 -5382
rect 434194 -5702 434226 -5466
rect 434462 -5702 434546 -5466
rect 434782 -5702 434814 -5466
rect 434194 -5734 434814 -5702
rect 432794 -6342 432826 -6106
rect 433062 -6342 433146 -6106
rect 433382 -6342 433414 -6106
rect 432794 -6426 433414 -6342
rect 432794 -6662 432826 -6426
rect 433062 -6662 433146 -6426
rect 433382 -6662 433414 -6426
rect 432794 -7654 433414 -6662
rect 437914 -7066 438534 13000
rect 439314 10894 439934 13000
rect 439314 10658 439346 10894
rect 439582 10658 439666 10894
rect 439902 10658 439934 10894
rect 439314 10574 439934 10658
rect 439314 10338 439346 10574
rect 439582 10338 439666 10574
rect 439902 10338 439934 10574
rect 439314 -4186 439934 10338
rect 440714 -3226 441334 13000
rect 442114 3454 442734 13000
rect 442114 3218 442146 3454
rect 442382 3218 442466 3454
rect 442702 3218 442734 3454
rect 442114 3134 442734 3218
rect 442114 2898 442146 3134
rect 442382 2898 442466 3134
rect 442702 2898 442734 3134
rect 442114 -346 442734 2898
rect 442114 -582 442146 -346
rect 442382 -582 442466 -346
rect 442702 -582 442734 -346
rect 442114 -666 442734 -582
rect 442114 -902 442146 -666
rect 442382 -902 442466 -666
rect 442702 -902 442734 -666
rect 442114 -1894 442734 -902
rect 440714 -3462 440746 -3226
rect 440982 -3462 441066 -3226
rect 441302 -3462 441334 -3226
rect 440714 -3546 441334 -3462
rect 440714 -3782 440746 -3546
rect 440982 -3782 441066 -3546
rect 441302 -3782 441334 -3546
rect 440714 -3814 441334 -3782
rect 439314 -4422 439346 -4186
rect 439582 -4422 439666 -4186
rect 439902 -4422 439934 -4186
rect 439314 -4506 439934 -4422
rect 439314 -4742 439346 -4506
rect 439582 -4742 439666 -4506
rect 439902 -4742 439934 -4506
rect 439314 -5734 439934 -4742
rect 437914 -7302 437946 -7066
rect 438182 -7302 438266 -7066
rect 438502 -7302 438534 -7066
rect 437914 -7386 438534 -7302
rect 437914 -7622 437946 -7386
rect 438182 -7622 438266 -7386
rect 438502 -7622 438534 -7386
rect 437914 -7654 438534 -7622
rect 443034 -6106 443654 13000
rect 444434 -5146 445054 13000
rect 445834 7174 446454 13000
rect 445834 6938 445866 7174
rect 446102 6938 446186 7174
rect 446422 6938 446454 7174
rect 445834 6854 446454 6938
rect 445834 6618 445866 6854
rect 446102 6618 446186 6854
rect 446422 6618 446454 6854
rect 445834 -2266 446454 6618
rect 447234 -1306 447854 13000
rect 447234 -1542 447266 -1306
rect 447502 -1542 447586 -1306
rect 447822 -1542 447854 -1306
rect 447234 -1626 447854 -1542
rect 447234 -1862 447266 -1626
rect 447502 -1862 447586 -1626
rect 447822 -1862 447854 -1626
rect 447234 -1894 447854 -1862
rect 445834 -2502 445866 -2266
rect 446102 -2502 446186 -2266
rect 446422 -2502 446454 -2266
rect 445834 -2586 446454 -2502
rect 445834 -2822 445866 -2586
rect 446102 -2822 446186 -2586
rect 446422 -2822 446454 -2586
rect 445834 -3814 446454 -2822
rect 444434 -5382 444466 -5146
rect 444702 -5382 444786 -5146
rect 445022 -5382 445054 -5146
rect 444434 -5466 445054 -5382
rect 444434 -5702 444466 -5466
rect 444702 -5702 444786 -5466
rect 445022 -5702 445054 -5466
rect 444434 -5734 445054 -5702
rect 443034 -6342 443066 -6106
rect 443302 -6342 443386 -6106
rect 443622 -6342 443654 -6106
rect 443034 -6426 443654 -6342
rect 443034 -6662 443066 -6426
rect 443302 -6662 443386 -6426
rect 443622 -6662 443654 -6426
rect 443034 -7654 443654 -6662
rect 448154 -7066 448774 13000
rect 449554 10894 450174 13000
rect 449554 10658 449586 10894
rect 449822 10658 449906 10894
rect 450142 10658 450174 10894
rect 449554 10574 450174 10658
rect 449554 10338 449586 10574
rect 449822 10338 449906 10574
rect 450142 10338 450174 10574
rect 449554 -4186 450174 10338
rect 450954 -3226 451574 13000
rect 452354 3454 452974 13000
rect 452354 3218 452386 3454
rect 452622 3218 452706 3454
rect 452942 3218 452974 3454
rect 452354 3134 452974 3218
rect 452354 2898 452386 3134
rect 452622 2898 452706 3134
rect 452942 2898 452974 3134
rect 452354 -346 452974 2898
rect 452354 -582 452386 -346
rect 452622 -582 452706 -346
rect 452942 -582 452974 -346
rect 452354 -666 452974 -582
rect 452354 -902 452386 -666
rect 452622 -902 452706 -666
rect 452942 -902 452974 -666
rect 452354 -1894 452974 -902
rect 450954 -3462 450986 -3226
rect 451222 -3462 451306 -3226
rect 451542 -3462 451574 -3226
rect 450954 -3546 451574 -3462
rect 450954 -3782 450986 -3546
rect 451222 -3782 451306 -3546
rect 451542 -3782 451574 -3546
rect 450954 -3814 451574 -3782
rect 449554 -4422 449586 -4186
rect 449822 -4422 449906 -4186
rect 450142 -4422 450174 -4186
rect 449554 -4506 450174 -4422
rect 449554 -4742 449586 -4506
rect 449822 -4742 449906 -4506
rect 450142 -4742 450174 -4506
rect 449554 -5734 450174 -4742
rect 448154 -7302 448186 -7066
rect 448422 -7302 448506 -7066
rect 448742 -7302 448774 -7066
rect 448154 -7386 448774 -7302
rect 448154 -7622 448186 -7386
rect 448422 -7622 448506 -7386
rect 448742 -7622 448774 -7386
rect 448154 -7654 448774 -7622
rect 453274 -6106 453894 13000
rect 454674 -5146 455294 13000
rect 456074 7174 456694 13000
rect 456074 6938 456106 7174
rect 456342 6938 456426 7174
rect 456662 6938 456694 7174
rect 456074 6854 456694 6938
rect 456074 6618 456106 6854
rect 456342 6618 456426 6854
rect 456662 6618 456694 6854
rect 456074 -2266 456694 6618
rect 457474 -1306 458094 13000
rect 457474 -1542 457506 -1306
rect 457742 -1542 457826 -1306
rect 458062 -1542 458094 -1306
rect 457474 -1626 458094 -1542
rect 457474 -1862 457506 -1626
rect 457742 -1862 457826 -1626
rect 458062 -1862 458094 -1626
rect 457474 -1894 458094 -1862
rect 456074 -2502 456106 -2266
rect 456342 -2502 456426 -2266
rect 456662 -2502 456694 -2266
rect 456074 -2586 456694 -2502
rect 456074 -2822 456106 -2586
rect 456342 -2822 456426 -2586
rect 456662 -2822 456694 -2586
rect 456074 -3814 456694 -2822
rect 454674 -5382 454706 -5146
rect 454942 -5382 455026 -5146
rect 455262 -5382 455294 -5146
rect 454674 -5466 455294 -5382
rect 454674 -5702 454706 -5466
rect 454942 -5702 455026 -5466
rect 455262 -5702 455294 -5466
rect 454674 -5734 455294 -5702
rect 453274 -6342 453306 -6106
rect 453542 -6342 453626 -6106
rect 453862 -6342 453894 -6106
rect 453274 -6426 453894 -6342
rect 453274 -6662 453306 -6426
rect 453542 -6662 453626 -6426
rect 453862 -6662 453894 -6426
rect 453274 -7654 453894 -6662
rect 458394 -7066 459014 13000
rect 459794 10894 460414 13000
rect 459794 10658 459826 10894
rect 460062 10658 460146 10894
rect 460382 10658 460414 10894
rect 459794 10574 460414 10658
rect 459794 10338 459826 10574
rect 460062 10338 460146 10574
rect 460382 10338 460414 10574
rect 459794 -4186 460414 10338
rect 461194 -3226 461814 13000
rect 462594 3454 463214 13000
rect 462594 3218 462626 3454
rect 462862 3218 462946 3454
rect 463182 3218 463214 3454
rect 462594 3134 463214 3218
rect 462594 2898 462626 3134
rect 462862 2898 462946 3134
rect 463182 2898 463214 3134
rect 462594 -346 463214 2898
rect 462594 -582 462626 -346
rect 462862 -582 462946 -346
rect 463182 -582 463214 -346
rect 462594 -666 463214 -582
rect 462594 -902 462626 -666
rect 462862 -902 462946 -666
rect 463182 -902 463214 -666
rect 462594 -1894 463214 -902
rect 461194 -3462 461226 -3226
rect 461462 -3462 461546 -3226
rect 461782 -3462 461814 -3226
rect 461194 -3546 461814 -3462
rect 461194 -3782 461226 -3546
rect 461462 -3782 461546 -3546
rect 461782 -3782 461814 -3546
rect 461194 -3814 461814 -3782
rect 459794 -4422 459826 -4186
rect 460062 -4422 460146 -4186
rect 460382 -4422 460414 -4186
rect 459794 -4506 460414 -4422
rect 459794 -4742 459826 -4506
rect 460062 -4742 460146 -4506
rect 460382 -4742 460414 -4506
rect 459794 -5734 460414 -4742
rect 458394 -7302 458426 -7066
rect 458662 -7302 458746 -7066
rect 458982 -7302 459014 -7066
rect 458394 -7386 459014 -7302
rect 458394 -7622 458426 -7386
rect 458662 -7622 458746 -7386
rect 458982 -7622 459014 -7386
rect 458394 -7654 459014 -7622
rect 463514 -6106 464134 13000
rect 464914 -5146 465534 13000
rect 466314 7174 466934 13000
rect 466314 6938 466346 7174
rect 466582 6938 466666 7174
rect 466902 6938 466934 7174
rect 466314 6854 466934 6938
rect 466314 6618 466346 6854
rect 466582 6618 466666 6854
rect 466902 6618 466934 6854
rect 466314 -2266 466934 6618
rect 467714 -1306 468334 13000
rect 467714 -1542 467746 -1306
rect 467982 -1542 468066 -1306
rect 468302 -1542 468334 -1306
rect 467714 -1626 468334 -1542
rect 467714 -1862 467746 -1626
rect 467982 -1862 468066 -1626
rect 468302 -1862 468334 -1626
rect 467714 -1894 468334 -1862
rect 466314 -2502 466346 -2266
rect 466582 -2502 466666 -2266
rect 466902 -2502 466934 -2266
rect 466314 -2586 466934 -2502
rect 466314 -2822 466346 -2586
rect 466582 -2822 466666 -2586
rect 466902 -2822 466934 -2586
rect 466314 -3814 466934 -2822
rect 464914 -5382 464946 -5146
rect 465182 -5382 465266 -5146
rect 465502 -5382 465534 -5146
rect 464914 -5466 465534 -5382
rect 464914 -5702 464946 -5466
rect 465182 -5702 465266 -5466
rect 465502 -5702 465534 -5466
rect 464914 -5734 465534 -5702
rect 463514 -6342 463546 -6106
rect 463782 -6342 463866 -6106
rect 464102 -6342 464134 -6106
rect 463514 -6426 464134 -6342
rect 463514 -6662 463546 -6426
rect 463782 -6662 463866 -6426
rect 464102 -6662 464134 -6426
rect 463514 -7654 464134 -6662
rect 468634 -7066 469254 13000
rect 470034 10894 470654 13000
rect 470034 10658 470066 10894
rect 470302 10658 470386 10894
rect 470622 10658 470654 10894
rect 470034 10574 470654 10658
rect 470034 10338 470066 10574
rect 470302 10338 470386 10574
rect 470622 10338 470654 10574
rect 470034 -4186 470654 10338
rect 471434 -3226 472054 13000
rect 472834 3454 473454 13000
rect 472834 3218 472866 3454
rect 473102 3218 473186 3454
rect 473422 3218 473454 3454
rect 472834 3134 473454 3218
rect 472834 2898 472866 3134
rect 473102 2898 473186 3134
rect 473422 2898 473454 3134
rect 472834 -346 473454 2898
rect 472834 -582 472866 -346
rect 473102 -582 473186 -346
rect 473422 -582 473454 -346
rect 472834 -666 473454 -582
rect 472834 -902 472866 -666
rect 473102 -902 473186 -666
rect 473422 -902 473454 -666
rect 472834 -1894 473454 -902
rect 471434 -3462 471466 -3226
rect 471702 -3462 471786 -3226
rect 472022 -3462 472054 -3226
rect 471434 -3546 472054 -3462
rect 471434 -3782 471466 -3546
rect 471702 -3782 471786 -3546
rect 472022 -3782 472054 -3546
rect 471434 -3814 472054 -3782
rect 470034 -4422 470066 -4186
rect 470302 -4422 470386 -4186
rect 470622 -4422 470654 -4186
rect 470034 -4506 470654 -4422
rect 470034 -4742 470066 -4506
rect 470302 -4742 470386 -4506
rect 470622 -4742 470654 -4506
rect 470034 -5734 470654 -4742
rect 468634 -7302 468666 -7066
rect 468902 -7302 468986 -7066
rect 469222 -7302 469254 -7066
rect 468634 -7386 469254 -7302
rect 468634 -7622 468666 -7386
rect 468902 -7622 468986 -7386
rect 469222 -7622 469254 -7386
rect 468634 -7654 469254 -7622
rect 473754 -6106 474374 13000
rect 475154 -5146 475774 13000
rect 476554 7174 477174 13000
rect 476554 6938 476586 7174
rect 476822 6938 476906 7174
rect 477142 6938 477174 7174
rect 476554 6854 477174 6938
rect 476554 6618 476586 6854
rect 476822 6618 476906 6854
rect 477142 6618 477174 6854
rect 476554 -2266 477174 6618
rect 477954 -1306 478574 13000
rect 477954 -1542 477986 -1306
rect 478222 -1542 478306 -1306
rect 478542 -1542 478574 -1306
rect 477954 -1626 478574 -1542
rect 477954 -1862 477986 -1626
rect 478222 -1862 478306 -1626
rect 478542 -1862 478574 -1626
rect 477954 -1894 478574 -1862
rect 476554 -2502 476586 -2266
rect 476822 -2502 476906 -2266
rect 477142 -2502 477174 -2266
rect 476554 -2586 477174 -2502
rect 476554 -2822 476586 -2586
rect 476822 -2822 476906 -2586
rect 477142 -2822 477174 -2586
rect 476554 -3814 477174 -2822
rect 475154 -5382 475186 -5146
rect 475422 -5382 475506 -5146
rect 475742 -5382 475774 -5146
rect 475154 -5466 475774 -5382
rect 475154 -5702 475186 -5466
rect 475422 -5702 475506 -5466
rect 475742 -5702 475774 -5466
rect 475154 -5734 475774 -5702
rect 473754 -6342 473786 -6106
rect 474022 -6342 474106 -6106
rect 474342 -6342 474374 -6106
rect 473754 -6426 474374 -6342
rect 473754 -6662 473786 -6426
rect 474022 -6662 474106 -6426
rect 474342 -6662 474374 -6426
rect 473754 -7654 474374 -6662
rect 478874 -7066 479494 13000
rect 480274 10894 480894 13000
rect 480274 10658 480306 10894
rect 480542 10658 480626 10894
rect 480862 10658 480894 10894
rect 480274 10574 480894 10658
rect 480274 10338 480306 10574
rect 480542 10338 480626 10574
rect 480862 10338 480894 10574
rect 480274 -4186 480894 10338
rect 481674 -3226 482294 13000
rect 483074 3454 483694 13000
rect 483074 3218 483106 3454
rect 483342 3218 483426 3454
rect 483662 3218 483694 3454
rect 483074 3134 483694 3218
rect 483074 2898 483106 3134
rect 483342 2898 483426 3134
rect 483662 2898 483694 3134
rect 483074 -346 483694 2898
rect 483074 -582 483106 -346
rect 483342 -582 483426 -346
rect 483662 -582 483694 -346
rect 483074 -666 483694 -582
rect 483074 -902 483106 -666
rect 483342 -902 483426 -666
rect 483662 -902 483694 -666
rect 483074 -1894 483694 -902
rect 481674 -3462 481706 -3226
rect 481942 -3462 482026 -3226
rect 482262 -3462 482294 -3226
rect 481674 -3546 482294 -3462
rect 481674 -3782 481706 -3546
rect 481942 -3782 482026 -3546
rect 482262 -3782 482294 -3546
rect 481674 -3814 482294 -3782
rect 480274 -4422 480306 -4186
rect 480542 -4422 480626 -4186
rect 480862 -4422 480894 -4186
rect 480274 -4506 480894 -4422
rect 480274 -4742 480306 -4506
rect 480542 -4742 480626 -4506
rect 480862 -4742 480894 -4506
rect 480274 -5734 480894 -4742
rect 478874 -7302 478906 -7066
rect 479142 -7302 479226 -7066
rect 479462 -7302 479494 -7066
rect 478874 -7386 479494 -7302
rect 478874 -7622 478906 -7386
rect 479142 -7622 479226 -7386
rect 479462 -7622 479494 -7386
rect 478874 -7654 479494 -7622
rect 483994 -6106 484614 13000
rect 485394 -5146 486014 13000
rect 486794 7174 487414 13000
rect 486794 6938 486826 7174
rect 487062 6938 487146 7174
rect 487382 6938 487414 7174
rect 486794 6854 487414 6938
rect 486794 6618 486826 6854
rect 487062 6618 487146 6854
rect 487382 6618 487414 6854
rect 486794 -2266 487414 6618
rect 488194 -1306 488814 13000
rect 488194 -1542 488226 -1306
rect 488462 -1542 488546 -1306
rect 488782 -1542 488814 -1306
rect 488194 -1626 488814 -1542
rect 488194 -1862 488226 -1626
rect 488462 -1862 488546 -1626
rect 488782 -1862 488814 -1626
rect 488194 -1894 488814 -1862
rect 486794 -2502 486826 -2266
rect 487062 -2502 487146 -2266
rect 487382 -2502 487414 -2266
rect 486794 -2586 487414 -2502
rect 486794 -2822 486826 -2586
rect 487062 -2822 487146 -2586
rect 487382 -2822 487414 -2586
rect 486794 -3814 487414 -2822
rect 485394 -5382 485426 -5146
rect 485662 -5382 485746 -5146
rect 485982 -5382 486014 -5146
rect 485394 -5466 486014 -5382
rect 485394 -5702 485426 -5466
rect 485662 -5702 485746 -5466
rect 485982 -5702 486014 -5466
rect 485394 -5734 486014 -5702
rect 483994 -6342 484026 -6106
rect 484262 -6342 484346 -6106
rect 484582 -6342 484614 -6106
rect 483994 -6426 484614 -6342
rect 483994 -6662 484026 -6426
rect 484262 -6662 484346 -6426
rect 484582 -6662 484614 -6426
rect 483994 -7654 484614 -6662
rect 489114 -7066 489734 13000
rect 490514 10894 491134 13000
rect 490514 10658 490546 10894
rect 490782 10658 490866 10894
rect 491102 10658 491134 10894
rect 490514 10574 491134 10658
rect 490514 10338 490546 10574
rect 490782 10338 490866 10574
rect 491102 10338 491134 10574
rect 490514 -4186 491134 10338
rect 491914 -3226 492534 13000
rect 493314 3454 493934 13000
rect 493314 3218 493346 3454
rect 493582 3218 493666 3454
rect 493902 3218 493934 3454
rect 493314 3134 493934 3218
rect 493314 2898 493346 3134
rect 493582 2898 493666 3134
rect 493902 2898 493934 3134
rect 493314 -346 493934 2898
rect 493314 -582 493346 -346
rect 493582 -582 493666 -346
rect 493902 -582 493934 -346
rect 493314 -666 493934 -582
rect 493314 -902 493346 -666
rect 493582 -902 493666 -666
rect 493902 -902 493934 -666
rect 493314 -1894 493934 -902
rect 491914 -3462 491946 -3226
rect 492182 -3462 492266 -3226
rect 492502 -3462 492534 -3226
rect 491914 -3546 492534 -3462
rect 491914 -3782 491946 -3546
rect 492182 -3782 492266 -3546
rect 492502 -3782 492534 -3546
rect 491914 -3814 492534 -3782
rect 490514 -4422 490546 -4186
rect 490782 -4422 490866 -4186
rect 491102 -4422 491134 -4186
rect 490514 -4506 491134 -4422
rect 490514 -4742 490546 -4506
rect 490782 -4742 490866 -4506
rect 491102 -4742 491134 -4506
rect 490514 -5734 491134 -4742
rect 489114 -7302 489146 -7066
rect 489382 -7302 489466 -7066
rect 489702 -7302 489734 -7066
rect 489114 -7386 489734 -7302
rect 489114 -7622 489146 -7386
rect 489382 -7622 489466 -7386
rect 489702 -7622 489734 -7386
rect 489114 -7654 489734 -7622
rect 494234 -6106 494854 13000
rect 495634 -5146 496254 13000
rect 497034 7174 497654 13000
rect 497034 6938 497066 7174
rect 497302 6938 497386 7174
rect 497622 6938 497654 7174
rect 497034 6854 497654 6938
rect 497034 6618 497066 6854
rect 497302 6618 497386 6854
rect 497622 6618 497654 6854
rect 497034 -2266 497654 6618
rect 498434 -1306 499054 13000
rect 498434 -1542 498466 -1306
rect 498702 -1542 498786 -1306
rect 499022 -1542 499054 -1306
rect 498434 -1626 499054 -1542
rect 498434 -1862 498466 -1626
rect 498702 -1862 498786 -1626
rect 499022 -1862 499054 -1626
rect 498434 -1894 499054 -1862
rect 497034 -2502 497066 -2266
rect 497302 -2502 497386 -2266
rect 497622 -2502 497654 -2266
rect 497034 -2586 497654 -2502
rect 497034 -2822 497066 -2586
rect 497302 -2822 497386 -2586
rect 497622 -2822 497654 -2586
rect 497034 -3814 497654 -2822
rect 495634 -5382 495666 -5146
rect 495902 -5382 495986 -5146
rect 496222 -5382 496254 -5146
rect 495634 -5466 496254 -5382
rect 495634 -5702 495666 -5466
rect 495902 -5702 495986 -5466
rect 496222 -5702 496254 -5466
rect 495634 -5734 496254 -5702
rect 494234 -6342 494266 -6106
rect 494502 -6342 494586 -6106
rect 494822 -6342 494854 -6106
rect 494234 -6426 494854 -6342
rect 494234 -6662 494266 -6426
rect 494502 -6662 494586 -6426
rect 494822 -6662 494854 -6426
rect 494234 -7654 494854 -6662
rect 499354 -7066 499974 13000
rect 500754 10894 501374 13000
rect 500754 10658 500786 10894
rect 501022 10658 501106 10894
rect 501342 10658 501374 10894
rect 500754 10574 501374 10658
rect 500754 10338 500786 10574
rect 501022 10338 501106 10574
rect 501342 10338 501374 10574
rect 500754 -4186 501374 10338
rect 502154 -3226 502774 13000
rect 503554 3454 504174 13000
rect 503554 3218 503586 3454
rect 503822 3218 503906 3454
rect 504142 3218 504174 3454
rect 503554 3134 504174 3218
rect 503554 2898 503586 3134
rect 503822 2898 503906 3134
rect 504142 2898 504174 3134
rect 503554 -346 504174 2898
rect 503554 -582 503586 -346
rect 503822 -582 503906 -346
rect 504142 -582 504174 -346
rect 503554 -666 504174 -582
rect 503554 -902 503586 -666
rect 503822 -902 503906 -666
rect 504142 -902 504174 -666
rect 503554 -1894 504174 -902
rect 502154 -3462 502186 -3226
rect 502422 -3462 502506 -3226
rect 502742 -3462 502774 -3226
rect 502154 -3546 502774 -3462
rect 502154 -3782 502186 -3546
rect 502422 -3782 502506 -3546
rect 502742 -3782 502774 -3546
rect 502154 -3814 502774 -3782
rect 500754 -4422 500786 -4186
rect 501022 -4422 501106 -4186
rect 501342 -4422 501374 -4186
rect 500754 -4506 501374 -4422
rect 500754 -4742 500786 -4506
rect 501022 -4742 501106 -4506
rect 501342 -4742 501374 -4506
rect 500754 -5734 501374 -4742
rect 499354 -7302 499386 -7066
rect 499622 -7302 499706 -7066
rect 499942 -7302 499974 -7066
rect 499354 -7386 499974 -7302
rect 499354 -7622 499386 -7386
rect 499622 -7622 499706 -7386
rect 499942 -7622 499974 -7386
rect 499354 -7654 499974 -7622
rect 504474 -6106 505094 13000
rect 505874 -5146 506494 13000
rect 507274 7174 507894 13000
rect 507274 6938 507306 7174
rect 507542 6938 507626 7174
rect 507862 6938 507894 7174
rect 507274 6854 507894 6938
rect 507274 6618 507306 6854
rect 507542 6618 507626 6854
rect 507862 6618 507894 6854
rect 507274 -2266 507894 6618
rect 508674 -1306 509294 13000
rect 508674 -1542 508706 -1306
rect 508942 -1542 509026 -1306
rect 509262 -1542 509294 -1306
rect 508674 -1626 509294 -1542
rect 508674 -1862 508706 -1626
rect 508942 -1862 509026 -1626
rect 509262 -1862 509294 -1626
rect 508674 -1894 509294 -1862
rect 507274 -2502 507306 -2266
rect 507542 -2502 507626 -2266
rect 507862 -2502 507894 -2266
rect 507274 -2586 507894 -2502
rect 507274 -2822 507306 -2586
rect 507542 -2822 507626 -2586
rect 507862 -2822 507894 -2586
rect 507274 -3814 507894 -2822
rect 505874 -5382 505906 -5146
rect 506142 -5382 506226 -5146
rect 506462 -5382 506494 -5146
rect 505874 -5466 506494 -5382
rect 505874 -5702 505906 -5466
rect 506142 -5702 506226 -5466
rect 506462 -5702 506494 -5466
rect 505874 -5734 506494 -5702
rect 504474 -6342 504506 -6106
rect 504742 -6342 504826 -6106
rect 505062 -6342 505094 -6106
rect 504474 -6426 505094 -6342
rect 504474 -6662 504506 -6426
rect 504742 -6662 504826 -6426
rect 505062 -6662 505094 -6426
rect 504474 -7654 505094 -6662
rect 509594 -7066 510214 13000
rect 510994 10894 511614 13000
rect 510994 10658 511026 10894
rect 511262 10658 511346 10894
rect 511582 10658 511614 10894
rect 510994 10574 511614 10658
rect 510994 10338 511026 10574
rect 511262 10338 511346 10574
rect 511582 10338 511614 10574
rect 510994 -4186 511614 10338
rect 512394 -3226 513014 13000
rect 513794 3454 514414 13000
rect 513794 3218 513826 3454
rect 514062 3218 514146 3454
rect 514382 3218 514414 3454
rect 513794 3134 514414 3218
rect 513794 2898 513826 3134
rect 514062 2898 514146 3134
rect 514382 2898 514414 3134
rect 513794 -346 514414 2898
rect 513794 -582 513826 -346
rect 514062 -582 514146 -346
rect 514382 -582 514414 -346
rect 513794 -666 514414 -582
rect 513794 -902 513826 -666
rect 514062 -902 514146 -666
rect 514382 -902 514414 -666
rect 513794 -1894 514414 -902
rect 512394 -3462 512426 -3226
rect 512662 -3462 512746 -3226
rect 512982 -3462 513014 -3226
rect 512394 -3546 513014 -3462
rect 512394 -3782 512426 -3546
rect 512662 -3782 512746 -3546
rect 512982 -3782 513014 -3546
rect 512394 -3814 513014 -3782
rect 510994 -4422 511026 -4186
rect 511262 -4422 511346 -4186
rect 511582 -4422 511614 -4186
rect 510994 -4506 511614 -4422
rect 510994 -4742 511026 -4506
rect 511262 -4742 511346 -4506
rect 511582 -4742 511614 -4506
rect 510994 -5734 511614 -4742
rect 509594 -7302 509626 -7066
rect 509862 -7302 509946 -7066
rect 510182 -7302 510214 -7066
rect 509594 -7386 510214 -7302
rect 509594 -7622 509626 -7386
rect 509862 -7622 509946 -7386
rect 510182 -7622 510214 -7386
rect 509594 -7654 510214 -7622
rect 514714 -6106 515334 13000
rect 516114 -5146 516734 13000
rect 517514 7174 518134 13000
rect 517514 6938 517546 7174
rect 517782 6938 517866 7174
rect 518102 6938 518134 7174
rect 517514 6854 518134 6938
rect 517514 6618 517546 6854
rect 517782 6618 517866 6854
rect 518102 6618 518134 6854
rect 517514 -2266 518134 6618
rect 518914 -1306 519534 13000
rect 518914 -1542 518946 -1306
rect 519182 -1542 519266 -1306
rect 519502 -1542 519534 -1306
rect 518914 -1626 519534 -1542
rect 518914 -1862 518946 -1626
rect 519182 -1862 519266 -1626
rect 519502 -1862 519534 -1626
rect 518914 -1894 519534 -1862
rect 517514 -2502 517546 -2266
rect 517782 -2502 517866 -2266
rect 518102 -2502 518134 -2266
rect 517514 -2586 518134 -2502
rect 517514 -2822 517546 -2586
rect 517782 -2822 517866 -2586
rect 518102 -2822 518134 -2586
rect 517514 -3814 518134 -2822
rect 516114 -5382 516146 -5146
rect 516382 -5382 516466 -5146
rect 516702 -5382 516734 -5146
rect 516114 -5466 516734 -5382
rect 516114 -5702 516146 -5466
rect 516382 -5702 516466 -5466
rect 516702 -5702 516734 -5466
rect 516114 -5734 516734 -5702
rect 514714 -6342 514746 -6106
rect 514982 -6342 515066 -6106
rect 515302 -6342 515334 -6106
rect 514714 -6426 515334 -6342
rect 514714 -6662 514746 -6426
rect 514982 -6662 515066 -6426
rect 515302 -6662 515334 -6426
rect 514714 -7654 515334 -6662
rect 519834 -7066 520454 13000
rect 521234 10894 521854 13000
rect 521234 10658 521266 10894
rect 521502 10658 521586 10894
rect 521822 10658 521854 10894
rect 521234 10574 521854 10658
rect 521234 10338 521266 10574
rect 521502 10338 521586 10574
rect 521822 10338 521854 10574
rect 521234 -4186 521854 10338
rect 522634 -3226 523254 13000
rect 524034 3454 524654 13000
rect 524034 3218 524066 3454
rect 524302 3218 524386 3454
rect 524622 3218 524654 3454
rect 524034 3134 524654 3218
rect 524034 2898 524066 3134
rect 524302 2898 524386 3134
rect 524622 2898 524654 3134
rect 524034 -346 524654 2898
rect 524034 -582 524066 -346
rect 524302 -582 524386 -346
rect 524622 -582 524654 -346
rect 524034 -666 524654 -582
rect 524034 -902 524066 -666
rect 524302 -902 524386 -666
rect 524622 -902 524654 -666
rect 524034 -1894 524654 -902
rect 522634 -3462 522666 -3226
rect 522902 -3462 522986 -3226
rect 523222 -3462 523254 -3226
rect 522634 -3546 523254 -3462
rect 522634 -3782 522666 -3546
rect 522902 -3782 522986 -3546
rect 523222 -3782 523254 -3546
rect 522634 -3814 523254 -3782
rect 521234 -4422 521266 -4186
rect 521502 -4422 521586 -4186
rect 521822 -4422 521854 -4186
rect 521234 -4506 521854 -4422
rect 521234 -4742 521266 -4506
rect 521502 -4742 521586 -4506
rect 521822 -4742 521854 -4506
rect 521234 -5734 521854 -4742
rect 519834 -7302 519866 -7066
rect 520102 -7302 520186 -7066
rect 520422 -7302 520454 -7066
rect 519834 -7386 520454 -7302
rect 519834 -7622 519866 -7386
rect 520102 -7622 520186 -7386
rect 520422 -7622 520454 -7386
rect 519834 -7654 520454 -7622
rect 524954 -6106 525574 13000
rect 526354 -5146 526974 13000
rect 527754 7174 528374 13000
rect 527754 6938 527786 7174
rect 528022 6938 528106 7174
rect 528342 6938 528374 7174
rect 527754 6854 528374 6938
rect 527754 6618 527786 6854
rect 528022 6618 528106 6854
rect 528342 6618 528374 6854
rect 527754 -2266 528374 6618
rect 529154 -1306 529774 13000
rect 529154 -1542 529186 -1306
rect 529422 -1542 529506 -1306
rect 529742 -1542 529774 -1306
rect 529154 -1626 529774 -1542
rect 529154 -1862 529186 -1626
rect 529422 -1862 529506 -1626
rect 529742 -1862 529774 -1626
rect 529154 -1894 529774 -1862
rect 527754 -2502 527786 -2266
rect 528022 -2502 528106 -2266
rect 528342 -2502 528374 -2266
rect 527754 -2586 528374 -2502
rect 527754 -2822 527786 -2586
rect 528022 -2822 528106 -2586
rect 528342 -2822 528374 -2586
rect 527754 -3814 528374 -2822
rect 526354 -5382 526386 -5146
rect 526622 -5382 526706 -5146
rect 526942 -5382 526974 -5146
rect 526354 -5466 526974 -5382
rect 526354 -5702 526386 -5466
rect 526622 -5702 526706 -5466
rect 526942 -5702 526974 -5466
rect 526354 -5734 526974 -5702
rect 524954 -6342 524986 -6106
rect 525222 -6342 525306 -6106
rect 525542 -6342 525574 -6106
rect 524954 -6426 525574 -6342
rect 524954 -6662 524986 -6426
rect 525222 -6662 525306 -6426
rect 525542 -6662 525574 -6426
rect 524954 -7654 525574 -6662
rect 530074 -7066 530694 13000
rect 531474 10894 532094 13000
rect 531474 10658 531506 10894
rect 531742 10658 531826 10894
rect 532062 10658 532094 10894
rect 531474 10574 532094 10658
rect 531474 10338 531506 10574
rect 531742 10338 531826 10574
rect 532062 10338 532094 10574
rect 531474 -4186 532094 10338
rect 532874 -3226 533494 13000
rect 534274 3454 534894 13000
rect 534274 3218 534306 3454
rect 534542 3218 534626 3454
rect 534862 3218 534894 3454
rect 534274 3134 534894 3218
rect 534274 2898 534306 3134
rect 534542 2898 534626 3134
rect 534862 2898 534894 3134
rect 534274 -346 534894 2898
rect 534274 -582 534306 -346
rect 534542 -582 534626 -346
rect 534862 -582 534894 -346
rect 534274 -666 534894 -582
rect 534274 -902 534306 -666
rect 534542 -902 534626 -666
rect 534862 -902 534894 -666
rect 534274 -1894 534894 -902
rect 532874 -3462 532906 -3226
rect 533142 -3462 533226 -3226
rect 533462 -3462 533494 -3226
rect 532874 -3546 533494 -3462
rect 532874 -3782 532906 -3546
rect 533142 -3782 533226 -3546
rect 533462 -3782 533494 -3546
rect 532874 -3814 533494 -3782
rect 531474 -4422 531506 -4186
rect 531742 -4422 531826 -4186
rect 532062 -4422 532094 -4186
rect 531474 -4506 532094 -4422
rect 531474 -4742 531506 -4506
rect 531742 -4742 531826 -4506
rect 532062 -4742 532094 -4506
rect 531474 -5734 532094 -4742
rect 530074 -7302 530106 -7066
rect 530342 -7302 530426 -7066
rect 530662 -7302 530694 -7066
rect 530074 -7386 530694 -7302
rect 530074 -7622 530106 -7386
rect 530342 -7622 530426 -7386
rect 530662 -7622 530694 -7386
rect 530074 -7654 530694 -7622
rect 535194 -6106 535814 13000
rect 536594 -5146 537214 13000
rect 537994 7174 538614 13000
rect 537994 6938 538026 7174
rect 538262 6938 538346 7174
rect 538582 6938 538614 7174
rect 537994 6854 538614 6938
rect 537994 6618 538026 6854
rect 538262 6618 538346 6854
rect 538582 6618 538614 6854
rect 537994 -2266 538614 6618
rect 539394 -1306 540014 13000
rect 539394 -1542 539426 -1306
rect 539662 -1542 539746 -1306
rect 539982 -1542 540014 -1306
rect 539394 -1626 540014 -1542
rect 539394 -1862 539426 -1626
rect 539662 -1862 539746 -1626
rect 539982 -1862 540014 -1626
rect 539394 -1894 540014 -1862
rect 537994 -2502 538026 -2266
rect 538262 -2502 538346 -2266
rect 538582 -2502 538614 -2266
rect 537994 -2586 538614 -2502
rect 537994 -2822 538026 -2586
rect 538262 -2822 538346 -2586
rect 538582 -2822 538614 -2586
rect 537994 -3814 538614 -2822
rect 536594 -5382 536626 -5146
rect 536862 -5382 536946 -5146
rect 537182 -5382 537214 -5146
rect 536594 -5466 537214 -5382
rect 536594 -5702 536626 -5466
rect 536862 -5702 536946 -5466
rect 537182 -5702 537214 -5466
rect 536594 -5734 537214 -5702
rect 535194 -6342 535226 -6106
rect 535462 -6342 535546 -6106
rect 535782 -6342 535814 -6106
rect 535194 -6426 535814 -6342
rect 535194 -6662 535226 -6426
rect 535462 -6662 535546 -6426
rect 535782 -6662 535814 -6426
rect 535194 -7654 535814 -6662
rect 540314 -7066 540934 13000
rect 541714 10894 542334 46338
rect 541714 10658 541746 10894
rect 541982 10658 542066 10894
rect 542302 10658 542334 10894
rect 541714 10574 542334 10658
rect 541714 10338 541746 10574
rect 541982 10338 542066 10574
rect 542302 10338 542334 10574
rect 541714 -4186 542334 10338
rect 543114 707718 543734 707750
rect 543114 707482 543146 707718
rect 543382 707482 543466 707718
rect 543702 707482 543734 707718
rect 543114 707398 543734 707482
rect 543114 707162 543146 707398
rect 543382 707162 543466 707398
rect 543702 707162 543734 707398
rect 543114 673174 543734 707162
rect 543114 672938 543146 673174
rect 543382 672938 543466 673174
rect 543702 672938 543734 673174
rect 543114 672854 543734 672938
rect 543114 672618 543146 672854
rect 543382 672618 543466 672854
rect 543702 672618 543734 672854
rect 543114 637174 543734 672618
rect 543114 636938 543146 637174
rect 543382 636938 543466 637174
rect 543702 636938 543734 637174
rect 543114 636854 543734 636938
rect 543114 636618 543146 636854
rect 543382 636618 543466 636854
rect 543702 636618 543734 636854
rect 543114 601174 543734 636618
rect 543114 600938 543146 601174
rect 543382 600938 543466 601174
rect 543702 600938 543734 601174
rect 543114 600854 543734 600938
rect 543114 600618 543146 600854
rect 543382 600618 543466 600854
rect 543702 600618 543734 600854
rect 543114 565174 543734 600618
rect 543114 564938 543146 565174
rect 543382 564938 543466 565174
rect 543702 564938 543734 565174
rect 543114 564854 543734 564938
rect 543114 564618 543146 564854
rect 543382 564618 543466 564854
rect 543702 564618 543734 564854
rect 543114 529174 543734 564618
rect 543114 528938 543146 529174
rect 543382 528938 543466 529174
rect 543702 528938 543734 529174
rect 543114 528854 543734 528938
rect 543114 528618 543146 528854
rect 543382 528618 543466 528854
rect 543702 528618 543734 528854
rect 543114 493174 543734 528618
rect 543114 492938 543146 493174
rect 543382 492938 543466 493174
rect 543702 492938 543734 493174
rect 543114 492854 543734 492938
rect 543114 492618 543146 492854
rect 543382 492618 543466 492854
rect 543702 492618 543734 492854
rect 543114 457174 543734 492618
rect 543114 456938 543146 457174
rect 543382 456938 543466 457174
rect 543702 456938 543734 457174
rect 543114 456854 543734 456938
rect 543114 456618 543146 456854
rect 543382 456618 543466 456854
rect 543702 456618 543734 456854
rect 543114 421174 543734 456618
rect 543114 420938 543146 421174
rect 543382 420938 543466 421174
rect 543702 420938 543734 421174
rect 543114 420854 543734 420938
rect 543114 420618 543146 420854
rect 543382 420618 543466 420854
rect 543702 420618 543734 420854
rect 543114 385174 543734 420618
rect 543114 384938 543146 385174
rect 543382 384938 543466 385174
rect 543702 384938 543734 385174
rect 543114 384854 543734 384938
rect 543114 384618 543146 384854
rect 543382 384618 543466 384854
rect 543702 384618 543734 384854
rect 543114 349174 543734 384618
rect 543114 348938 543146 349174
rect 543382 348938 543466 349174
rect 543702 348938 543734 349174
rect 543114 348854 543734 348938
rect 543114 348618 543146 348854
rect 543382 348618 543466 348854
rect 543702 348618 543734 348854
rect 543114 313174 543734 348618
rect 543114 312938 543146 313174
rect 543382 312938 543466 313174
rect 543702 312938 543734 313174
rect 543114 312854 543734 312938
rect 543114 312618 543146 312854
rect 543382 312618 543466 312854
rect 543702 312618 543734 312854
rect 543114 277174 543734 312618
rect 543114 276938 543146 277174
rect 543382 276938 543466 277174
rect 543702 276938 543734 277174
rect 543114 276854 543734 276938
rect 543114 276618 543146 276854
rect 543382 276618 543466 276854
rect 543702 276618 543734 276854
rect 543114 241174 543734 276618
rect 543114 240938 543146 241174
rect 543382 240938 543466 241174
rect 543702 240938 543734 241174
rect 543114 240854 543734 240938
rect 543114 240618 543146 240854
rect 543382 240618 543466 240854
rect 543702 240618 543734 240854
rect 543114 205174 543734 240618
rect 543114 204938 543146 205174
rect 543382 204938 543466 205174
rect 543702 204938 543734 205174
rect 543114 204854 543734 204938
rect 543114 204618 543146 204854
rect 543382 204618 543466 204854
rect 543702 204618 543734 204854
rect 543114 169174 543734 204618
rect 543114 168938 543146 169174
rect 543382 168938 543466 169174
rect 543702 168938 543734 169174
rect 543114 168854 543734 168938
rect 543114 168618 543146 168854
rect 543382 168618 543466 168854
rect 543702 168618 543734 168854
rect 543114 133174 543734 168618
rect 543114 132938 543146 133174
rect 543382 132938 543466 133174
rect 543702 132938 543734 133174
rect 543114 132854 543734 132938
rect 543114 132618 543146 132854
rect 543382 132618 543466 132854
rect 543702 132618 543734 132854
rect 543114 97174 543734 132618
rect 543114 96938 543146 97174
rect 543382 96938 543466 97174
rect 543702 96938 543734 97174
rect 543114 96854 543734 96938
rect 543114 96618 543146 96854
rect 543382 96618 543466 96854
rect 543702 96618 543734 96854
rect 543114 61174 543734 96618
rect 543114 60938 543146 61174
rect 543382 60938 543466 61174
rect 543702 60938 543734 61174
rect 543114 60854 543734 60938
rect 543114 60618 543146 60854
rect 543382 60618 543466 60854
rect 543702 60618 543734 60854
rect 543114 25174 543734 60618
rect 543114 24938 543146 25174
rect 543382 24938 543466 25174
rect 543702 24938 543734 25174
rect 543114 24854 543734 24938
rect 543114 24618 543146 24854
rect 543382 24618 543466 24854
rect 543702 24618 543734 24854
rect 543114 -3226 543734 24618
rect 544514 704838 545134 705830
rect 544514 704602 544546 704838
rect 544782 704602 544866 704838
rect 545102 704602 545134 704838
rect 544514 704518 545134 704602
rect 544514 704282 544546 704518
rect 544782 704282 544866 704518
rect 545102 704282 545134 704518
rect 544514 687454 545134 704282
rect 544514 687218 544546 687454
rect 544782 687218 544866 687454
rect 545102 687218 545134 687454
rect 544514 687134 545134 687218
rect 544514 686898 544546 687134
rect 544782 686898 544866 687134
rect 545102 686898 545134 687134
rect 544514 651454 545134 686898
rect 544514 651218 544546 651454
rect 544782 651218 544866 651454
rect 545102 651218 545134 651454
rect 544514 651134 545134 651218
rect 544514 650898 544546 651134
rect 544782 650898 544866 651134
rect 545102 650898 545134 651134
rect 544514 615454 545134 650898
rect 544514 615218 544546 615454
rect 544782 615218 544866 615454
rect 545102 615218 545134 615454
rect 544514 615134 545134 615218
rect 544514 614898 544546 615134
rect 544782 614898 544866 615134
rect 545102 614898 545134 615134
rect 544514 579454 545134 614898
rect 544514 579218 544546 579454
rect 544782 579218 544866 579454
rect 545102 579218 545134 579454
rect 544514 579134 545134 579218
rect 544514 578898 544546 579134
rect 544782 578898 544866 579134
rect 545102 578898 545134 579134
rect 544514 543454 545134 578898
rect 544514 543218 544546 543454
rect 544782 543218 544866 543454
rect 545102 543218 545134 543454
rect 544514 543134 545134 543218
rect 544514 542898 544546 543134
rect 544782 542898 544866 543134
rect 545102 542898 545134 543134
rect 544514 507454 545134 542898
rect 544514 507218 544546 507454
rect 544782 507218 544866 507454
rect 545102 507218 545134 507454
rect 544514 507134 545134 507218
rect 544514 506898 544546 507134
rect 544782 506898 544866 507134
rect 545102 506898 545134 507134
rect 544514 471454 545134 506898
rect 544514 471218 544546 471454
rect 544782 471218 544866 471454
rect 545102 471218 545134 471454
rect 544514 471134 545134 471218
rect 544514 470898 544546 471134
rect 544782 470898 544866 471134
rect 545102 470898 545134 471134
rect 544514 435454 545134 470898
rect 544514 435218 544546 435454
rect 544782 435218 544866 435454
rect 545102 435218 545134 435454
rect 544514 435134 545134 435218
rect 544514 434898 544546 435134
rect 544782 434898 544866 435134
rect 545102 434898 545134 435134
rect 544514 399454 545134 434898
rect 544514 399218 544546 399454
rect 544782 399218 544866 399454
rect 545102 399218 545134 399454
rect 544514 399134 545134 399218
rect 544514 398898 544546 399134
rect 544782 398898 544866 399134
rect 545102 398898 545134 399134
rect 544514 363454 545134 398898
rect 544514 363218 544546 363454
rect 544782 363218 544866 363454
rect 545102 363218 545134 363454
rect 544514 363134 545134 363218
rect 544514 362898 544546 363134
rect 544782 362898 544866 363134
rect 545102 362898 545134 363134
rect 544514 327454 545134 362898
rect 544514 327218 544546 327454
rect 544782 327218 544866 327454
rect 545102 327218 545134 327454
rect 544514 327134 545134 327218
rect 544514 326898 544546 327134
rect 544782 326898 544866 327134
rect 545102 326898 545134 327134
rect 544514 291454 545134 326898
rect 544514 291218 544546 291454
rect 544782 291218 544866 291454
rect 545102 291218 545134 291454
rect 544514 291134 545134 291218
rect 544514 290898 544546 291134
rect 544782 290898 544866 291134
rect 545102 290898 545134 291134
rect 544514 255454 545134 290898
rect 544514 255218 544546 255454
rect 544782 255218 544866 255454
rect 545102 255218 545134 255454
rect 544514 255134 545134 255218
rect 544514 254898 544546 255134
rect 544782 254898 544866 255134
rect 545102 254898 545134 255134
rect 544514 219454 545134 254898
rect 544514 219218 544546 219454
rect 544782 219218 544866 219454
rect 545102 219218 545134 219454
rect 544514 219134 545134 219218
rect 544514 218898 544546 219134
rect 544782 218898 544866 219134
rect 545102 218898 545134 219134
rect 544514 183454 545134 218898
rect 544514 183218 544546 183454
rect 544782 183218 544866 183454
rect 545102 183218 545134 183454
rect 544514 183134 545134 183218
rect 544514 182898 544546 183134
rect 544782 182898 544866 183134
rect 545102 182898 545134 183134
rect 544514 147454 545134 182898
rect 544514 147218 544546 147454
rect 544782 147218 544866 147454
rect 545102 147218 545134 147454
rect 544514 147134 545134 147218
rect 544514 146898 544546 147134
rect 544782 146898 544866 147134
rect 545102 146898 545134 147134
rect 544514 111454 545134 146898
rect 544514 111218 544546 111454
rect 544782 111218 544866 111454
rect 545102 111218 545134 111454
rect 544514 111134 545134 111218
rect 544514 110898 544546 111134
rect 544782 110898 544866 111134
rect 545102 110898 545134 111134
rect 544514 75454 545134 110898
rect 544514 75218 544546 75454
rect 544782 75218 544866 75454
rect 545102 75218 545134 75454
rect 544514 75134 545134 75218
rect 544514 74898 544546 75134
rect 544782 74898 544866 75134
rect 545102 74898 545134 75134
rect 544514 39454 545134 74898
rect 544514 39218 544546 39454
rect 544782 39218 544866 39454
rect 545102 39218 545134 39454
rect 544514 39134 545134 39218
rect 544514 38898 544546 39134
rect 544782 38898 544866 39134
rect 545102 38898 545134 39134
rect 544514 3454 545134 38898
rect 544514 3218 544546 3454
rect 544782 3218 544866 3454
rect 545102 3218 545134 3454
rect 544514 3134 545134 3218
rect 544514 2898 544546 3134
rect 544782 2898 544866 3134
rect 545102 2898 545134 3134
rect 544514 -346 545134 2898
rect 544514 -582 544546 -346
rect 544782 -582 544866 -346
rect 545102 -582 545134 -346
rect 544514 -666 545134 -582
rect 544514 -902 544546 -666
rect 544782 -902 544866 -666
rect 545102 -902 545134 -666
rect 544514 -1894 545134 -902
rect 545434 698614 546054 710042
rect 550554 711558 551174 711590
rect 550554 711322 550586 711558
rect 550822 711322 550906 711558
rect 551142 711322 551174 711558
rect 550554 711238 551174 711322
rect 550554 711002 550586 711238
rect 550822 711002 550906 711238
rect 551142 711002 551174 711238
rect 545434 698378 545466 698614
rect 545702 698378 545786 698614
rect 546022 698378 546054 698614
rect 545434 698294 546054 698378
rect 545434 698058 545466 698294
rect 545702 698058 545786 698294
rect 546022 698058 546054 698294
rect 545434 662614 546054 698058
rect 545434 662378 545466 662614
rect 545702 662378 545786 662614
rect 546022 662378 546054 662614
rect 545434 662294 546054 662378
rect 545434 662058 545466 662294
rect 545702 662058 545786 662294
rect 546022 662058 546054 662294
rect 545434 626614 546054 662058
rect 545434 626378 545466 626614
rect 545702 626378 545786 626614
rect 546022 626378 546054 626614
rect 545434 626294 546054 626378
rect 545434 626058 545466 626294
rect 545702 626058 545786 626294
rect 546022 626058 546054 626294
rect 545434 590614 546054 626058
rect 545434 590378 545466 590614
rect 545702 590378 545786 590614
rect 546022 590378 546054 590614
rect 545434 590294 546054 590378
rect 545434 590058 545466 590294
rect 545702 590058 545786 590294
rect 546022 590058 546054 590294
rect 545434 554614 546054 590058
rect 545434 554378 545466 554614
rect 545702 554378 545786 554614
rect 546022 554378 546054 554614
rect 545434 554294 546054 554378
rect 545434 554058 545466 554294
rect 545702 554058 545786 554294
rect 546022 554058 546054 554294
rect 545434 518614 546054 554058
rect 545434 518378 545466 518614
rect 545702 518378 545786 518614
rect 546022 518378 546054 518614
rect 545434 518294 546054 518378
rect 545434 518058 545466 518294
rect 545702 518058 545786 518294
rect 546022 518058 546054 518294
rect 545434 482614 546054 518058
rect 545434 482378 545466 482614
rect 545702 482378 545786 482614
rect 546022 482378 546054 482614
rect 545434 482294 546054 482378
rect 545434 482058 545466 482294
rect 545702 482058 545786 482294
rect 546022 482058 546054 482294
rect 545434 446614 546054 482058
rect 545434 446378 545466 446614
rect 545702 446378 545786 446614
rect 546022 446378 546054 446614
rect 545434 446294 546054 446378
rect 545434 446058 545466 446294
rect 545702 446058 545786 446294
rect 546022 446058 546054 446294
rect 545434 410614 546054 446058
rect 545434 410378 545466 410614
rect 545702 410378 545786 410614
rect 546022 410378 546054 410614
rect 545434 410294 546054 410378
rect 545434 410058 545466 410294
rect 545702 410058 545786 410294
rect 546022 410058 546054 410294
rect 545434 374614 546054 410058
rect 545434 374378 545466 374614
rect 545702 374378 545786 374614
rect 546022 374378 546054 374614
rect 545434 374294 546054 374378
rect 545434 374058 545466 374294
rect 545702 374058 545786 374294
rect 546022 374058 546054 374294
rect 545434 338614 546054 374058
rect 545434 338378 545466 338614
rect 545702 338378 545786 338614
rect 546022 338378 546054 338614
rect 545434 338294 546054 338378
rect 545434 338058 545466 338294
rect 545702 338058 545786 338294
rect 546022 338058 546054 338294
rect 545434 302614 546054 338058
rect 545434 302378 545466 302614
rect 545702 302378 545786 302614
rect 546022 302378 546054 302614
rect 545434 302294 546054 302378
rect 545434 302058 545466 302294
rect 545702 302058 545786 302294
rect 546022 302058 546054 302294
rect 545434 266614 546054 302058
rect 545434 266378 545466 266614
rect 545702 266378 545786 266614
rect 546022 266378 546054 266614
rect 545434 266294 546054 266378
rect 545434 266058 545466 266294
rect 545702 266058 545786 266294
rect 546022 266058 546054 266294
rect 545434 230614 546054 266058
rect 545434 230378 545466 230614
rect 545702 230378 545786 230614
rect 546022 230378 546054 230614
rect 545434 230294 546054 230378
rect 545434 230058 545466 230294
rect 545702 230058 545786 230294
rect 546022 230058 546054 230294
rect 545434 194614 546054 230058
rect 545434 194378 545466 194614
rect 545702 194378 545786 194614
rect 546022 194378 546054 194614
rect 545434 194294 546054 194378
rect 545434 194058 545466 194294
rect 545702 194058 545786 194294
rect 546022 194058 546054 194294
rect 545434 158614 546054 194058
rect 545434 158378 545466 158614
rect 545702 158378 545786 158614
rect 546022 158378 546054 158614
rect 545434 158294 546054 158378
rect 545434 158058 545466 158294
rect 545702 158058 545786 158294
rect 546022 158058 546054 158294
rect 545434 122614 546054 158058
rect 545434 122378 545466 122614
rect 545702 122378 545786 122614
rect 546022 122378 546054 122614
rect 545434 122294 546054 122378
rect 545434 122058 545466 122294
rect 545702 122058 545786 122294
rect 546022 122058 546054 122294
rect 545434 86614 546054 122058
rect 545434 86378 545466 86614
rect 545702 86378 545786 86614
rect 546022 86378 546054 86614
rect 545434 86294 546054 86378
rect 545434 86058 545466 86294
rect 545702 86058 545786 86294
rect 546022 86058 546054 86294
rect 545434 50614 546054 86058
rect 545434 50378 545466 50614
rect 545702 50378 545786 50614
rect 546022 50378 546054 50614
rect 545434 50294 546054 50378
rect 545434 50058 545466 50294
rect 545702 50058 545786 50294
rect 546022 50058 546054 50294
rect 545434 14614 546054 50058
rect 545434 14378 545466 14614
rect 545702 14378 545786 14614
rect 546022 14378 546054 14614
rect 545434 14294 546054 14378
rect 545434 14058 545466 14294
rect 545702 14058 545786 14294
rect 546022 14058 546054 14294
rect 543114 -3462 543146 -3226
rect 543382 -3462 543466 -3226
rect 543702 -3462 543734 -3226
rect 543114 -3546 543734 -3462
rect 543114 -3782 543146 -3546
rect 543382 -3782 543466 -3546
rect 543702 -3782 543734 -3546
rect 543114 -3814 543734 -3782
rect 541714 -4422 541746 -4186
rect 541982 -4422 542066 -4186
rect 542302 -4422 542334 -4186
rect 541714 -4506 542334 -4422
rect 541714 -4742 541746 -4506
rect 541982 -4742 542066 -4506
rect 542302 -4742 542334 -4506
rect 541714 -5734 542334 -4742
rect 540314 -7302 540346 -7066
rect 540582 -7302 540666 -7066
rect 540902 -7302 540934 -7066
rect 540314 -7386 540934 -7302
rect 540314 -7622 540346 -7386
rect 540582 -7622 540666 -7386
rect 540902 -7622 540934 -7386
rect 540314 -7654 540934 -7622
rect 545434 -6106 546054 14058
rect 546834 709638 547454 709670
rect 546834 709402 546866 709638
rect 547102 709402 547186 709638
rect 547422 709402 547454 709638
rect 546834 709318 547454 709402
rect 546834 709082 546866 709318
rect 547102 709082 547186 709318
rect 547422 709082 547454 709318
rect 546834 676894 547454 709082
rect 546834 676658 546866 676894
rect 547102 676658 547186 676894
rect 547422 676658 547454 676894
rect 546834 676574 547454 676658
rect 546834 676338 546866 676574
rect 547102 676338 547186 676574
rect 547422 676338 547454 676574
rect 546834 640894 547454 676338
rect 546834 640658 546866 640894
rect 547102 640658 547186 640894
rect 547422 640658 547454 640894
rect 546834 640574 547454 640658
rect 546834 640338 546866 640574
rect 547102 640338 547186 640574
rect 547422 640338 547454 640574
rect 546834 604894 547454 640338
rect 546834 604658 546866 604894
rect 547102 604658 547186 604894
rect 547422 604658 547454 604894
rect 546834 604574 547454 604658
rect 546834 604338 546866 604574
rect 547102 604338 547186 604574
rect 547422 604338 547454 604574
rect 546834 568894 547454 604338
rect 546834 568658 546866 568894
rect 547102 568658 547186 568894
rect 547422 568658 547454 568894
rect 546834 568574 547454 568658
rect 546834 568338 546866 568574
rect 547102 568338 547186 568574
rect 547422 568338 547454 568574
rect 546834 532894 547454 568338
rect 546834 532658 546866 532894
rect 547102 532658 547186 532894
rect 547422 532658 547454 532894
rect 546834 532574 547454 532658
rect 546834 532338 546866 532574
rect 547102 532338 547186 532574
rect 547422 532338 547454 532574
rect 546834 496894 547454 532338
rect 546834 496658 546866 496894
rect 547102 496658 547186 496894
rect 547422 496658 547454 496894
rect 546834 496574 547454 496658
rect 546834 496338 546866 496574
rect 547102 496338 547186 496574
rect 547422 496338 547454 496574
rect 546834 460894 547454 496338
rect 546834 460658 546866 460894
rect 547102 460658 547186 460894
rect 547422 460658 547454 460894
rect 546834 460574 547454 460658
rect 546834 460338 546866 460574
rect 547102 460338 547186 460574
rect 547422 460338 547454 460574
rect 546834 424894 547454 460338
rect 546834 424658 546866 424894
rect 547102 424658 547186 424894
rect 547422 424658 547454 424894
rect 546834 424574 547454 424658
rect 546834 424338 546866 424574
rect 547102 424338 547186 424574
rect 547422 424338 547454 424574
rect 546834 388894 547454 424338
rect 546834 388658 546866 388894
rect 547102 388658 547186 388894
rect 547422 388658 547454 388894
rect 546834 388574 547454 388658
rect 546834 388338 546866 388574
rect 547102 388338 547186 388574
rect 547422 388338 547454 388574
rect 546834 352894 547454 388338
rect 546834 352658 546866 352894
rect 547102 352658 547186 352894
rect 547422 352658 547454 352894
rect 546834 352574 547454 352658
rect 546834 352338 546866 352574
rect 547102 352338 547186 352574
rect 547422 352338 547454 352574
rect 546834 316894 547454 352338
rect 546834 316658 546866 316894
rect 547102 316658 547186 316894
rect 547422 316658 547454 316894
rect 546834 316574 547454 316658
rect 546834 316338 546866 316574
rect 547102 316338 547186 316574
rect 547422 316338 547454 316574
rect 546834 280894 547454 316338
rect 546834 280658 546866 280894
rect 547102 280658 547186 280894
rect 547422 280658 547454 280894
rect 546834 280574 547454 280658
rect 546834 280338 546866 280574
rect 547102 280338 547186 280574
rect 547422 280338 547454 280574
rect 546834 244894 547454 280338
rect 546834 244658 546866 244894
rect 547102 244658 547186 244894
rect 547422 244658 547454 244894
rect 546834 244574 547454 244658
rect 546834 244338 546866 244574
rect 547102 244338 547186 244574
rect 547422 244338 547454 244574
rect 546834 208894 547454 244338
rect 546834 208658 546866 208894
rect 547102 208658 547186 208894
rect 547422 208658 547454 208894
rect 546834 208574 547454 208658
rect 546834 208338 546866 208574
rect 547102 208338 547186 208574
rect 547422 208338 547454 208574
rect 546834 172894 547454 208338
rect 546834 172658 546866 172894
rect 547102 172658 547186 172894
rect 547422 172658 547454 172894
rect 546834 172574 547454 172658
rect 546834 172338 546866 172574
rect 547102 172338 547186 172574
rect 547422 172338 547454 172574
rect 546834 136894 547454 172338
rect 546834 136658 546866 136894
rect 547102 136658 547186 136894
rect 547422 136658 547454 136894
rect 546834 136574 547454 136658
rect 546834 136338 546866 136574
rect 547102 136338 547186 136574
rect 547422 136338 547454 136574
rect 546834 100894 547454 136338
rect 546834 100658 546866 100894
rect 547102 100658 547186 100894
rect 547422 100658 547454 100894
rect 546834 100574 547454 100658
rect 546834 100338 546866 100574
rect 547102 100338 547186 100574
rect 547422 100338 547454 100574
rect 546834 64894 547454 100338
rect 546834 64658 546866 64894
rect 547102 64658 547186 64894
rect 547422 64658 547454 64894
rect 546834 64574 547454 64658
rect 546834 64338 546866 64574
rect 547102 64338 547186 64574
rect 547422 64338 547454 64574
rect 546834 28894 547454 64338
rect 546834 28658 546866 28894
rect 547102 28658 547186 28894
rect 547422 28658 547454 28894
rect 546834 28574 547454 28658
rect 546834 28338 546866 28574
rect 547102 28338 547186 28574
rect 547422 28338 547454 28574
rect 546834 -5146 547454 28338
rect 548234 706758 548854 707750
rect 548234 706522 548266 706758
rect 548502 706522 548586 706758
rect 548822 706522 548854 706758
rect 548234 706438 548854 706522
rect 548234 706202 548266 706438
rect 548502 706202 548586 706438
rect 548822 706202 548854 706438
rect 548234 691174 548854 706202
rect 548234 690938 548266 691174
rect 548502 690938 548586 691174
rect 548822 690938 548854 691174
rect 548234 690854 548854 690938
rect 548234 690618 548266 690854
rect 548502 690618 548586 690854
rect 548822 690618 548854 690854
rect 548234 655174 548854 690618
rect 548234 654938 548266 655174
rect 548502 654938 548586 655174
rect 548822 654938 548854 655174
rect 548234 654854 548854 654938
rect 548234 654618 548266 654854
rect 548502 654618 548586 654854
rect 548822 654618 548854 654854
rect 548234 619174 548854 654618
rect 548234 618938 548266 619174
rect 548502 618938 548586 619174
rect 548822 618938 548854 619174
rect 548234 618854 548854 618938
rect 548234 618618 548266 618854
rect 548502 618618 548586 618854
rect 548822 618618 548854 618854
rect 548234 583174 548854 618618
rect 548234 582938 548266 583174
rect 548502 582938 548586 583174
rect 548822 582938 548854 583174
rect 548234 582854 548854 582938
rect 548234 582618 548266 582854
rect 548502 582618 548586 582854
rect 548822 582618 548854 582854
rect 548234 547174 548854 582618
rect 548234 546938 548266 547174
rect 548502 546938 548586 547174
rect 548822 546938 548854 547174
rect 548234 546854 548854 546938
rect 548234 546618 548266 546854
rect 548502 546618 548586 546854
rect 548822 546618 548854 546854
rect 548234 511174 548854 546618
rect 548234 510938 548266 511174
rect 548502 510938 548586 511174
rect 548822 510938 548854 511174
rect 548234 510854 548854 510938
rect 548234 510618 548266 510854
rect 548502 510618 548586 510854
rect 548822 510618 548854 510854
rect 548234 475174 548854 510618
rect 548234 474938 548266 475174
rect 548502 474938 548586 475174
rect 548822 474938 548854 475174
rect 548234 474854 548854 474938
rect 548234 474618 548266 474854
rect 548502 474618 548586 474854
rect 548822 474618 548854 474854
rect 548234 439174 548854 474618
rect 548234 438938 548266 439174
rect 548502 438938 548586 439174
rect 548822 438938 548854 439174
rect 548234 438854 548854 438938
rect 548234 438618 548266 438854
rect 548502 438618 548586 438854
rect 548822 438618 548854 438854
rect 548234 403174 548854 438618
rect 548234 402938 548266 403174
rect 548502 402938 548586 403174
rect 548822 402938 548854 403174
rect 548234 402854 548854 402938
rect 548234 402618 548266 402854
rect 548502 402618 548586 402854
rect 548822 402618 548854 402854
rect 548234 367174 548854 402618
rect 548234 366938 548266 367174
rect 548502 366938 548586 367174
rect 548822 366938 548854 367174
rect 548234 366854 548854 366938
rect 548234 366618 548266 366854
rect 548502 366618 548586 366854
rect 548822 366618 548854 366854
rect 548234 331174 548854 366618
rect 548234 330938 548266 331174
rect 548502 330938 548586 331174
rect 548822 330938 548854 331174
rect 548234 330854 548854 330938
rect 548234 330618 548266 330854
rect 548502 330618 548586 330854
rect 548822 330618 548854 330854
rect 548234 295174 548854 330618
rect 548234 294938 548266 295174
rect 548502 294938 548586 295174
rect 548822 294938 548854 295174
rect 548234 294854 548854 294938
rect 548234 294618 548266 294854
rect 548502 294618 548586 294854
rect 548822 294618 548854 294854
rect 548234 259174 548854 294618
rect 548234 258938 548266 259174
rect 548502 258938 548586 259174
rect 548822 258938 548854 259174
rect 548234 258854 548854 258938
rect 548234 258618 548266 258854
rect 548502 258618 548586 258854
rect 548822 258618 548854 258854
rect 548234 223174 548854 258618
rect 548234 222938 548266 223174
rect 548502 222938 548586 223174
rect 548822 222938 548854 223174
rect 548234 222854 548854 222938
rect 548234 222618 548266 222854
rect 548502 222618 548586 222854
rect 548822 222618 548854 222854
rect 548234 187174 548854 222618
rect 548234 186938 548266 187174
rect 548502 186938 548586 187174
rect 548822 186938 548854 187174
rect 548234 186854 548854 186938
rect 548234 186618 548266 186854
rect 548502 186618 548586 186854
rect 548822 186618 548854 186854
rect 548234 151174 548854 186618
rect 548234 150938 548266 151174
rect 548502 150938 548586 151174
rect 548822 150938 548854 151174
rect 548234 150854 548854 150938
rect 548234 150618 548266 150854
rect 548502 150618 548586 150854
rect 548822 150618 548854 150854
rect 548234 115174 548854 150618
rect 548234 114938 548266 115174
rect 548502 114938 548586 115174
rect 548822 114938 548854 115174
rect 548234 114854 548854 114938
rect 548234 114618 548266 114854
rect 548502 114618 548586 114854
rect 548822 114618 548854 114854
rect 548234 79174 548854 114618
rect 548234 78938 548266 79174
rect 548502 78938 548586 79174
rect 548822 78938 548854 79174
rect 548234 78854 548854 78938
rect 548234 78618 548266 78854
rect 548502 78618 548586 78854
rect 548822 78618 548854 78854
rect 548234 43174 548854 78618
rect 548234 42938 548266 43174
rect 548502 42938 548586 43174
rect 548822 42938 548854 43174
rect 548234 42854 548854 42938
rect 548234 42618 548266 42854
rect 548502 42618 548586 42854
rect 548822 42618 548854 42854
rect 548234 7174 548854 42618
rect 548234 6938 548266 7174
rect 548502 6938 548586 7174
rect 548822 6938 548854 7174
rect 548234 6854 548854 6938
rect 548234 6618 548266 6854
rect 548502 6618 548586 6854
rect 548822 6618 548854 6854
rect 548234 -2266 548854 6618
rect 549634 705798 550254 705830
rect 549634 705562 549666 705798
rect 549902 705562 549986 705798
rect 550222 705562 550254 705798
rect 549634 705478 550254 705562
rect 549634 705242 549666 705478
rect 549902 705242 549986 705478
rect 550222 705242 550254 705478
rect 549634 669454 550254 705242
rect 549634 669218 549666 669454
rect 549902 669218 549986 669454
rect 550222 669218 550254 669454
rect 549634 669134 550254 669218
rect 549634 668898 549666 669134
rect 549902 668898 549986 669134
rect 550222 668898 550254 669134
rect 549634 633454 550254 668898
rect 549634 633218 549666 633454
rect 549902 633218 549986 633454
rect 550222 633218 550254 633454
rect 549634 633134 550254 633218
rect 549634 632898 549666 633134
rect 549902 632898 549986 633134
rect 550222 632898 550254 633134
rect 549634 597454 550254 632898
rect 549634 597218 549666 597454
rect 549902 597218 549986 597454
rect 550222 597218 550254 597454
rect 549634 597134 550254 597218
rect 549634 596898 549666 597134
rect 549902 596898 549986 597134
rect 550222 596898 550254 597134
rect 549634 561454 550254 596898
rect 549634 561218 549666 561454
rect 549902 561218 549986 561454
rect 550222 561218 550254 561454
rect 549634 561134 550254 561218
rect 549634 560898 549666 561134
rect 549902 560898 549986 561134
rect 550222 560898 550254 561134
rect 549634 525454 550254 560898
rect 549634 525218 549666 525454
rect 549902 525218 549986 525454
rect 550222 525218 550254 525454
rect 549634 525134 550254 525218
rect 549634 524898 549666 525134
rect 549902 524898 549986 525134
rect 550222 524898 550254 525134
rect 549634 489454 550254 524898
rect 549634 489218 549666 489454
rect 549902 489218 549986 489454
rect 550222 489218 550254 489454
rect 549634 489134 550254 489218
rect 549634 488898 549666 489134
rect 549902 488898 549986 489134
rect 550222 488898 550254 489134
rect 549634 453454 550254 488898
rect 549634 453218 549666 453454
rect 549902 453218 549986 453454
rect 550222 453218 550254 453454
rect 549634 453134 550254 453218
rect 549634 452898 549666 453134
rect 549902 452898 549986 453134
rect 550222 452898 550254 453134
rect 549634 417454 550254 452898
rect 549634 417218 549666 417454
rect 549902 417218 549986 417454
rect 550222 417218 550254 417454
rect 549634 417134 550254 417218
rect 549634 416898 549666 417134
rect 549902 416898 549986 417134
rect 550222 416898 550254 417134
rect 549634 381454 550254 416898
rect 549634 381218 549666 381454
rect 549902 381218 549986 381454
rect 550222 381218 550254 381454
rect 549634 381134 550254 381218
rect 549634 380898 549666 381134
rect 549902 380898 549986 381134
rect 550222 380898 550254 381134
rect 549634 345454 550254 380898
rect 549634 345218 549666 345454
rect 549902 345218 549986 345454
rect 550222 345218 550254 345454
rect 549634 345134 550254 345218
rect 549634 344898 549666 345134
rect 549902 344898 549986 345134
rect 550222 344898 550254 345134
rect 549634 309454 550254 344898
rect 549634 309218 549666 309454
rect 549902 309218 549986 309454
rect 550222 309218 550254 309454
rect 549634 309134 550254 309218
rect 549634 308898 549666 309134
rect 549902 308898 549986 309134
rect 550222 308898 550254 309134
rect 549634 273454 550254 308898
rect 549634 273218 549666 273454
rect 549902 273218 549986 273454
rect 550222 273218 550254 273454
rect 549634 273134 550254 273218
rect 549634 272898 549666 273134
rect 549902 272898 549986 273134
rect 550222 272898 550254 273134
rect 549634 237454 550254 272898
rect 549634 237218 549666 237454
rect 549902 237218 549986 237454
rect 550222 237218 550254 237454
rect 549634 237134 550254 237218
rect 549634 236898 549666 237134
rect 549902 236898 549986 237134
rect 550222 236898 550254 237134
rect 549634 201454 550254 236898
rect 549634 201218 549666 201454
rect 549902 201218 549986 201454
rect 550222 201218 550254 201454
rect 549634 201134 550254 201218
rect 549634 200898 549666 201134
rect 549902 200898 549986 201134
rect 550222 200898 550254 201134
rect 549634 165454 550254 200898
rect 549634 165218 549666 165454
rect 549902 165218 549986 165454
rect 550222 165218 550254 165454
rect 549634 165134 550254 165218
rect 549634 164898 549666 165134
rect 549902 164898 549986 165134
rect 550222 164898 550254 165134
rect 549634 129454 550254 164898
rect 549634 129218 549666 129454
rect 549902 129218 549986 129454
rect 550222 129218 550254 129454
rect 549634 129134 550254 129218
rect 549634 128898 549666 129134
rect 549902 128898 549986 129134
rect 550222 128898 550254 129134
rect 549634 93454 550254 128898
rect 549634 93218 549666 93454
rect 549902 93218 549986 93454
rect 550222 93218 550254 93454
rect 549634 93134 550254 93218
rect 549634 92898 549666 93134
rect 549902 92898 549986 93134
rect 550222 92898 550254 93134
rect 549634 57454 550254 92898
rect 549634 57218 549666 57454
rect 549902 57218 549986 57454
rect 550222 57218 550254 57454
rect 549634 57134 550254 57218
rect 549634 56898 549666 57134
rect 549902 56898 549986 57134
rect 550222 56898 550254 57134
rect 549634 21454 550254 56898
rect 549634 21218 549666 21454
rect 549902 21218 549986 21454
rect 550222 21218 550254 21454
rect 549634 21134 550254 21218
rect 549634 20898 549666 21134
rect 549902 20898 549986 21134
rect 550222 20898 550254 21134
rect 549634 -1306 550254 20898
rect 549634 -1542 549666 -1306
rect 549902 -1542 549986 -1306
rect 550222 -1542 550254 -1306
rect 549634 -1626 550254 -1542
rect 549634 -1862 549666 -1626
rect 549902 -1862 549986 -1626
rect 550222 -1862 550254 -1626
rect 549634 -1894 550254 -1862
rect 550554 680614 551174 711002
rect 555674 710598 556294 711590
rect 555674 710362 555706 710598
rect 555942 710362 556026 710598
rect 556262 710362 556294 710598
rect 555674 710278 556294 710362
rect 555674 710042 555706 710278
rect 555942 710042 556026 710278
rect 556262 710042 556294 710278
rect 550554 680378 550586 680614
rect 550822 680378 550906 680614
rect 551142 680378 551174 680614
rect 550554 680294 551174 680378
rect 550554 680058 550586 680294
rect 550822 680058 550906 680294
rect 551142 680058 551174 680294
rect 550554 644614 551174 680058
rect 550554 644378 550586 644614
rect 550822 644378 550906 644614
rect 551142 644378 551174 644614
rect 550554 644294 551174 644378
rect 550554 644058 550586 644294
rect 550822 644058 550906 644294
rect 551142 644058 551174 644294
rect 550554 608614 551174 644058
rect 550554 608378 550586 608614
rect 550822 608378 550906 608614
rect 551142 608378 551174 608614
rect 550554 608294 551174 608378
rect 550554 608058 550586 608294
rect 550822 608058 550906 608294
rect 551142 608058 551174 608294
rect 550554 572614 551174 608058
rect 550554 572378 550586 572614
rect 550822 572378 550906 572614
rect 551142 572378 551174 572614
rect 550554 572294 551174 572378
rect 550554 572058 550586 572294
rect 550822 572058 550906 572294
rect 551142 572058 551174 572294
rect 550554 536614 551174 572058
rect 550554 536378 550586 536614
rect 550822 536378 550906 536614
rect 551142 536378 551174 536614
rect 550554 536294 551174 536378
rect 550554 536058 550586 536294
rect 550822 536058 550906 536294
rect 551142 536058 551174 536294
rect 550554 500614 551174 536058
rect 550554 500378 550586 500614
rect 550822 500378 550906 500614
rect 551142 500378 551174 500614
rect 550554 500294 551174 500378
rect 550554 500058 550586 500294
rect 550822 500058 550906 500294
rect 551142 500058 551174 500294
rect 550554 464614 551174 500058
rect 550554 464378 550586 464614
rect 550822 464378 550906 464614
rect 551142 464378 551174 464614
rect 550554 464294 551174 464378
rect 550554 464058 550586 464294
rect 550822 464058 550906 464294
rect 551142 464058 551174 464294
rect 550554 428614 551174 464058
rect 550554 428378 550586 428614
rect 550822 428378 550906 428614
rect 551142 428378 551174 428614
rect 550554 428294 551174 428378
rect 550554 428058 550586 428294
rect 550822 428058 550906 428294
rect 551142 428058 551174 428294
rect 550554 392614 551174 428058
rect 550554 392378 550586 392614
rect 550822 392378 550906 392614
rect 551142 392378 551174 392614
rect 550554 392294 551174 392378
rect 550554 392058 550586 392294
rect 550822 392058 550906 392294
rect 551142 392058 551174 392294
rect 550554 356614 551174 392058
rect 550554 356378 550586 356614
rect 550822 356378 550906 356614
rect 551142 356378 551174 356614
rect 550554 356294 551174 356378
rect 550554 356058 550586 356294
rect 550822 356058 550906 356294
rect 551142 356058 551174 356294
rect 550554 320614 551174 356058
rect 550554 320378 550586 320614
rect 550822 320378 550906 320614
rect 551142 320378 551174 320614
rect 550554 320294 551174 320378
rect 550554 320058 550586 320294
rect 550822 320058 550906 320294
rect 551142 320058 551174 320294
rect 550554 284614 551174 320058
rect 550554 284378 550586 284614
rect 550822 284378 550906 284614
rect 551142 284378 551174 284614
rect 550554 284294 551174 284378
rect 550554 284058 550586 284294
rect 550822 284058 550906 284294
rect 551142 284058 551174 284294
rect 550554 248614 551174 284058
rect 550554 248378 550586 248614
rect 550822 248378 550906 248614
rect 551142 248378 551174 248614
rect 550554 248294 551174 248378
rect 550554 248058 550586 248294
rect 550822 248058 550906 248294
rect 551142 248058 551174 248294
rect 550554 212614 551174 248058
rect 550554 212378 550586 212614
rect 550822 212378 550906 212614
rect 551142 212378 551174 212614
rect 550554 212294 551174 212378
rect 550554 212058 550586 212294
rect 550822 212058 550906 212294
rect 551142 212058 551174 212294
rect 550554 176614 551174 212058
rect 550554 176378 550586 176614
rect 550822 176378 550906 176614
rect 551142 176378 551174 176614
rect 550554 176294 551174 176378
rect 550554 176058 550586 176294
rect 550822 176058 550906 176294
rect 551142 176058 551174 176294
rect 550554 140614 551174 176058
rect 550554 140378 550586 140614
rect 550822 140378 550906 140614
rect 551142 140378 551174 140614
rect 550554 140294 551174 140378
rect 550554 140058 550586 140294
rect 550822 140058 550906 140294
rect 551142 140058 551174 140294
rect 550554 104614 551174 140058
rect 550554 104378 550586 104614
rect 550822 104378 550906 104614
rect 551142 104378 551174 104614
rect 550554 104294 551174 104378
rect 550554 104058 550586 104294
rect 550822 104058 550906 104294
rect 551142 104058 551174 104294
rect 550554 68614 551174 104058
rect 550554 68378 550586 68614
rect 550822 68378 550906 68614
rect 551142 68378 551174 68614
rect 550554 68294 551174 68378
rect 550554 68058 550586 68294
rect 550822 68058 550906 68294
rect 551142 68058 551174 68294
rect 550554 32614 551174 68058
rect 550554 32378 550586 32614
rect 550822 32378 550906 32614
rect 551142 32378 551174 32614
rect 550554 32294 551174 32378
rect 550554 32058 550586 32294
rect 550822 32058 550906 32294
rect 551142 32058 551174 32294
rect 548234 -2502 548266 -2266
rect 548502 -2502 548586 -2266
rect 548822 -2502 548854 -2266
rect 548234 -2586 548854 -2502
rect 548234 -2822 548266 -2586
rect 548502 -2822 548586 -2586
rect 548822 -2822 548854 -2586
rect 548234 -3814 548854 -2822
rect 546834 -5382 546866 -5146
rect 547102 -5382 547186 -5146
rect 547422 -5382 547454 -5146
rect 546834 -5466 547454 -5382
rect 546834 -5702 546866 -5466
rect 547102 -5702 547186 -5466
rect 547422 -5702 547454 -5466
rect 546834 -5734 547454 -5702
rect 545434 -6342 545466 -6106
rect 545702 -6342 545786 -6106
rect 546022 -6342 546054 -6106
rect 545434 -6426 546054 -6342
rect 545434 -6662 545466 -6426
rect 545702 -6662 545786 -6426
rect 546022 -6662 546054 -6426
rect 545434 -7654 546054 -6662
rect 550554 -7066 551174 32058
rect 551954 708678 552574 709670
rect 551954 708442 551986 708678
rect 552222 708442 552306 708678
rect 552542 708442 552574 708678
rect 551954 708358 552574 708442
rect 551954 708122 551986 708358
rect 552222 708122 552306 708358
rect 552542 708122 552574 708358
rect 551954 694894 552574 708122
rect 551954 694658 551986 694894
rect 552222 694658 552306 694894
rect 552542 694658 552574 694894
rect 551954 694574 552574 694658
rect 551954 694338 551986 694574
rect 552222 694338 552306 694574
rect 552542 694338 552574 694574
rect 551954 658894 552574 694338
rect 551954 658658 551986 658894
rect 552222 658658 552306 658894
rect 552542 658658 552574 658894
rect 551954 658574 552574 658658
rect 551954 658338 551986 658574
rect 552222 658338 552306 658574
rect 552542 658338 552574 658574
rect 551954 622894 552574 658338
rect 551954 622658 551986 622894
rect 552222 622658 552306 622894
rect 552542 622658 552574 622894
rect 551954 622574 552574 622658
rect 551954 622338 551986 622574
rect 552222 622338 552306 622574
rect 552542 622338 552574 622574
rect 551954 586894 552574 622338
rect 551954 586658 551986 586894
rect 552222 586658 552306 586894
rect 552542 586658 552574 586894
rect 551954 586574 552574 586658
rect 551954 586338 551986 586574
rect 552222 586338 552306 586574
rect 552542 586338 552574 586574
rect 551954 550894 552574 586338
rect 551954 550658 551986 550894
rect 552222 550658 552306 550894
rect 552542 550658 552574 550894
rect 551954 550574 552574 550658
rect 551954 550338 551986 550574
rect 552222 550338 552306 550574
rect 552542 550338 552574 550574
rect 551954 514894 552574 550338
rect 551954 514658 551986 514894
rect 552222 514658 552306 514894
rect 552542 514658 552574 514894
rect 551954 514574 552574 514658
rect 551954 514338 551986 514574
rect 552222 514338 552306 514574
rect 552542 514338 552574 514574
rect 551954 478894 552574 514338
rect 551954 478658 551986 478894
rect 552222 478658 552306 478894
rect 552542 478658 552574 478894
rect 551954 478574 552574 478658
rect 551954 478338 551986 478574
rect 552222 478338 552306 478574
rect 552542 478338 552574 478574
rect 551954 442894 552574 478338
rect 551954 442658 551986 442894
rect 552222 442658 552306 442894
rect 552542 442658 552574 442894
rect 551954 442574 552574 442658
rect 551954 442338 551986 442574
rect 552222 442338 552306 442574
rect 552542 442338 552574 442574
rect 551954 406894 552574 442338
rect 551954 406658 551986 406894
rect 552222 406658 552306 406894
rect 552542 406658 552574 406894
rect 551954 406574 552574 406658
rect 551954 406338 551986 406574
rect 552222 406338 552306 406574
rect 552542 406338 552574 406574
rect 551954 370894 552574 406338
rect 551954 370658 551986 370894
rect 552222 370658 552306 370894
rect 552542 370658 552574 370894
rect 551954 370574 552574 370658
rect 551954 370338 551986 370574
rect 552222 370338 552306 370574
rect 552542 370338 552574 370574
rect 551954 334894 552574 370338
rect 551954 334658 551986 334894
rect 552222 334658 552306 334894
rect 552542 334658 552574 334894
rect 551954 334574 552574 334658
rect 551954 334338 551986 334574
rect 552222 334338 552306 334574
rect 552542 334338 552574 334574
rect 551954 298894 552574 334338
rect 551954 298658 551986 298894
rect 552222 298658 552306 298894
rect 552542 298658 552574 298894
rect 551954 298574 552574 298658
rect 551954 298338 551986 298574
rect 552222 298338 552306 298574
rect 552542 298338 552574 298574
rect 551954 262894 552574 298338
rect 551954 262658 551986 262894
rect 552222 262658 552306 262894
rect 552542 262658 552574 262894
rect 551954 262574 552574 262658
rect 551954 262338 551986 262574
rect 552222 262338 552306 262574
rect 552542 262338 552574 262574
rect 551954 226894 552574 262338
rect 551954 226658 551986 226894
rect 552222 226658 552306 226894
rect 552542 226658 552574 226894
rect 551954 226574 552574 226658
rect 551954 226338 551986 226574
rect 552222 226338 552306 226574
rect 552542 226338 552574 226574
rect 551954 190894 552574 226338
rect 551954 190658 551986 190894
rect 552222 190658 552306 190894
rect 552542 190658 552574 190894
rect 551954 190574 552574 190658
rect 551954 190338 551986 190574
rect 552222 190338 552306 190574
rect 552542 190338 552574 190574
rect 551954 154894 552574 190338
rect 551954 154658 551986 154894
rect 552222 154658 552306 154894
rect 552542 154658 552574 154894
rect 551954 154574 552574 154658
rect 551954 154338 551986 154574
rect 552222 154338 552306 154574
rect 552542 154338 552574 154574
rect 551954 118894 552574 154338
rect 551954 118658 551986 118894
rect 552222 118658 552306 118894
rect 552542 118658 552574 118894
rect 551954 118574 552574 118658
rect 551954 118338 551986 118574
rect 552222 118338 552306 118574
rect 552542 118338 552574 118574
rect 551954 82894 552574 118338
rect 551954 82658 551986 82894
rect 552222 82658 552306 82894
rect 552542 82658 552574 82894
rect 551954 82574 552574 82658
rect 551954 82338 551986 82574
rect 552222 82338 552306 82574
rect 552542 82338 552574 82574
rect 551954 46894 552574 82338
rect 551954 46658 551986 46894
rect 552222 46658 552306 46894
rect 552542 46658 552574 46894
rect 551954 46574 552574 46658
rect 551954 46338 551986 46574
rect 552222 46338 552306 46574
rect 552542 46338 552574 46574
rect 551954 10894 552574 46338
rect 551954 10658 551986 10894
rect 552222 10658 552306 10894
rect 552542 10658 552574 10894
rect 551954 10574 552574 10658
rect 551954 10338 551986 10574
rect 552222 10338 552306 10574
rect 552542 10338 552574 10574
rect 551954 -4186 552574 10338
rect 553354 707718 553974 707750
rect 553354 707482 553386 707718
rect 553622 707482 553706 707718
rect 553942 707482 553974 707718
rect 553354 707398 553974 707482
rect 553354 707162 553386 707398
rect 553622 707162 553706 707398
rect 553942 707162 553974 707398
rect 553354 673174 553974 707162
rect 553354 672938 553386 673174
rect 553622 672938 553706 673174
rect 553942 672938 553974 673174
rect 553354 672854 553974 672938
rect 553354 672618 553386 672854
rect 553622 672618 553706 672854
rect 553942 672618 553974 672854
rect 553354 637174 553974 672618
rect 553354 636938 553386 637174
rect 553622 636938 553706 637174
rect 553942 636938 553974 637174
rect 553354 636854 553974 636938
rect 553354 636618 553386 636854
rect 553622 636618 553706 636854
rect 553942 636618 553974 636854
rect 553354 601174 553974 636618
rect 553354 600938 553386 601174
rect 553622 600938 553706 601174
rect 553942 600938 553974 601174
rect 553354 600854 553974 600938
rect 553354 600618 553386 600854
rect 553622 600618 553706 600854
rect 553942 600618 553974 600854
rect 553354 565174 553974 600618
rect 553354 564938 553386 565174
rect 553622 564938 553706 565174
rect 553942 564938 553974 565174
rect 553354 564854 553974 564938
rect 553354 564618 553386 564854
rect 553622 564618 553706 564854
rect 553942 564618 553974 564854
rect 553354 529174 553974 564618
rect 553354 528938 553386 529174
rect 553622 528938 553706 529174
rect 553942 528938 553974 529174
rect 553354 528854 553974 528938
rect 553354 528618 553386 528854
rect 553622 528618 553706 528854
rect 553942 528618 553974 528854
rect 553354 493174 553974 528618
rect 553354 492938 553386 493174
rect 553622 492938 553706 493174
rect 553942 492938 553974 493174
rect 553354 492854 553974 492938
rect 553354 492618 553386 492854
rect 553622 492618 553706 492854
rect 553942 492618 553974 492854
rect 553354 457174 553974 492618
rect 553354 456938 553386 457174
rect 553622 456938 553706 457174
rect 553942 456938 553974 457174
rect 553354 456854 553974 456938
rect 553354 456618 553386 456854
rect 553622 456618 553706 456854
rect 553942 456618 553974 456854
rect 553354 421174 553974 456618
rect 553354 420938 553386 421174
rect 553622 420938 553706 421174
rect 553942 420938 553974 421174
rect 553354 420854 553974 420938
rect 553354 420618 553386 420854
rect 553622 420618 553706 420854
rect 553942 420618 553974 420854
rect 553354 385174 553974 420618
rect 553354 384938 553386 385174
rect 553622 384938 553706 385174
rect 553942 384938 553974 385174
rect 553354 384854 553974 384938
rect 553354 384618 553386 384854
rect 553622 384618 553706 384854
rect 553942 384618 553974 384854
rect 553354 349174 553974 384618
rect 553354 348938 553386 349174
rect 553622 348938 553706 349174
rect 553942 348938 553974 349174
rect 553354 348854 553974 348938
rect 553354 348618 553386 348854
rect 553622 348618 553706 348854
rect 553942 348618 553974 348854
rect 553354 313174 553974 348618
rect 553354 312938 553386 313174
rect 553622 312938 553706 313174
rect 553942 312938 553974 313174
rect 553354 312854 553974 312938
rect 553354 312618 553386 312854
rect 553622 312618 553706 312854
rect 553942 312618 553974 312854
rect 553354 277174 553974 312618
rect 553354 276938 553386 277174
rect 553622 276938 553706 277174
rect 553942 276938 553974 277174
rect 553354 276854 553974 276938
rect 553354 276618 553386 276854
rect 553622 276618 553706 276854
rect 553942 276618 553974 276854
rect 553354 241174 553974 276618
rect 553354 240938 553386 241174
rect 553622 240938 553706 241174
rect 553942 240938 553974 241174
rect 553354 240854 553974 240938
rect 553354 240618 553386 240854
rect 553622 240618 553706 240854
rect 553942 240618 553974 240854
rect 553354 205174 553974 240618
rect 553354 204938 553386 205174
rect 553622 204938 553706 205174
rect 553942 204938 553974 205174
rect 553354 204854 553974 204938
rect 553354 204618 553386 204854
rect 553622 204618 553706 204854
rect 553942 204618 553974 204854
rect 553354 169174 553974 204618
rect 553354 168938 553386 169174
rect 553622 168938 553706 169174
rect 553942 168938 553974 169174
rect 553354 168854 553974 168938
rect 553354 168618 553386 168854
rect 553622 168618 553706 168854
rect 553942 168618 553974 168854
rect 553354 133174 553974 168618
rect 553354 132938 553386 133174
rect 553622 132938 553706 133174
rect 553942 132938 553974 133174
rect 553354 132854 553974 132938
rect 553354 132618 553386 132854
rect 553622 132618 553706 132854
rect 553942 132618 553974 132854
rect 553354 97174 553974 132618
rect 553354 96938 553386 97174
rect 553622 96938 553706 97174
rect 553942 96938 553974 97174
rect 553354 96854 553974 96938
rect 553354 96618 553386 96854
rect 553622 96618 553706 96854
rect 553942 96618 553974 96854
rect 553354 61174 553974 96618
rect 553354 60938 553386 61174
rect 553622 60938 553706 61174
rect 553942 60938 553974 61174
rect 553354 60854 553974 60938
rect 553354 60618 553386 60854
rect 553622 60618 553706 60854
rect 553942 60618 553974 60854
rect 553354 25174 553974 60618
rect 553354 24938 553386 25174
rect 553622 24938 553706 25174
rect 553942 24938 553974 25174
rect 553354 24854 553974 24938
rect 553354 24618 553386 24854
rect 553622 24618 553706 24854
rect 553942 24618 553974 24854
rect 553354 -3226 553974 24618
rect 554754 704838 555374 705830
rect 554754 704602 554786 704838
rect 555022 704602 555106 704838
rect 555342 704602 555374 704838
rect 554754 704518 555374 704602
rect 554754 704282 554786 704518
rect 555022 704282 555106 704518
rect 555342 704282 555374 704518
rect 554754 687454 555374 704282
rect 554754 687218 554786 687454
rect 555022 687218 555106 687454
rect 555342 687218 555374 687454
rect 554754 687134 555374 687218
rect 554754 686898 554786 687134
rect 555022 686898 555106 687134
rect 555342 686898 555374 687134
rect 554754 651454 555374 686898
rect 554754 651218 554786 651454
rect 555022 651218 555106 651454
rect 555342 651218 555374 651454
rect 554754 651134 555374 651218
rect 554754 650898 554786 651134
rect 555022 650898 555106 651134
rect 555342 650898 555374 651134
rect 554754 615454 555374 650898
rect 554754 615218 554786 615454
rect 555022 615218 555106 615454
rect 555342 615218 555374 615454
rect 554754 615134 555374 615218
rect 554754 614898 554786 615134
rect 555022 614898 555106 615134
rect 555342 614898 555374 615134
rect 554754 579454 555374 614898
rect 554754 579218 554786 579454
rect 555022 579218 555106 579454
rect 555342 579218 555374 579454
rect 554754 579134 555374 579218
rect 554754 578898 554786 579134
rect 555022 578898 555106 579134
rect 555342 578898 555374 579134
rect 554754 543454 555374 578898
rect 554754 543218 554786 543454
rect 555022 543218 555106 543454
rect 555342 543218 555374 543454
rect 554754 543134 555374 543218
rect 554754 542898 554786 543134
rect 555022 542898 555106 543134
rect 555342 542898 555374 543134
rect 554754 507454 555374 542898
rect 554754 507218 554786 507454
rect 555022 507218 555106 507454
rect 555342 507218 555374 507454
rect 554754 507134 555374 507218
rect 554754 506898 554786 507134
rect 555022 506898 555106 507134
rect 555342 506898 555374 507134
rect 554754 471454 555374 506898
rect 554754 471218 554786 471454
rect 555022 471218 555106 471454
rect 555342 471218 555374 471454
rect 554754 471134 555374 471218
rect 554754 470898 554786 471134
rect 555022 470898 555106 471134
rect 555342 470898 555374 471134
rect 554754 435454 555374 470898
rect 554754 435218 554786 435454
rect 555022 435218 555106 435454
rect 555342 435218 555374 435454
rect 554754 435134 555374 435218
rect 554754 434898 554786 435134
rect 555022 434898 555106 435134
rect 555342 434898 555374 435134
rect 554754 399454 555374 434898
rect 554754 399218 554786 399454
rect 555022 399218 555106 399454
rect 555342 399218 555374 399454
rect 554754 399134 555374 399218
rect 554754 398898 554786 399134
rect 555022 398898 555106 399134
rect 555342 398898 555374 399134
rect 554754 363454 555374 398898
rect 554754 363218 554786 363454
rect 555022 363218 555106 363454
rect 555342 363218 555374 363454
rect 554754 363134 555374 363218
rect 554754 362898 554786 363134
rect 555022 362898 555106 363134
rect 555342 362898 555374 363134
rect 554754 327454 555374 362898
rect 554754 327218 554786 327454
rect 555022 327218 555106 327454
rect 555342 327218 555374 327454
rect 554754 327134 555374 327218
rect 554754 326898 554786 327134
rect 555022 326898 555106 327134
rect 555342 326898 555374 327134
rect 554754 291454 555374 326898
rect 554754 291218 554786 291454
rect 555022 291218 555106 291454
rect 555342 291218 555374 291454
rect 554754 291134 555374 291218
rect 554754 290898 554786 291134
rect 555022 290898 555106 291134
rect 555342 290898 555374 291134
rect 554754 255454 555374 290898
rect 554754 255218 554786 255454
rect 555022 255218 555106 255454
rect 555342 255218 555374 255454
rect 554754 255134 555374 255218
rect 554754 254898 554786 255134
rect 555022 254898 555106 255134
rect 555342 254898 555374 255134
rect 554754 219454 555374 254898
rect 554754 219218 554786 219454
rect 555022 219218 555106 219454
rect 555342 219218 555374 219454
rect 554754 219134 555374 219218
rect 554754 218898 554786 219134
rect 555022 218898 555106 219134
rect 555342 218898 555374 219134
rect 554754 183454 555374 218898
rect 554754 183218 554786 183454
rect 555022 183218 555106 183454
rect 555342 183218 555374 183454
rect 554754 183134 555374 183218
rect 554754 182898 554786 183134
rect 555022 182898 555106 183134
rect 555342 182898 555374 183134
rect 554754 147454 555374 182898
rect 554754 147218 554786 147454
rect 555022 147218 555106 147454
rect 555342 147218 555374 147454
rect 554754 147134 555374 147218
rect 554754 146898 554786 147134
rect 555022 146898 555106 147134
rect 555342 146898 555374 147134
rect 554754 111454 555374 146898
rect 554754 111218 554786 111454
rect 555022 111218 555106 111454
rect 555342 111218 555374 111454
rect 554754 111134 555374 111218
rect 554754 110898 554786 111134
rect 555022 110898 555106 111134
rect 555342 110898 555374 111134
rect 554754 75454 555374 110898
rect 554754 75218 554786 75454
rect 555022 75218 555106 75454
rect 555342 75218 555374 75454
rect 554754 75134 555374 75218
rect 554754 74898 554786 75134
rect 555022 74898 555106 75134
rect 555342 74898 555374 75134
rect 554754 39454 555374 74898
rect 554754 39218 554786 39454
rect 555022 39218 555106 39454
rect 555342 39218 555374 39454
rect 554754 39134 555374 39218
rect 554754 38898 554786 39134
rect 555022 38898 555106 39134
rect 555342 38898 555374 39134
rect 554754 3454 555374 38898
rect 554754 3218 554786 3454
rect 555022 3218 555106 3454
rect 555342 3218 555374 3454
rect 554754 3134 555374 3218
rect 554754 2898 554786 3134
rect 555022 2898 555106 3134
rect 555342 2898 555374 3134
rect 554754 -346 555374 2898
rect 554754 -582 554786 -346
rect 555022 -582 555106 -346
rect 555342 -582 555374 -346
rect 554754 -666 555374 -582
rect 554754 -902 554786 -666
rect 555022 -902 555106 -666
rect 555342 -902 555374 -666
rect 554754 -1894 555374 -902
rect 555674 698614 556294 710042
rect 560794 711558 561414 711590
rect 560794 711322 560826 711558
rect 561062 711322 561146 711558
rect 561382 711322 561414 711558
rect 560794 711238 561414 711322
rect 560794 711002 560826 711238
rect 561062 711002 561146 711238
rect 561382 711002 561414 711238
rect 555674 698378 555706 698614
rect 555942 698378 556026 698614
rect 556262 698378 556294 698614
rect 555674 698294 556294 698378
rect 555674 698058 555706 698294
rect 555942 698058 556026 698294
rect 556262 698058 556294 698294
rect 555674 662614 556294 698058
rect 555674 662378 555706 662614
rect 555942 662378 556026 662614
rect 556262 662378 556294 662614
rect 555674 662294 556294 662378
rect 555674 662058 555706 662294
rect 555942 662058 556026 662294
rect 556262 662058 556294 662294
rect 555674 626614 556294 662058
rect 555674 626378 555706 626614
rect 555942 626378 556026 626614
rect 556262 626378 556294 626614
rect 555674 626294 556294 626378
rect 555674 626058 555706 626294
rect 555942 626058 556026 626294
rect 556262 626058 556294 626294
rect 555674 590614 556294 626058
rect 555674 590378 555706 590614
rect 555942 590378 556026 590614
rect 556262 590378 556294 590614
rect 555674 590294 556294 590378
rect 555674 590058 555706 590294
rect 555942 590058 556026 590294
rect 556262 590058 556294 590294
rect 555674 554614 556294 590058
rect 555674 554378 555706 554614
rect 555942 554378 556026 554614
rect 556262 554378 556294 554614
rect 555674 554294 556294 554378
rect 555674 554058 555706 554294
rect 555942 554058 556026 554294
rect 556262 554058 556294 554294
rect 555674 518614 556294 554058
rect 555674 518378 555706 518614
rect 555942 518378 556026 518614
rect 556262 518378 556294 518614
rect 555674 518294 556294 518378
rect 555674 518058 555706 518294
rect 555942 518058 556026 518294
rect 556262 518058 556294 518294
rect 555674 482614 556294 518058
rect 555674 482378 555706 482614
rect 555942 482378 556026 482614
rect 556262 482378 556294 482614
rect 555674 482294 556294 482378
rect 555674 482058 555706 482294
rect 555942 482058 556026 482294
rect 556262 482058 556294 482294
rect 555674 446614 556294 482058
rect 555674 446378 555706 446614
rect 555942 446378 556026 446614
rect 556262 446378 556294 446614
rect 555674 446294 556294 446378
rect 555674 446058 555706 446294
rect 555942 446058 556026 446294
rect 556262 446058 556294 446294
rect 555674 410614 556294 446058
rect 555674 410378 555706 410614
rect 555942 410378 556026 410614
rect 556262 410378 556294 410614
rect 555674 410294 556294 410378
rect 555674 410058 555706 410294
rect 555942 410058 556026 410294
rect 556262 410058 556294 410294
rect 555674 374614 556294 410058
rect 555674 374378 555706 374614
rect 555942 374378 556026 374614
rect 556262 374378 556294 374614
rect 555674 374294 556294 374378
rect 555674 374058 555706 374294
rect 555942 374058 556026 374294
rect 556262 374058 556294 374294
rect 555674 338614 556294 374058
rect 555674 338378 555706 338614
rect 555942 338378 556026 338614
rect 556262 338378 556294 338614
rect 555674 338294 556294 338378
rect 555674 338058 555706 338294
rect 555942 338058 556026 338294
rect 556262 338058 556294 338294
rect 555674 302614 556294 338058
rect 555674 302378 555706 302614
rect 555942 302378 556026 302614
rect 556262 302378 556294 302614
rect 555674 302294 556294 302378
rect 555674 302058 555706 302294
rect 555942 302058 556026 302294
rect 556262 302058 556294 302294
rect 555674 266614 556294 302058
rect 555674 266378 555706 266614
rect 555942 266378 556026 266614
rect 556262 266378 556294 266614
rect 555674 266294 556294 266378
rect 555674 266058 555706 266294
rect 555942 266058 556026 266294
rect 556262 266058 556294 266294
rect 555674 230614 556294 266058
rect 555674 230378 555706 230614
rect 555942 230378 556026 230614
rect 556262 230378 556294 230614
rect 555674 230294 556294 230378
rect 555674 230058 555706 230294
rect 555942 230058 556026 230294
rect 556262 230058 556294 230294
rect 555674 194614 556294 230058
rect 555674 194378 555706 194614
rect 555942 194378 556026 194614
rect 556262 194378 556294 194614
rect 555674 194294 556294 194378
rect 555674 194058 555706 194294
rect 555942 194058 556026 194294
rect 556262 194058 556294 194294
rect 555674 158614 556294 194058
rect 555674 158378 555706 158614
rect 555942 158378 556026 158614
rect 556262 158378 556294 158614
rect 555674 158294 556294 158378
rect 555674 158058 555706 158294
rect 555942 158058 556026 158294
rect 556262 158058 556294 158294
rect 555674 122614 556294 158058
rect 555674 122378 555706 122614
rect 555942 122378 556026 122614
rect 556262 122378 556294 122614
rect 555674 122294 556294 122378
rect 555674 122058 555706 122294
rect 555942 122058 556026 122294
rect 556262 122058 556294 122294
rect 555674 86614 556294 122058
rect 555674 86378 555706 86614
rect 555942 86378 556026 86614
rect 556262 86378 556294 86614
rect 555674 86294 556294 86378
rect 555674 86058 555706 86294
rect 555942 86058 556026 86294
rect 556262 86058 556294 86294
rect 555674 50614 556294 86058
rect 555674 50378 555706 50614
rect 555942 50378 556026 50614
rect 556262 50378 556294 50614
rect 555674 50294 556294 50378
rect 555674 50058 555706 50294
rect 555942 50058 556026 50294
rect 556262 50058 556294 50294
rect 555674 14614 556294 50058
rect 555674 14378 555706 14614
rect 555942 14378 556026 14614
rect 556262 14378 556294 14614
rect 555674 14294 556294 14378
rect 555674 14058 555706 14294
rect 555942 14058 556026 14294
rect 556262 14058 556294 14294
rect 553354 -3462 553386 -3226
rect 553622 -3462 553706 -3226
rect 553942 -3462 553974 -3226
rect 553354 -3546 553974 -3462
rect 553354 -3782 553386 -3546
rect 553622 -3782 553706 -3546
rect 553942 -3782 553974 -3546
rect 553354 -3814 553974 -3782
rect 551954 -4422 551986 -4186
rect 552222 -4422 552306 -4186
rect 552542 -4422 552574 -4186
rect 551954 -4506 552574 -4422
rect 551954 -4742 551986 -4506
rect 552222 -4742 552306 -4506
rect 552542 -4742 552574 -4506
rect 551954 -5734 552574 -4742
rect 550554 -7302 550586 -7066
rect 550822 -7302 550906 -7066
rect 551142 -7302 551174 -7066
rect 550554 -7386 551174 -7302
rect 550554 -7622 550586 -7386
rect 550822 -7622 550906 -7386
rect 551142 -7622 551174 -7386
rect 550554 -7654 551174 -7622
rect 555674 -6106 556294 14058
rect 557074 709638 557694 709670
rect 557074 709402 557106 709638
rect 557342 709402 557426 709638
rect 557662 709402 557694 709638
rect 557074 709318 557694 709402
rect 557074 709082 557106 709318
rect 557342 709082 557426 709318
rect 557662 709082 557694 709318
rect 557074 676894 557694 709082
rect 557074 676658 557106 676894
rect 557342 676658 557426 676894
rect 557662 676658 557694 676894
rect 557074 676574 557694 676658
rect 557074 676338 557106 676574
rect 557342 676338 557426 676574
rect 557662 676338 557694 676574
rect 557074 640894 557694 676338
rect 557074 640658 557106 640894
rect 557342 640658 557426 640894
rect 557662 640658 557694 640894
rect 557074 640574 557694 640658
rect 557074 640338 557106 640574
rect 557342 640338 557426 640574
rect 557662 640338 557694 640574
rect 557074 604894 557694 640338
rect 557074 604658 557106 604894
rect 557342 604658 557426 604894
rect 557662 604658 557694 604894
rect 557074 604574 557694 604658
rect 557074 604338 557106 604574
rect 557342 604338 557426 604574
rect 557662 604338 557694 604574
rect 557074 568894 557694 604338
rect 557074 568658 557106 568894
rect 557342 568658 557426 568894
rect 557662 568658 557694 568894
rect 557074 568574 557694 568658
rect 557074 568338 557106 568574
rect 557342 568338 557426 568574
rect 557662 568338 557694 568574
rect 557074 532894 557694 568338
rect 557074 532658 557106 532894
rect 557342 532658 557426 532894
rect 557662 532658 557694 532894
rect 557074 532574 557694 532658
rect 557074 532338 557106 532574
rect 557342 532338 557426 532574
rect 557662 532338 557694 532574
rect 557074 496894 557694 532338
rect 557074 496658 557106 496894
rect 557342 496658 557426 496894
rect 557662 496658 557694 496894
rect 557074 496574 557694 496658
rect 557074 496338 557106 496574
rect 557342 496338 557426 496574
rect 557662 496338 557694 496574
rect 557074 460894 557694 496338
rect 557074 460658 557106 460894
rect 557342 460658 557426 460894
rect 557662 460658 557694 460894
rect 557074 460574 557694 460658
rect 557074 460338 557106 460574
rect 557342 460338 557426 460574
rect 557662 460338 557694 460574
rect 557074 424894 557694 460338
rect 557074 424658 557106 424894
rect 557342 424658 557426 424894
rect 557662 424658 557694 424894
rect 557074 424574 557694 424658
rect 557074 424338 557106 424574
rect 557342 424338 557426 424574
rect 557662 424338 557694 424574
rect 557074 388894 557694 424338
rect 557074 388658 557106 388894
rect 557342 388658 557426 388894
rect 557662 388658 557694 388894
rect 557074 388574 557694 388658
rect 557074 388338 557106 388574
rect 557342 388338 557426 388574
rect 557662 388338 557694 388574
rect 557074 352894 557694 388338
rect 557074 352658 557106 352894
rect 557342 352658 557426 352894
rect 557662 352658 557694 352894
rect 557074 352574 557694 352658
rect 557074 352338 557106 352574
rect 557342 352338 557426 352574
rect 557662 352338 557694 352574
rect 557074 316894 557694 352338
rect 557074 316658 557106 316894
rect 557342 316658 557426 316894
rect 557662 316658 557694 316894
rect 557074 316574 557694 316658
rect 557074 316338 557106 316574
rect 557342 316338 557426 316574
rect 557662 316338 557694 316574
rect 557074 280894 557694 316338
rect 557074 280658 557106 280894
rect 557342 280658 557426 280894
rect 557662 280658 557694 280894
rect 557074 280574 557694 280658
rect 557074 280338 557106 280574
rect 557342 280338 557426 280574
rect 557662 280338 557694 280574
rect 557074 244894 557694 280338
rect 557074 244658 557106 244894
rect 557342 244658 557426 244894
rect 557662 244658 557694 244894
rect 557074 244574 557694 244658
rect 557074 244338 557106 244574
rect 557342 244338 557426 244574
rect 557662 244338 557694 244574
rect 557074 208894 557694 244338
rect 557074 208658 557106 208894
rect 557342 208658 557426 208894
rect 557662 208658 557694 208894
rect 557074 208574 557694 208658
rect 557074 208338 557106 208574
rect 557342 208338 557426 208574
rect 557662 208338 557694 208574
rect 557074 172894 557694 208338
rect 557074 172658 557106 172894
rect 557342 172658 557426 172894
rect 557662 172658 557694 172894
rect 557074 172574 557694 172658
rect 557074 172338 557106 172574
rect 557342 172338 557426 172574
rect 557662 172338 557694 172574
rect 557074 136894 557694 172338
rect 557074 136658 557106 136894
rect 557342 136658 557426 136894
rect 557662 136658 557694 136894
rect 557074 136574 557694 136658
rect 557074 136338 557106 136574
rect 557342 136338 557426 136574
rect 557662 136338 557694 136574
rect 557074 100894 557694 136338
rect 557074 100658 557106 100894
rect 557342 100658 557426 100894
rect 557662 100658 557694 100894
rect 557074 100574 557694 100658
rect 557074 100338 557106 100574
rect 557342 100338 557426 100574
rect 557662 100338 557694 100574
rect 557074 64894 557694 100338
rect 557074 64658 557106 64894
rect 557342 64658 557426 64894
rect 557662 64658 557694 64894
rect 557074 64574 557694 64658
rect 557074 64338 557106 64574
rect 557342 64338 557426 64574
rect 557662 64338 557694 64574
rect 557074 28894 557694 64338
rect 557074 28658 557106 28894
rect 557342 28658 557426 28894
rect 557662 28658 557694 28894
rect 557074 28574 557694 28658
rect 557074 28338 557106 28574
rect 557342 28338 557426 28574
rect 557662 28338 557694 28574
rect 557074 -5146 557694 28338
rect 558474 706758 559094 707750
rect 558474 706522 558506 706758
rect 558742 706522 558826 706758
rect 559062 706522 559094 706758
rect 558474 706438 559094 706522
rect 558474 706202 558506 706438
rect 558742 706202 558826 706438
rect 559062 706202 559094 706438
rect 558474 691174 559094 706202
rect 558474 690938 558506 691174
rect 558742 690938 558826 691174
rect 559062 690938 559094 691174
rect 558474 690854 559094 690938
rect 558474 690618 558506 690854
rect 558742 690618 558826 690854
rect 559062 690618 559094 690854
rect 558474 655174 559094 690618
rect 558474 654938 558506 655174
rect 558742 654938 558826 655174
rect 559062 654938 559094 655174
rect 558474 654854 559094 654938
rect 558474 654618 558506 654854
rect 558742 654618 558826 654854
rect 559062 654618 559094 654854
rect 558474 619174 559094 654618
rect 558474 618938 558506 619174
rect 558742 618938 558826 619174
rect 559062 618938 559094 619174
rect 558474 618854 559094 618938
rect 558474 618618 558506 618854
rect 558742 618618 558826 618854
rect 559062 618618 559094 618854
rect 558474 583174 559094 618618
rect 558474 582938 558506 583174
rect 558742 582938 558826 583174
rect 559062 582938 559094 583174
rect 558474 582854 559094 582938
rect 558474 582618 558506 582854
rect 558742 582618 558826 582854
rect 559062 582618 559094 582854
rect 558474 547174 559094 582618
rect 558474 546938 558506 547174
rect 558742 546938 558826 547174
rect 559062 546938 559094 547174
rect 558474 546854 559094 546938
rect 558474 546618 558506 546854
rect 558742 546618 558826 546854
rect 559062 546618 559094 546854
rect 558474 511174 559094 546618
rect 558474 510938 558506 511174
rect 558742 510938 558826 511174
rect 559062 510938 559094 511174
rect 558474 510854 559094 510938
rect 558474 510618 558506 510854
rect 558742 510618 558826 510854
rect 559062 510618 559094 510854
rect 558474 475174 559094 510618
rect 558474 474938 558506 475174
rect 558742 474938 558826 475174
rect 559062 474938 559094 475174
rect 558474 474854 559094 474938
rect 558474 474618 558506 474854
rect 558742 474618 558826 474854
rect 559062 474618 559094 474854
rect 558474 439174 559094 474618
rect 558474 438938 558506 439174
rect 558742 438938 558826 439174
rect 559062 438938 559094 439174
rect 558474 438854 559094 438938
rect 558474 438618 558506 438854
rect 558742 438618 558826 438854
rect 559062 438618 559094 438854
rect 558474 403174 559094 438618
rect 558474 402938 558506 403174
rect 558742 402938 558826 403174
rect 559062 402938 559094 403174
rect 558474 402854 559094 402938
rect 558474 402618 558506 402854
rect 558742 402618 558826 402854
rect 559062 402618 559094 402854
rect 558474 367174 559094 402618
rect 558474 366938 558506 367174
rect 558742 366938 558826 367174
rect 559062 366938 559094 367174
rect 558474 366854 559094 366938
rect 558474 366618 558506 366854
rect 558742 366618 558826 366854
rect 559062 366618 559094 366854
rect 558474 331174 559094 366618
rect 558474 330938 558506 331174
rect 558742 330938 558826 331174
rect 559062 330938 559094 331174
rect 558474 330854 559094 330938
rect 558474 330618 558506 330854
rect 558742 330618 558826 330854
rect 559062 330618 559094 330854
rect 558474 295174 559094 330618
rect 558474 294938 558506 295174
rect 558742 294938 558826 295174
rect 559062 294938 559094 295174
rect 558474 294854 559094 294938
rect 558474 294618 558506 294854
rect 558742 294618 558826 294854
rect 559062 294618 559094 294854
rect 558474 259174 559094 294618
rect 558474 258938 558506 259174
rect 558742 258938 558826 259174
rect 559062 258938 559094 259174
rect 558474 258854 559094 258938
rect 558474 258618 558506 258854
rect 558742 258618 558826 258854
rect 559062 258618 559094 258854
rect 558474 223174 559094 258618
rect 558474 222938 558506 223174
rect 558742 222938 558826 223174
rect 559062 222938 559094 223174
rect 558474 222854 559094 222938
rect 558474 222618 558506 222854
rect 558742 222618 558826 222854
rect 559062 222618 559094 222854
rect 558474 187174 559094 222618
rect 558474 186938 558506 187174
rect 558742 186938 558826 187174
rect 559062 186938 559094 187174
rect 558474 186854 559094 186938
rect 558474 186618 558506 186854
rect 558742 186618 558826 186854
rect 559062 186618 559094 186854
rect 558474 151174 559094 186618
rect 558474 150938 558506 151174
rect 558742 150938 558826 151174
rect 559062 150938 559094 151174
rect 558474 150854 559094 150938
rect 558474 150618 558506 150854
rect 558742 150618 558826 150854
rect 559062 150618 559094 150854
rect 558474 115174 559094 150618
rect 558474 114938 558506 115174
rect 558742 114938 558826 115174
rect 559062 114938 559094 115174
rect 558474 114854 559094 114938
rect 558474 114618 558506 114854
rect 558742 114618 558826 114854
rect 559062 114618 559094 114854
rect 558474 79174 559094 114618
rect 558474 78938 558506 79174
rect 558742 78938 558826 79174
rect 559062 78938 559094 79174
rect 558474 78854 559094 78938
rect 558474 78618 558506 78854
rect 558742 78618 558826 78854
rect 559062 78618 559094 78854
rect 558474 43174 559094 78618
rect 558474 42938 558506 43174
rect 558742 42938 558826 43174
rect 559062 42938 559094 43174
rect 558474 42854 559094 42938
rect 558474 42618 558506 42854
rect 558742 42618 558826 42854
rect 559062 42618 559094 42854
rect 558474 7174 559094 42618
rect 558474 6938 558506 7174
rect 558742 6938 558826 7174
rect 559062 6938 559094 7174
rect 558474 6854 559094 6938
rect 558474 6618 558506 6854
rect 558742 6618 558826 6854
rect 559062 6618 559094 6854
rect 558474 -2266 559094 6618
rect 559874 705798 560494 705830
rect 559874 705562 559906 705798
rect 560142 705562 560226 705798
rect 560462 705562 560494 705798
rect 559874 705478 560494 705562
rect 559874 705242 559906 705478
rect 560142 705242 560226 705478
rect 560462 705242 560494 705478
rect 559874 669454 560494 705242
rect 559874 669218 559906 669454
rect 560142 669218 560226 669454
rect 560462 669218 560494 669454
rect 559874 669134 560494 669218
rect 559874 668898 559906 669134
rect 560142 668898 560226 669134
rect 560462 668898 560494 669134
rect 559874 633454 560494 668898
rect 559874 633218 559906 633454
rect 560142 633218 560226 633454
rect 560462 633218 560494 633454
rect 559874 633134 560494 633218
rect 559874 632898 559906 633134
rect 560142 632898 560226 633134
rect 560462 632898 560494 633134
rect 559874 597454 560494 632898
rect 559874 597218 559906 597454
rect 560142 597218 560226 597454
rect 560462 597218 560494 597454
rect 559874 597134 560494 597218
rect 559874 596898 559906 597134
rect 560142 596898 560226 597134
rect 560462 596898 560494 597134
rect 559874 561454 560494 596898
rect 559874 561218 559906 561454
rect 560142 561218 560226 561454
rect 560462 561218 560494 561454
rect 559874 561134 560494 561218
rect 559874 560898 559906 561134
rect 560142 560898 560226 561134
rect 560462 560898 560494 561134
rect 559874 525454 560494 560898
rect 559874 525218 559906 525454
rect 560142 525218 560226 525454
rect 560462 525218 560494 525454
rect 559874 525134 560494 525218
rect 559874 524898 559906 525134
rect 560142 524898 560226 525134
rect 560462 524898 560494 525134
rect 559874 489454 560494 524898
rect 559874 489218 559906 489454
rect 560142 489218 560226 489454
rect 560462 489218 560494 489454
rect 559874 489134 560494 489218
rect 559874 488898 559906 489134
rect 560142 488898 560226 489134
rect 560462 488898 560494 489134
rect 559874 453454 560494 488898
rect 559874 453218 559906 453454
rect 560142 453218 560226 453454
rect 560462 453218 560494 453454
rect 559874 453134 560494 453218
rect 559874 452898 559906 453134
rect 560142 452898 560226 453134
rect 560462 452898 560494 453134
rect 559874 417454 560494 452898
rect 559874 417218 559906 417454
rect 560142 417218 560226 417454
rect 560462 417218 560494 417454
rect 559874 417134 560494 417218
rect 559874 416898 559906 417134
rect 560142 416898 560226 417134
rect 560462 416898 560494 417134
rect 559874 381454 560494 416898
rect 559874 381218 559906 381454
rect 560142 381218 560226 381454
rect 560462 381218 560494 381454
rect 559874 381134 560494 381218
rect 559874 380898 559906 381134
rect 560142 380898 560226 381134
rect 560462 380898 560494 381134
rect 559874 345454 560494 380898
rect 559874 345218 559906 345454
rect 560142 345218 560226 345454
rect 560462 345218 560494 345454
rect 559874 345134 560494 345218
rect 559874 344898 559906 345134
rect 560142 344898 560226 345134
rect 560462 344898 560494 345134
rect 559874 309454 560494 344898
rect 559874 309218 559906 309454
rect 560142 309218 560226 309454
rect 560462 309218 560494 309454
rect 559874 309134 560494 309218
rect 559874 308898 559906 309134
rect 560142 308898 560226 309134
rect 560462 308898 560494 309134
rect 559874 273454 560494 308898
rect 559874 273218 559906 273454
rect 560142 273218 560226 273454
rect 560462 273218 560494 273454
rect 559874 273134 560494 273218
rect 559874 272898 559906 273134
rect 560142 272898 560226 273134
rect 560462 272898 560494 273134
rect 559874 237454 560494 272898
rect 559874 237218 559906 237454
rect 560142 237218 560226 237454
rect 560462 237218 560494 237454
rect 559874 237134 560494 237218
rect 559874 236898 559906 237134
rect 560142 236898 560226 237134
rect 560462 236898 560494 237134
rect 559874 201454 560494 236898
rect 559874 201218 559906 201454
rect 560142 201218 560226 201454
rect 560462 201218 560494 201454
rect 559874 201134 560494 201218
rect 559874 200898 559906 201134
rect 560142 200898 560226 201134
rect 560462 200898 560494 201134
rect 559874 165454 560494 200898
rect 559874 165218 559906 165454
rect 560142 165218 560226 165454
rect 560462 165218 560494 165454
rect 559874 165134 560494 165218
rect 559874 164898 559906 165134
rect 560142 164898 560226 165134
rect 560462 164898 560494 165134
rect 559874 129454 560494 164898
rect 559874 129218 559906 129454
rect 560142 129218 560226 129454
rect 560462 129218 560494 129454
rect 559874 129134 560494 129218
rect 559874 128898 559906 129134
rect 560142 128898 560226 129134
rect 560462 128898 560494 129134
rect 559874 93454 560494 128898
rect 559874 93218 559906 93454
rect 560142 93218 560226 93454
rect 560462 93218 560494 93454
rect 559874 93134 560494 93218
rect 559874 92898 559906 93134
rect 560142 92898 560226 93134
rect 560462 92898 560494 93134
rect 559874 57454 560494 92898
rect 559874 57218 559906 57454
rect 560142 57218 560226 57454
rect 560462 57218 560494 57454
rect 559874 57134 560494 57218
rect 559874 56898 559906 57134
rect 560142 56898 560226 57134
rect 560462 56898 560494 57134
rect 559874 21454 560494 56898
rect 559874 21218 559906 21454
rect 560142 21218 560226 21454
rect 560462 21218 560494 21454
rect 559874 21134 560494 21218
rect 559874 20898 559906 21134
rect 560142 20898 560226 21134
rect 560462 20898 560494 21134
rect 559874 -1306 560494 20898
rect 559874 -1542 559906 -1306
rect 560142 -1542 560226 -1306
rect 560462 -1542 560494 -1306
rect 559874 -1626 560494 -1542
rect 559874 -1862 559906 -1626
rect 560142 -1862 560226 -1626
rect 560462 -1862 560494 -1626
rect 559874 -1894 560494 -1862
rect 560794 680614 561414 711002
rect 565914 710598 566534 711590
rect 565914 710362 565946 710598
rect 566182 710362 566266 710598
rect 566502 710362 566534 710598
rect 565914 710278 566534 710362
rect 565914 710042 565946 710278
rect 566182 710042 566266 710278
rect 566502 710042 566534 710278
rect 560794 680378 560826 680614
rect 561062 680378 561146 680614
rect 561382 680378 561414 680614
rect 560794 680294 561414 680378
rect 560794 680058 560826 680294
rect 561062 680058 561146 680294
rect 561382 680058 561414 680294
rect 560794 644614 561414 680058
rect 560794 644378 560826 644614
rect 561062 644378 561146 644614
rect 561382 644378 561414 644614
rect 560794 644294 561414 644378
rect 560794 644058 560826 644294
rect 561062 644058 561146 644294
rect 561382 644058 561414 644294
rect 560794 608614 561414 644058
rect 560794 608378 560826 608614
rect 561062 608378 561146 608614
rect 561382 608378 561414 608614
rect 560794 608294 561414 608378
rect 560794 608058 560826 608294
rect 561062 608058 561146 608294
rect 561382 608058 561414 608294
rect 560794 572614 561414 608058
rect 560794 572378 560826 572614
rect 561062 572378 561146 572614
rect 561382 572378 561414 572614
rect 560794 572294 561414 572378
rect 560794 572058 560826 572294
rect 561062 572058 561146 572294
rect 561382 572058 561414 572294
rect 560794 536614 561414 572058
rect 560794 536378 560826 536614
rect 561062 536378 561146 536614
rect 561382 536378 561414 536614
rect 560794 536294 561414 536378
rect 560794 536058 560826 536294
rect 561062 536058 561146 536294
rect 561382 536058 561414 536294
rect 560794 500614 561414 536058
rect 560794 500378 560826 500614
rect 561062 500378 561146 500614
rect 561382 500378 561414 500614
rect 560794 500294 561414 500378
rect 560794 500058 560826 500294
rect 561062 500058 561146 500294
rect 561382 500058 561414 500294
rect 560794 464614 561414 500058
rect 560794 464378 560826 464614
rect 561062 464378 561146 464614
rect 561382 464378 561414 464614
rect 560794 464294 561414 464378
rect 560794 464058 560826 464294
rect 561062 464058 561146 464294
rect 561382 464058 561414 464294
rect 560794 428614 561414 464058
rect 560794 428378 560826 428614
rect 561062 428378 561146 428614
rect 561382 428378 561414 428614
rect 560794 428294 561414 428378
rect 560794 428058 560826 428294
rect 561062 428058 561146 428294
rect 561382 428058 561414 428294
rect 560794 392614 561414 428058
rect 560794 392378 560826 392614
rect 561062 392378 561146 392614
rect 561382 392378 561414 392614
rect 560794 392294 561414 392378
rect 560794 392058 560826 392294
rect 561062 392058 561146 392294
rect 561382 392058 561414 392294
rect 560794 356614 561414 392058
rect 560794 356378 560826 356614
rect 561062 356378 561146 356614
rect 561382 356378 561414 356614
rect 560794 356294 561414 356378
rect 560794 356058 560826 356294
rect 561062 356058 561146 356294
rect 561382 356058 561414 356294
rect 560794 320614 561414 356058
rect 560794 320378 560826 320614
rect 561062 320378 561146 320614
rect 561382 320378 561414 320614
rect 560794 320294 561414 320378
rect 560794 320058 560826 320294
rect 561062 320058 561146 320294
rect 561382 320058 561414 320294
rect 560794 284614 561414 320058
rect 560794 284378 560826 284614
rect 561062 284378 561146 284614
rect 561382 284378 561414 284614
rect 560794 284294 561414 284378
rect 560794 284058 560826 284294
rect 561062 284058 561146 284294
rect 561382 284058 561414 284294
rect 560794 248614 561414 284058
rect 560794 248378 560826 248614
rect 561062 248378 561146 248614
rect 561382 248378 561414 248614
rect 560794 248294 561414 248378
rect 560794 248058 560826 248294
rect 561062 248058 561146 248294
rect 561382 248058 561414 248294
rect 560794 212614 561414 248058
rect 560794 212378 560826 212614
rect 561062 212378 561146 212614
rect 561382 212378 561414 212614
rect 560794 212294 561414 212378
rect 560794 212058 560826 212294
rect 561062 212058 561146 212294
rect 561382 212058 561414 212294
rect 560794 176614 561414 212058
rect 560794 176378 560826 176614
rect 561062 176378 561146 176614
rect 561382 176378 561414 176614
rect 560794 176294 561414 176378
rect 560794 176058 560826 176294
rect 561062 176058 561146 176294
rect 561382 176058 561414 176294
rect 560794 140614 561414 176058
rect 560794 140378 560826 140614
rect 561062 140378 561146 140614
rect 561382 140378 561414 140614
rect 560794 140294 561414 140378
rect 560794 140058 560826 140294
rect 561062 140058 561146 140294
rect 561382 140058 561414 140294
rect 560794 104614 561414 140058
rect 560794 104378 560826 104614
rect 561062 104378 561146 104614
rect 561382 104378 561414 104614
rect 560794 104294 561414 104378
rect 560794 104058 560826 104294
rect 561062 104058 561146 104294
rect 561382 104058 561414 104294
rect 560794 68614 561414 104058
rect 560794 68378 560826 68614
rect 561062 68378 561146 68614
rect 561382 68378 561414 68614
rect 560794 68294 561414 68378
rect 560794 68058 560826 68294
rect 561062 68058 561146 68294
rect 561382 68058 561414 68294
rect 560794 32614 561414 68058
rect 560794 32378 560826 32614
rect 561062 32378 561146 32614
rect 561382 32378 561414 32614
rect 560794 32294 561414 32378
rect 560794 32058 560826 32294
rect 561062 32058 561146 32294
rect 561382 32058 561414 32294
rect 558474 -2502 558506 -2266
rect 558742 -2502 558826 -2266
rect 559062 -2502 559094 -2266
rect 558474 -2586 559094 -2502
rect 558474 -2822 558506 -2586
rect 558742 -2822 558826 -2586
rect 559062 -2822 559094 -2586
rect 558474 -3814 559094 -2822
rect 557074 -5382 557106 -5146
rect 557342 -5382 557426 -5146
rect 557662 -5382 557694 -5146
rect 557074 -5466 557694 -5382
rect 557074 -5702 557106 -5466
rect 557342 -5702 557426 -5466
rect 557662 -5702 557694 -5466
rect 557074 -5734 557694 -5702
rect 555674 -6342 555706 -6106
rect 555942 -6342 556026 -6106
rect 556262 -6342 556294 -6106
rect 555674 -6426 556294 -6342
rect 555674 -6662 555706 -6426
rect 555942 -6662 556026 -6426
rect 556262 -6662 556294 -6426
rect 555674 -7654 556294 -6662
rect 560794 -7066 561414 32058
rect 562194 708678 562814 709670
rect 562194 708442 562226 708678
rect 562462 708442 562546 708678
rect 562782 708442 562814 708678
rect 562194 708358 562814 708442
rect 562194 708122 562226 708358
rect 562462 708122 562546 708358
rect 562782 708122 562814 708358
rect 562194 694894 562814 708122
rect 562194 694658 562226 694894
rect 562462 694658 562546 694894
rect 562782 694658 562814 694894
rect 562194 694574 562814 694658
rect 562194 694338 562226 694574
rect 562462 694338 562546 694574
rect 562782 694338 562814 694574
rect 562194 658894 562814 694338
rect 562194 658658 562226 658894
rect 562462 658658 562546 658894
rect 562782 658658 562814 658894
rect 562194 658574 562814 658658
rect 562194 658338 562226 658574
rect 562462 658338 562546 658574
rect 562782 658338 562814 658574
rect 562194 622894 562814 658338
rect 562194 622658 562226 622894
rect 562462 622658 562546 622894
rect 562782 622658 562814 622894
rect 562194 622574 562814 622658
rect 562194 622338 562226 622574
rect 562462 622338 562546 622574
rect 562782 622338 562814 622574
rect 562194 586894 562814 622338
rect 562194 586658 562226 586894
rect 562462 586658 562546 586894
rect 562782 586658 562814 586894
rect 562194 586574 562814 586658
rect 562194 586338 562226 586574
rect 562462 586338 562546 586574
rect 562782 586338 562814 586574
rect 562194 550894 562814 586338
rect 562194 550658 562226 550894
rect 562462 550658 562546 550894
rect 562782 550658 562814 550894
rect 562194 550574 562814 550658
rect 562194 550338 562226 550574
rect 562462 550338 562546 550574
rect 562782 550338 562814 550574
rect 562194 514894 562814 550338
rect 562194 514658 562226 514894
rect 562462 514658 562546 514894
rect 562782 514658 562814 514894
rect 562194 514574 562814 514658
rect 562194 514338 562226 514574
rect 562462 514338 562546 514574
rect 562782 514338 562814 514574
rect 562194 478894 562814 514338
rect 562194 478658 562226 478894
rect 562462 478658 562546 478894
rect 562782 478658 562814 478894
rect 562194 478574 562814 478658
rect 562194 478338 562226 478574
rect 562462 478338 562546 478574
rect 562782 478338 562814 478574
rect 562194 442894 562814 478338
rect 562194 442658 562226 442894
rect 562462 442658 562546 442894
rect 562782 442658 562814 442894
rect 562194 442574 562814 442658
rect 562194 442338 562226 442574
rect 562462 442338 562546 442574
rect 562782 442338 562814 442574
rect 562194 406894 562814 442338
rect 562194 406658 562226 406894
rect 562462 406658 562546 406894
rect 562782 406658 562814 406894
rect 562194 406574 562814 406658
rect 562194 406338 562226 406574
rect 562462 406338 562546 406574
rect 562782 406338 562814 406574
rect 562194 370894 562814 406338
rect 562194 370658 562226 370894
rect 562462 370658 562546 370894
rect 562782 370658 562814 370894
rect 562194 370574 562814 370658
rect 562194 370338 562226 370574
rect 562462 370338 562546 370574
rect 562782 370338 562814 370574
rect 562194 334894 562814 370338
rect 562194 334658 562226 334894
rect 562462 334658 562546 334894
rect 562782 334658 562814 334894
rect 562194 334574 562814 334658
rect 562194 334338 562226 334574
rect 562462 334338 562546 334574
rect 562782 334338 562814 334574
rect 562194 298894 562814 334338
rect 562194 298658 562226 298894
rect 562462 298658 562546 298894
rect 562782 298658 562814 298894
rect 562194 298574 562814 298658
rect 562194 298338 562226 298574
rect 562462 298338 562546 298574
rect 562782 298338 562814 298574
rect 562194 262894 562814 298338
rect 562194 262658 562226 262894
rect 562462 262658 562546 262894
rect 562782 262658 562814 262894
rect 562194 262574 562814 262658
rect 562194 262338 562226 262574
rect 562462 262338 562546 262574
rect 562782 262338 562814 262574
rect 562194 226894 562814 262338
rect 562194 226658 562226 226894
rect 562462 226658 562546 226894
rect 562782 226658 562814 226894
rect 562194 226574 562814 226658
rect 562194 226338 562226 226574
rect 562462 226338 562546 226574
rect 562782 226338 562814 226574
rect 562194 190894 562814 226338
rect 562194 190658 562226 190894
rect 562462 190658 562546 190894
rect 562782 190658 562814 190894
rect 562194 190574 562814 190658
rect 562194 190338 562226 190574
rect 562462 190338 562546 190574
rect 562782 190338 562814 190574
rect 562194 154894 562814 190338
rect 562194 154658 562226 154894
rect 562462 154658 562546 154894
rect 562782 154658 562814 154894
rect 562194 154574 562814 154658
rect 562194 154338 562226 154574
rect 562462 154338 562546 154574
rect 562782 154338 562814 154574
rect 562194 118894 562814 154338
rect 562194 118658 562226 118894
rect 562462 118658 562546 118894
rect 562782 118658 562814 118894
rect 562194 118574 562814 118658
rect 562194 118338 562226 118574
rect 562462 118338 562546 118574
rect 562782 118338 562814 118574
rect 562194 82894 562814 118338
rect 562194 82658 562226 82894
rect 562462 82658 562546 82894
rect 562782 82658 562814 82894
rect 562194 82574 562814 82658
rect 562194 82338 562226 82574
rect 562462 82338 562546 82574
rect 562782 82338 562814 82574
rect 562194 46894 562814 82338
rect 562194 46658 562226 46894
rect 562462 46658 562546 46894
rect 562782 46658 562814 46894
rect 562194 46574 562814 46658
rect 562194 46338 562226 46574
rect 562462 46338 562546 46574
rect 562782 46338 562814 46574
rect 562194 10894 562814 46338
rect 562194 10658 562226 10894
rect 562462 10658 562546 10894
rect 562782 10658 562814 10894
rect 562194 10574 562814 10658
rect 562194 10338 562226 10574
rect 562462 10338 562546 10574
rect 562782 10338 562814 10574
rect 562194 -4186 562814 10338
rect 563594 707718 564214 707750
rect 563594 707482 563626 707718
rect 563862 707482 563946 707718
rect 564182 707482 564214 707718
rect 563594 707398 564214 707482
rect 563594 707162 563626 707398
rect 563862 707162 563946 707398
rect 564182 707162 564214 707398
rect 563594 673174 564214 707162
rect 563594 672938 563626 673174
rect 563862 672938 563946 673174
rect 564182 672938 564214 673174
rect 563594 672854 564214 672938
rect 563594 672618 563626 672854
rect 563862 672618 563946 672854
rect 564182 672618 564214 672854
rect 563594 637174 564214 672618
rect 563594 636938 563626 637174
rect 563862 636938 563946 637174
rect 564182 636938 564214 637174
rect 563594 636854 564214 636938
rect 563594 636618 563626 636854
rect 563862 636618 563946 636854
rect 564182 636618 564214 636854
rect 563594 601174 564214 636618
rect 563594 600938 563626 601174
rect 563862 600938 563946 601174
rect 564182 600938 564214 601174
rect 563594 600854 564214 600938
rect 563594 600618 563626 600854
rect 563862 600618 563946 600854
rect 564182 600618 564214 600854
rect 563594 565174 564214 600618
rect 563594 564938 563626 565174
rect 563862 564938 563946 565174
rect 564182 564938 564214 565174
rect 563594 564854 564214 564938
rect 563594 564618 563626 564854
rect 563862 564618 563946 564854
rect 564182 564618 564214 564854
rect 563594 529174 564214 564618
rect 563594 528938 563626 529174
rect 563862 528938 563946 529174
rect 564182 528938 564214 529174
rect 563594 528854 564214 528938
rect 563594 528618 563626 528854
rect 563862 528618 563946 528854
rect 564182 528618 564214 528854
rect 563594 493174 564214 528618
rect 563594 492938 563626 493174
rect 563862 492938 563946 493174
rect 564182 492938 564214 493174
rect 563594 492854 564214 492938
rect 563594 492618 563626 492854
rect 563862 492618 563946 492854
rect 564182 492618 564214 492854
rect 563594 457174 564214 492618
rect 563594 456938 563626 457174
rect 563862 456938 563946 457174
rect 564182 456938 564214 457174
rect 563594 456854 564214 456938
rect 563594 456618 563626 456854
rect 563862 456618 563946 456854
rect 564182 456618 564214 456854
rect 563594 421174 564214 456618
rect 563594 420938 563626 421174
rect 563862 420938 563946 421174
rect 564182 420938 564214 421174
rect 563594 420854 564214 420938
rect 563594 420618 563626 420854
rect 563862 420618 563946 420854
rect 564182 420618 564214 420854
rect 563594 385174 564214 420618
rect 563594 384938 563626 385174
rect 563862 384938 563946 385174
rect 564182 384938 564214 385174
rect 563594 384854 564214 384938
rect 563594 384618 563626 384854
rect 563862 384618 563946 384854
rect 564182 384618 564214 384854
rect 563594 349174 564214 384618
rect 563594 348938 563626 349174
rect 563862 348938 563946 349174
rect 564182 348938 564214 349174
rect 563594 348854 564214 348938
rect 563594 348618 563626 348854
rect 563862 348618 563946 348854
rect 564182 348618 564214 348854
rect 563594 313174 564214 348618
rect 563594 312938 563626 313174
rect 563862 312938 563946 313174
rect 564182 312938 564214 313174
rect 563594 312854 564214 312938
rect 563594 312618 563626 312854
rect 563862 312618 563946 312854
rect 564182 312618 564214 312854
rect 563594 277174 564214 312618
rect 563594 276938 563626 277174
rect 563862 276938 563946 277174
rect 564182 276938 564214 277174
rect 563594 276854 564214 276938
rect 563594 276618 563626 276854
rect 563862 276618 563946 276854
rect 564182 276618 564214 276854
rect 563594 241174 564214 276618
rect 563594 240938 563626 241174
rect 563862 240938 563946 241174
rect 564182 240938 564214 241174
rect 563594 240854 564214 240938
rect 563594 240618 563626 240854
rect 563862 240618 563946 240854
rect 564182 240618 564214 240854
rect 563594 205174 564214 240618
rect 563594 204938 563626 205174
rect 563862 204938 563946 205174
rect 564182 204938 564214 205174
rect 563594 204854 564214 204938
rect 563594 204618 563626 204854
rect 563862 204618 563946 204854
rect 564182 204618 564214 204854
rect 563594 169174 564214 204618
rect 563594 168938 563626 169174
rect 563862 168938 563946 169174
rect 564182 168938 564214 169174
rect 563594 168854 564214 168938
rect 563594 168618 563626 168854
rect 563862 168618 563946 168854
rect 564182 168618 564214 168854
rect 563594 133174 564214 168618
rect 563594 132938 563626 133174
rect 563862 132938 563946 133174
rect 564182 132938 564214 133174
rect 563594 132854 564214 132938
rect 563594 132618 563626 132854
rect 563862 132618 563946 132854
rect 564182 132618 564214 132854
rect 563594 97174 564214 132618
rect 563594 96938 563626 97174
rect 563862 96938 563946 97174
rect 564182 96938 564214 97174
rect 563594 96854 564214 96938
rect 563594 96618 563626 96854
rect 563862 96618 563946 96854
rect 564182 96618 564214 96854
rect 563594 61174 564214 96618
rect 563594 60938 563626 61174
rect 563862 60938 563946 61174
rect 564182 60938 564214 61174
rect 563594 60854 564214 60938
rect 563594 60618 563626 60854
rect 563862 60618 563946 60854
rect 564182 60618 564214 60854
rect 563594 25174 564214 60618
rect 563594 24938 563626 25174
rect 563862 24938 563946 25174
rect 564182 24938 564214 25174
rect 563594 24854 564214 24938
rect 563594 24618 563626 24854
rect 563862 24618 563946 24854
rect 564182 24618 564214 24854
rect 563594 -3226 564214 24618
rect 564994 704838 565614 705830
rect 564994 704602 565026 704838
rect 565262 704602 565346 704838
rect 565582 704602 565614 704838
rect 564994 704518 565614 704602
rect 564994 704282 565026 704518
rect 565262 704282 565346 704518
rect 565582 704282 565614 704518
rect 564994 687454 565614 704282
rect 564994 687218 565026 687454
rect 565262 687218 565346 687454
rect 565582 687218 565614 687454
rect 564994 687134 565614 687218
rect 564994 686898 565026 687134
rect 565262 686898 565346 687134
rect 565582 686898 565614 687134
rect 564994 651454 565614 686898
rect 564994 651218 565026 651454
rect 565262 651218 565346 651454
rect 565582 651218 565614 651454
rect 564994 651134 565614 651218
rect 564994 650898 565026 651134
rect 565262 650898 565346 651134
rect 565582 650898 565614 651134
rect 564994 615454 565614 650898
rect 564994 615218 565026 615454
rect 565262 615218 565346 615454
rect 565582 615218 565614 615454
rect 564994 615134 565614 615218
rect 564994 614898 565026 615134
rect 565262 614898 565346 615134
rect 565582 614898 565614 615134
rect 564994 579454 565614 614898
rect 564994 579218 565026 579454
rect 565262 579218 565346 579454
rect 565582 579218 565614 579454
rect 564994 579134 565614 579218
rect 564994 578898 565026 579134
rect 565262 578898 565346 579134
rect 565582 578898 565614 579134
rect 564994 543454 565614 578898
rect 564994 543218 565026 543454
rect 565262 543218 565346 543454
rect 565582 543218 565614 543454
rect 564994 543134 565614 543218
rect 564994 542898 565026 543134
rect 565262 542898 565346 543134
rect 565582 542898 565614 543134
rect 564994 507454 565614 542898
rect 564994 507218 565026 507454
rect 565262 507218 565346 507454
rect 565582 507218 565614 507454
rect 564994 507134 565614 507218
rect 564994 506898 565026 507134
rect 565262 506898 565346 507134
rect 565582 506898 565614 507134
rect 564994 471454 565614 506898
rect 564994 471218 565026 471454
rect 565262 471218 565346 471454
rect 565582 471218 565614 471454
rect 564994 471134 565614 471218
rect 564994 470898 565026 471134
rect 565262 470898 565346 471134
rect 565582 470898 565614 471134
rect 564994 435454 565614 470898
rect 564994 435218 565026 435454
rect 565262 435218 565346 435454
rect 565582 435218 565614 435454
rect 564994 435134 565614 435218
rect 564994 434898 565026 435134
rect 565262 434898 565346 435134
rect 565582 434898 565614 435134
rect 564994 399454 565614 434898
rect 564994 399218 565026 399454
rect 565262 399218 565346 399454
rect 565582 399218 565614 399454
rect 564994 399134 565614 399218
rect 564994 398898 565026 399134
rect 565262 398898 565346 399134
rect 565582 398898 565614 399134
rect 564994 363454 565614 398898
rect 564994 363218 565026 363454
rect 565262 363218 565346 363454
rect 565582 363218 565614 363454
rect 564994 363134 565614 363218
rect 564994 362898 565026 363134
rect 565262 362898 565346 363134
rect 565582 362898 565614 363134
rect 564994 327454 565614 362898
rect 564994 327218 565026 327454
rect 565262 327218 565346 327454
rect 565582 327218 565614 327454
rect 564994 327134 565614 327218
rect 564994 326898 565026 327134
rect 565262 326898 565346 327134
rect 565582 326898 565614 327134
rect 564994 291454 565614 326898
rect 564994 291218 565026 291454
rect 565262 291218 565346 291454
rect 565582 291218 565614 291454
rect 564994 291134 565614 291218
rect 564994 290898 565026 291134
rect 565262 290898 565346 291134
rect 565582 290898 565614 291134
rect 564994 255454 565614 290898
rect 564994 255218 565026 255454
rect 565262 255218 565346 255454
rect 565582 255218 565614 255454
rect 564994 255134 565614 255218
rect 564994 254898 565026 255134
rect 565262 254898 565346 255134
rect 565582 254898 565614 255134
rect 564994 219454 565614 254898
rect 564994 219218 565026 219454
rect 565262 219218 565346 219454
rect 565582 219218 565614 219454
rect 564994 219134 565614 219218
rect 564994 218898 565026 219134
rect 565262 218898 565346 219134
rect 565582 218898 565614 219134
rect 564994 183454 565614 218898
rect 564994 183218 565026 183454
rect 565262 183218 565346 183454
rect 565582 183218 565614 183454
rect 564994 183134 565614 183218
rect 564994 182898 565026 183134
rect 565262 182898 565346 183134
rect 565582 182898 565614 183134
rect 564994 147454 565614 182898
rect 564994 147218 565026 147454
rect 565262 147218 565346 147454
rect 565582 147218 565614 147454
rect 564994 147134 565614 147218
rect 564994 146898 565026 147134
rect 565262 146898 565346 147134
rect 565582 146898 565614 147134
rect 564994 111454 565614 146898
rect 564994 111218 565026 111454
rect 565262 111218 565346 111454
rect 565582 111218 565614 111454
rect 564994 111134 565614 111218
rect 564994 110898 565026 111134
rect 565262 110898 565346 111134
rect 565582 110898 565614 111134
rect 564994 75454 565614 110898
rect 564994 75218 565026 75454
rect 565262 75218 565346 75454
rect 565582 75218 565614 75454
rect 564994 75134 565614 75218
rect 564994 74898 565026 75134
rect 565262 74898 565346 75134
rect 565582 74898 565614 75134
rect 564994 39454 565614 74898
rect 564994 39218 565026 39454
rect 565262 39218 565346 39454
rect 565582 39218 565614 39454
rect 564994 39134 565614 39218
rect 564994 38898 565026 39134
rect 565262 38898 565346 39134
rect 565582 38898 565614 39134
rect 564994 3454 565614 38898
rect 564994 3218 565026 3454
rect 565262 3218 565346 3454
rect 565582 3218 565614 3454
rect 564994 3134 565614 3218
rect 564994 2898 565026 3134
rect 565262 2898 565346 3134
rect 565582 2898 565614 3134
rect 564994 -346 565614 2898
rect 564994 -582 565026 -346
rect 565262 -582 565346 -346
rect 565582 -582 565614 -346
rect 564994 -666 565614 -582
rect 564994 -902 565026 -666
rect 565262 -902 565346 -666
rect 565582 -902 565614 -666
rect 564994 -1894 565614 -902
rect 565914 698614 566534 710042
rect 571034 711558 571654 711590
rect 571034 711322 571066 711558
rect 571302 711322 571386 711558
rect 571622 711322 571654 711558
rect 571034 711238 571654 711322
rect 571034 711002 571066 711238
rect 571302 711002 571386 711238
rect 571622 711002 571654 711238
rect 565914 698378 565946 698614
rect 566182 698378 566266 698614
rect 566502 698378 566534 698614
rect 565914 698294 566534 698378
rect 565914 698058 565946 698294
rect 566182 698058 566266 698294
rect 566502 698058 566534 698294
rect 565914 662614 566534 698058
rect 565914 662378 565946 662614
rect 566182 662378 566266 662614
rect 566502 662378 566534 662614
rect 565914 662294 566534 662378
rect 565914 662058 565946 662294
rect 566182 662058 566266 662294
rect 566502 662058 566534 662294
rect 565914 626614 566534 662058
rect 565914 626378 565946 626614
rect 566182 626378 566266 626614
rect 566502 626378 566534 626614
rect 565914 626294 566534 626378
rect 565914 626058 565946 626294
rect 566182 626058 566266 626294
rect 566502 626058 566534 626294
rect 565914 590614 566534 626058
rect 565914 590378 565946 590614
rect 566182 590378 566266 590614
rect 566502 590378 566534 590614
rect 565914 590294 566534 590378
rect 565914 590058 565946 590294
rect 566182 590058 566266 590294
rect 566502 590058 566534 590294
rect 565914 554614 566534 590058
rect 565914 554378 565946 554614
rect 566182 554378 566266 554614
rect 566502 554378 566534 554614
rect 565914 554294 566534 554378
rect 565914 554058 565946 554294
rect 566182 554058 566266 554294
rect 566502 554058 566534 554294
rect 565914 518614 566534 554058
rect 565914 518378 565946 518614
rect 566182 518378 566266 518614
rect 566502 518378 566534 518614
rect 565914 518294 566534 518378
rect 565914 518058 565946 518294
rect 566182 518058 566266 518294
rect 566502 518058 566534 518294
rect 565914 482614 566534 518058
rect 565914 482378 565946 482614
rect 566182 482378 566266 482614
rect 566502 482378 566534 482614
rect 565914 482294 566534 482378
rect 565914 482058 565946 482294
rect 566182 482058 566266 482294
rect 566502 482058 566534 482294
rect 565914 446614 566534 482058
rect 565914 446378 565946 446614
rect 566182 446378 566266 446614
rect 566502 446378 566534 446614
rect 565914 446294 566534 446378
rect 565914 446058 565946 446294
rect 566182 446058 566266 446294
rect 566502 446058 566534 446294
rect 565914 410614 566534 446058
rect 565914 410378 565946 410614
rect 566182 410378 566266 410614
rect 566502 410378 566534 410614
rect 565914 410294 566534 410378
rect 565914 410058 565946 410294
rect 566182 410058 566266 410294
rect 566502 410058 566534 410294
rect 565914 374614 566534 410058
rect 565914 374378 565946 374614
rect 566182 374378 566266 374614
rect 566502 374378 566534 374614
rect 565914 374294 566534 374378
rect 565914 374058 565946 374294
rect 566182 374058 566266 374294
rect 566502 374058 566534 374294
rect 565914 338614 566534 374058
rect 565914 338378 565946 338614
rect 566182 338378 566266 338614
rect 566502 338378 566534 338614
rect 565914 338294 566534 338378
rect 565914 338058 565946 338294
rect 566182 338058 566266 338294
rect 566502 338058 566534 338294
rect 565914 302614 566534 338058
rect 565914 302378 565946 302614
rect 566182 302378 566266 302614
rect 566502 302378 566534 302614
rect 565914 302294 566534 302378
rect 565914 302058 565946 302294
rect 566182 302058 566266 302294
rect 566502 302058 566534 302294
rect 565914 266614 566534 302058
rect 565914 266378 565946 266614
rect 566182 266378 566266 266614
rect 566502 266378 566534 266614
rect 565914 266294 566534 266378
rect 565914 266058 565946 266294
rect 566182 266058 566266 266294
rect 566502 266058 566534 266294
rect 565914 230614 566534 266058
rect 565914 230378 565946 230614
rect 566182 230378 566266 230614
rect 566502 230378 566534 230614
rect 565914 230294 566534 230378
rect 565914 230058 565946 230294
rect 566182 230058 566266 230294
rect 566502 230058 566534 230294
rect 565914 194614 566534 230058
rect 565914 194378 565946 194614
rect 566182 194378 566266 194614
rect 566502 194378 566534 194614
rect 565914 194294 566534 194378
rect 565914 194058 565946 194294
rect 566182 194058 566266 194294
rect 566502 194058 566534 194294
rect 565914 158614 566534 194058
rect 565914 158378 565946 158614
rect 566182 158378 566266 158614
rect 566502 158378 566534 158614
rect 565914 158294 566534 158378
rect 565914 158058 565946 158294
rect 566182 158058 566266 158294
rect 566502 158058 566534 158294
rect 565914 122614 566534 158058
rect 565914 122378 565946 122614
rect 566182 122378 566266 122614
rect 566502 122378 566534 122614
rect 565914 122294 566534 122378
rect 565914 122058 565946 122294
rect 566182 122058 566266 122294
rect 566502 122058 566534 122294
rect 565914 86614 566534 122058
rect 565914 86378 565946 86614
rect 566182 86378 566266 86614
rect 566502 86378 566534 86614
rect 565914 86294 566534 86378
rect 565914 86058 565946 86294
rect 566182 86058 566266 86294
rect 566502 86058 566534 86294
rect 565914 50614 566534 86058
rect 565914 50378 565946 50614
rect 566182 50378 566266 50614
rect 566502 50378 566534 50614
rect 565914 50294 566534 50378
rect 565914 50058 565946 50294
rect 566182 50058 566266 50294
rect 566502 50058 566534 50294
rect 565914 14614 566534 50058
rect 565914 14378 565946 14614
rect 566182 14378 566266 14614
rect 566502 14378 566534 14614
rect 565914 14294 566534 14378
rect 565914 14058 565946 14294
rect 566182 14058 566266 14294
rect 566502 14058 566534 14294
rect 563594 -3462 563626 -3226
rect 563862 -3462 563946 -3226
rect 564182 -3462 564214 -3226
rect 563594 -3546 564214 -3462
rect 563594 -3782 563626 -3546
rect 563862 -3782 563946 -3546
rect 564182 -3782 564214 -3546
rect 563594 -3814 564214 -3782
rect 562194 -4422 562226 -4186
rect 562462 -4422 562546 -4186
rect 562782 -4422 562814 -4186
rect 562194 -4506 562814 -4422
rect 562194 -4742 562226 -4506
rect 562462 -4742 562546 -4506
rect 562782 -4742 562814 -4506
rect 562194 -5734 562814 -4742
rect 560794 -7302 560826 -7066
rect 561062 -7302 561146 -7066
rect 561382 -7302 561414 -7066
rect 560794 -7386 561414 -7302
rect 560794 -7622 560826 -7386
rect 561062 -7622 561146 -7386
rect 561382 -7622 561414 -7386
rect 560794 -7654 561414 -7622
rect 565914 -6106 566534 14058
rect 567314 709638 567934 709670
rect 567314 709402 567346 709638
rect 567582 709402 567666 709638
rect 567902 709402 567934 709638
rect 567314 709318 567934 709402
rect 567314 709082 567346 709318
rect 567582 709082 567666 709318
rect 567902 709082 567934 709318
rect 567314 676894 567934 709082
rect 567314 676658 567346 676894
rect 567582 676658 567666 676894
rect 567902 676658 567934 676894
rect 567314 676574 567934 676658
rect 567314 676338 567346 676574
rect 567582 676338 567666 676574
rect 567902 676338 567934 676574
rect 567314 640894 567934 676338
rect 567314 640658 567346 640894
rect 567582 640658 567666 640894
rect 567902 640658 567934 640894
rect 567314 640574 567934 640658
rect 567314 640338 567346 640574
rect 567582 640338 567666 640574
rect 567902 640338 567934 640574
rect 567314 604894 567934 640338
rect 567314 604658 567346 604894
rect 567582 604658 567666 604894
rect 567902 604658 567934 604894
rect 567314 604574 567934 604658
rect 567314 604338 567346 604574
rect 567582 604338 567666 604574
rect 567902 604338 567934 604574
rect 567314 568894 567934 604338
rect 567314 568658 567346 568894
rect 567582 568658 567666 568894
rect 567902 568658 567934 568894
rect 567314 568574 567934 568658
rect 567314 568338 567346 568574
rect 567582 568338 567666 568574
rect 567902 568338 567934 568574
rect 567314 532894 567934 568338
rect 567314 532658 567346 532894
rect 567582 532658 567666 532894
rect 567902 532658 567934 532894
rect 567314 532574 567934 532658
rect 567314 532338 567346 532574
rect 567582 532338 567666 532574
rect 567902 532338 567934 532574
rect 567314 496894 567934 532338
rect 567314 496658 567346 496894
rect 567582 496658 567666 496894
rect 567902 496658 567934 496894
rect 567314 496574 567934 496658
rect 567314 496338 567346 496574
rect 567582 496338 567666 496574
rect 567902 496338 567934 496574
rect 567314 460894 567934 496338
rect 567314 460658 567346 460894
rect 567582 460658 567666 460894
rect 567902 460658 567934 460894
rect 567314 460574 567934 460658
rect 567314 460338 567346 460574
rect 567582 460338 567666 460574
rect 567902 460338 567934 460574
rect 567314 424894 567934 460338
rect 567314 424658 567346 424894
rect 567582 424658 567666 424894
rect 567902 424658 567934 424894
rect 567314 424574 567934 424658
rect 567314 424338 567346 424574
rect 567582 424338 567666 424574
rect 567902 424338 567934 424574
rect 567314 388894 567934 424338
rect 567314 388658 567346 388894
rect 567582 388658 567666 388894
rect 567902 388658 567934 388894
rect 567314 388574 567934 388658
rect 567314 388338 567346 388574
rect 567582 388338 567666 388574
rect 567902 388338 567934 388574
rect 567314 352894 567934 388338
rect 567314 352658 567346 352894
rect 567582 352658 567666 352894
rect 567902 352658 567934 352894
rect 567314 352574 567934 352658
rect 567314 352338 567346 352574
rect 567582 352338 567666 352574
rect 567902 352338 567934 352574
rect 567314 316894 567934 352338
rect 567314 316658 567346 316894
rect 567582 316658 567666 316894
rect 567902 316658 567934 316894
rect 567314 316574 567934 316658
rect 567314 316338 567346 316574
rect 567582 316338 567666 316574
rect 567902 316338 567934 316574
rect 567314 280894 567934 316338
rect 567314 280658 567346 280894
rect 567582 280658 567666 280894
rect 567902 280658 567934 280894
rect 567314 280574 567934 280658
rect 567314 280338 567346 280574
rect 567582 280338 567666 280574
rect 567902 280338 567934 280574
rect 567314 244894 567934 280338
rect 567314 244658 567346 244894
rect 567582 244658 567666 244894
rect 567902 244658 567934 244894
rect 567314 244574 567934 244658
rect 567314 244338 567346 244574
rect 567582 244338 567666 244574
rect 567902 244338 567934 244574
rect 567314 208894 567934 244338
rect 567314 208658 567346 208894
rect 567582 208658 567666 208894
rect 567902 208658 567934 208894
rect 567314 208574 567934 208658
rect 567314 208338 567346 208574
rect 567582 208338 567666 208574
rect 567902 208338 567934 208574
rect 567314 172894 567934 208338
rect 567314 172658 567346 172894
rect 567582 172658 567666 172894
rect 567902 172658 567934 172894
rect 567314 172574 567934 172658
rect 567314 172338 567346 172574
rect 567582 172338 567666 172574
rect 567902 172338 567934 172574
rect 567314 136894 567934 172338
rect 567314 136658 567346 136894
rect 567582 136658 567666 136894
rect 567902 136658 567934 136894
rect 567314 136574 567934 136658
rect 567314 136338 567346 136574
rect 567582 136338 567666 136574
rect 567902 136338 567934 136574
rect 567314 100894 567934 136338
rect 567314 100658 567346 100894
rect 567582 100658 567666 100894
rect 567902 100658 567934 100894
rect 567314 100574 567934 100658
rect 567314 100338 567346 100574
rect 567582 100338 567666 100574
rect 567902 100338 567934 100574
rect 567314 64894 567934 100338
rect 567314 64658 567346 64894
rect 567582 64658 567666 64894
rect 567902 64658 567934 64894
rect 567314 64574 567934 64658
rect 567314 64338 567346 64574
rect 567582 64338 567666 64574
rect 567902 64338 567934 64574
rect 567314 28894 567934 64338
rect 567314 28658 567346 28894
rect 567582 28658 567666 28894
rect 567902 28658 567934 28894
rect 567314 28574 567934 28658
rect 567314 28338 567346 28574
rect 567582 28338 567666 28574
rect 567902 28338 567934 28574
rect 567314 -5146 567934 28338
rect 568714 706758 569334 707750
rect 568714 706522 568746 706758
rect 568982 706522 569066 706758
rect 569302 706522 569334 706758
rect 568714 706438 569334 706522
rect 568714 706202 568746 706438
rect 568982 706202 569066 706438
rect 569302 706202 569334 706438
rect 568714 691174 569334 706202
rect 568714 690938 568746 691174
rect 568982 690938 569066 691174
rect 569302 690938 569334 691174
rect 568714 690854 569334 690938
rect 568714 690618 568746 690854
rect 568982 690618 569066 690854
rect 569302 690618 569334 690854
rect 568714 655174 569334 690618
rect 568714 654938 568746 655174
rect 568982 654938 569066 655174
rect 569302 654938 569334 655174
rect 568714 654854 569334 654938
rect 568714 654618 568746 654854
rect 568982 654618 569066 654854
rect 569302 654618 569334 654854
rect 568714 619174 569334 654618
rect 568714 618938 568746 619174
rect 568982 618938 569066 619174
rect 569302 618938 569334 619174
rect 568714 618854 569334 618938
rect 568714 618618 568746 618854
rect 568982 618618 569066 618854
rect 569302 618618 569334 618854
rect 568714 583174 569334 618618
rect 568714 582938 568746 583174
rect 568982 582938 569066 583174
rect 569302 582938 569334 583174
rect 568714 582854 569334 582938
rect 568714 582618 568746 582854
rect 568982 582618 569066 582854
rect 569302 582618 569334 582854
rect 568714 547174 569334 582618
rect 568714 546938 568746 547174
rect 568982 546938 569066 547174
rect 569302 546938 569334 547174
rect 568714 546854 569334 546938
rect 568714 546618 568746 546854
rect 568982 546618 569066 546854
rect 569302 546618 569334 546854
rect 568714 511174 569334 546618
rect 568714 510938 568746 511174
rect 568982 510938 569066 511174
rect 569302 510938 569334 511174
rect 568714 510854 569334 510938
rect 568714 510618 568746 510854
rect 568982 510618 569066 510854
rect 569302 510618 569334 510854
rect 568714 475174 569334 510618
rect 568714 474938 568746 475174
rect 568982 474938 569066 475174
rect 569302 474938 569334 475174
rect 568714 474854 569334 474938
rect 568714 474618 568746 474854
rect 568982 474618 569066 474854
rect 569302 474618 569334 474854
rect 568714 439174 569334 474618
rect 568714 438938 568746 439174
rect 568982 438938 569066 439174
rect 569302 438938 569334 439174
rect 568714 438854 569334 438938
rect 568714 438618 568746 438854
rect 568982 438618 569066 438854
rect 569302 438618 569334 438854
rect 568714 403174 569334 438618
rect 568714 402938 568746 403174
rect 568982 402938 569066 403174
rect 569302 402938 569334 403174
rect 568714 402854 569334 402938
rect 568714 402618 568746 402854
rect 568982 402618 569066 402854
rect 569302 402618 569334 402854
rect 568714 367174 569334 402618
rect 568714 366938 568746 367174
rect 568982 366938 569066 367174
rect 569302 366938 569334 367174
rect 568714 366854 569334 366938
rect 568714 366618 568746 366854
rect 568982 366618 569066 366854
rect 569302 366618 569334 366854
rect 568714 331174 569334 366618
rect 568714 330938 568746 331174
rect 568982 330938 569066 331174
rect 569302 330938 569334 331174
rect 568714 330854 569334 330938
rect 568714 330618 568746 330854
rect 568982 330618 569066 330854
rect 569302 330618 569334 330854
rect 568714 295174 569334 330618
rect 568714 294938 568746 295174
rect 568982 294938 569066 295174
rect 569302 294938 569334 295174
rect 568714 294854 569334 294938
rect 568714 294618 568746 294854
rect 568982 294618 569066 294854
rect 569302 294618 569334 294854
rect 568714 259174 569334 294618
rect 568714 258938 568746 259174
rect 568982 258938 569066 259174
rect 569302 258938 569334 259174
rect 568714 258854 569334 258938
rect 568714 258618 568746 258854
rect 568982 258618 569066 258854
rect 569302 258618 569334 258854
rect 568714 223174 569334 258618
rect 568714 222938 568746 223174
rect 568982 222938 569066 223174
rect 569302 222938 569334 223174
rect 568714 222854 569334 222938
rect 568714 222618 568746 222854
rect 568982 222618 569066 222854
rect 569302 222618 569334 222854
rect 568714 187174 569334 222618
rect 568714 186938 568746 187174
rect 568982 186938 569066 187174
rect 569302 186938 569334 187174
rect 568714 186854 569334 186938
rect 568714 186618 568746 186854
rect 568982 186618 569066 186854
rect 569302 186618 569334 186854
rect 568714 151174 569334 186618
rect 568714 150938 568746 151174
rect 568982 150938 569066 151174
rect 569302 150938 569334 151174
rect 568714 150854 569334 150938
rect 568714 150618 568746 150854
rect 568982 150618 569066 150854
rect 569302 150618 569334 150854
rect 568714 115174 569334 150618
rect 568714 114938 568746 115174
rect 568982 114938 569066 115174
rect 569302 114938 569334 115174
rect 568714 114854 569334 114938
rect 568714 114618 568746 114854
rect 568982 114618 569066 114854
rect 569302 114618 569334 114854
rect 568714 79174 569334 114618
rect 568714 78938 568746 79174
rect 568982 78938 569066 79174
rect 569302 78938 569334 79174
rect 568714 78854 569334 78938
rect 568714 78618 568746 78854
rect 568982 78618 569066 78854
rect 569302 78618 569334 78854
rect 568714 43174 569334 78618
rect 568714 42938 568746 43174
rect 568982 42938 569066 43174
rect 569302 42938 569334 43174
rect 568714 42854 569334 42938
rect 568714 42618 568746 42854
rect 568982 42618 569066 42854
rect 569302 42618 569334 42854
rect 568714 7174 569334 42618
rect 568714 6938 568746 7174
rect 568982 6938 569066 7174
rect 569302 6938 569334 7174
rect 568714 6854 569334 6938
rect 568714 6618 568746 6854
rect 568982 6618 569066 6854
rect 569302 6618 569334 6854
rect 568714 -2266 569334 6618
rect 570114 705798 570734 705830
rect 570114 705562 570146 705798
rect 570382 705562 570466 705798
rect 570702 705562 570734 705798
rect 570114 705478 570734 705562
rect 570114 705242 570146 705478
rect 570382 705242 570466 705478
rect 570702 705242 570734 705478
rect 570114 669454 570734 705242
rect 570114 669218 570146 669454
rect 570382 669218 570466 669454
rect 570702 669218 570734 669454
rect 570114 669134 570734 669218
rect 570114 668898 570146 669134
rect 570382 668898 570466 669134
rect 570702 668898 570734 669134
rect 570114 633454 570734 668898
rect 570114 633218 570146 633454
rect 570382 633218 570466 633454
rect 570702 633218 570734 633454
rect 570114 633134 570734 633218
rect 570114 632898 570146 633134
rect 570382 632898 570466 633134
rect 570702 632898 570734 633134
rect 570114 597454 570734 632898
rect 570114 597218 570146 597454
rect 570382 597218 570466 597454
rect 570702 597218 570734 597454
rect 570114 597134 570734 597218
rect 570114 596898 570146 597134
rect 570382 596898 570466 597134
rect 570702 596898 570734 597134
rect 570114 561454 570734 596898
rect 570114 561218 570146 561454
rect 570382 561218 570466 561454
rect 570702 561218 570734 561454
rect 570114 561134 570734 561218
rect 570114 560898 570146 561134
rect 570382 560898 570466 561134
rect 570702 560898 570734 561134
rect 570114 525454 570734 560898
rect 570114 525218 570146 525454
rect 570382 525218 570466 525454
rect 570702 525218 570734 525454
rect 570114 525134 570734 525218
rect 570114 524898 570146 525134
rect 570382 524898 570466 525134
rect 570702 524898 570734 525134
rect 570114 489454 570734 524898
rect 570114 489218 570146 489454
rect 570382 489218 570466 489454
rect 570702 489218 570734 489454
rect 570114 489134 570734 489218
rect 570114 488898 570146 489134
rect 570382 488898 570466 489134
rect 570702 488898 570734 489134
rect 570114 453454 570734 488898
rect 570114 453218 570146 453454
rect 570382 453218 570466 453454
rect 570702 453218 570734 453454
rect 570114 453134 570734 453218
rect 570114 452898 570146 453134
rect 570382 452898 570466 453134
rect 570702 452898 570734 453134
rect 570114 417454 570734 452898
rect 570114 417218 570146 417454
rect 570382 417218 570466 417454
rect 570702 417218 570734 417454
rect 570114 417134 570734 417218
rect 570114 416898 570146 417134
rect 570382 416898 570466 417134
rect 570702 416898 570734 417134
rect 570114 381454 570734 416898
rect 570114 381218 570146 381454
rect 570382 381218 570466 381454
rect 570702 381218 570734 381454
rect 570114 381134 570734 381218
rect 570114 380898 570146 381134
rect 570382 380898 570466 381134
rect 570702 380898 570734 381134
rect 570114 345454 570734 380898
rect 570114 345218 570146 345454
rect 570382 345218 570466 345454
rect 570702 345218 570734 345454
rect 570114 345134 570734 345218
rect 570114 344898 570146 345134
rect 570382 344898 570466 345134
rect 570702 344898 570734 345134
rect 570114 309454 570734 344898
rect 570114 309218 570146 309454
rect 570382 309218 570466 309454
rect 570702 309218 570734 309454
rect 570114 309134 570734 309218
rect 570114 308898 570146 309134
rect 570382 308898 570466 309134
rect 570702 308898 570734 309134
rect 570114 273454 570734 308898
rect 570114 273218 570146 273454
rect 570382 273218 570466 273454
rect 570702 273218 570734 273454
rect 570114 273134 570734 273218
rect 570114 272898 570146 273134
rect 570382 272898 570466 273134
rect 570702 272898 570734 273134
rect 570114 237454 570734 272898
rect 570114 237218 570146 237454
rect 570382 237218 570466 237454
rect 570702 237218 570734 237454
rect 570114 237134 570734 237218
rect 570114 236898 570146 237134
rect 570382 236898 570466 237134
rect 570702 236898 570734 237134
rect 570114 201454 570734 236898
rect 570114 201218 570146 201454
rect 570382 201218 570466 201454
rect 570702 201218 570734 201454
rect 570114 201134 570734 201218
rect 570114 200898 570146 201134
rect 570382 200898 570466 201134
rect 570702 200898 570734 201134
rect 570114 165454 570734 200898
rect 570114 165218 570146 165454
rect 570382 165218 570466 165454
rect 570702 165218 570734 165454
rect 570114 165134 570734 165218
rect 570114 164898 570146 165134
rect 570382 164898 570466 165134
rect 570702 164898 570734 165134
rect 570114 129454 570734 164898
rect 570114 129218 570146 129454
rect 570382 129218 570466 129454
rect 570702 129218 570734 129454
rect 570114 129134 570734 129218
rect 570114 128898 570146 129134
rect 570382 128898 570466 129134
rect 570702 128898 570734 129134
rect 570114 93454 570734 128898
rect 570114 93218 570146 93454
rect 570382 93218 570466 93454
rect 570702 93218 570734 93454
rect 570114 93134 570734 93218
rect 570114 92898 570146 93134
rect 570382 92898 570466 93134
rect 570702 92898 570734 93134
rect 570114 57454 570734 92898
rect 570114 57218 570146 57454
rect 570382 57218 570466 57454
rect 570702 57218 570734 57454
rect 570114 57134 570734 57218
rect 570114 56898 570146 57134
rect 570382 56898 570466 57134
rect 570702 56898 570734 57134
rect 570114 21454 570734 56898
rect 570114 21218 570146 21454
rect 570382 21218 570466 21454
rect 570702 21218 570734 21454
rect 570114 21134 570734 21218
rect 570114 20898 570146 21134
rect 570382 20898 570466 21134
rect 570702 20898 570734 21134
rect 570114 -1306 570734 20898
rect 570114 -1542 570146 -1306
rect 570382 -1542 570466 -1306
rect 570702 -1542 570734 -1306
rect 570114 -1626 570734 -1542
rect 570114 -1862 570146 -1626
rect 570382 -1862 570466 -1626
rect 570702 -1862 570734 -1626
rect 570114 -1894 570734 -1862
rect 571034 680614 571654 711002
rect 576154 710598 576774 711590
rect 576154 710362 576186 710598
rect 576422 710362 576506 710598
rect 576742 710362 576774 710598
rect 576154 710278 576774 710362
rect 576154 710042 576186 710278
rect 576422 710042 576506 710278
rect 576742 710042 576774 710278
rect 571034 680378 571066 680614
rect 571302 680378 571386 680614
rect 571622 680378 571654 680614
rect 571034 680294 571654 680378
rect 571034 680058 571066 680294
rect 571302 680058 571386 680294
rect 571622 680058 571654 680294
rect 571034 644614 571654 680058
rect 571034 644378 571066 644614
rect 571302 644378 571386 644614
rect 571622 644378 571654 644614
rect 571034 644294 571654 644378
rect 571034 644058 571066 644294
rect 571302 644058 571386 644294
rect 571622 644058 571654 644294
rect 571034 608614 571654 644058
rect 571034 608378 571066 608614
rect 571302 608378 571386 608614
rect 571622 608378 571654 608614
rect 571034 608294 571654 608378
rect 571034 608058 571066 608294
rect 571302 608058 571386 608294
rect 571622 608058 571654 608294
rect 571034 572614 571654 608058
rect 571034 572378 571066 572614
rect 571302 572378 571386 572614
rect 571622 572378 571654 572614
rect 571034 572294 571654 572378
rect 571034 572058 571066 572294
rect 571302 572058 571386 572294
rect 571622 572058 571654 572294
rect 571034 536614 571654 572058
rect 571034 536378 571066 536614
rect 571302 536378 571386 536614
rect 571622 536378 571654 536614
rect 571034 536294 571654 536378
rect 571034 536058 571066 536294
rect 571302 536058 571386 536294
rect 571622 536058 571654 536294
rect 571034 500614 571654 536058
rect 571034 500378 571066 500614
rect 571302 500378 571386 500614
rect 571622 500378 571654 500614
rect 571034 500294 571654 500378
rect 571034 500058 571066 500294
rect 571302 500058 571386 500294
rect 571622 500058 571654 500294
rect 571034 464614 571654 500058
rect 571034 464378 571066 464614
rect 571302 464378 571386 464614
rect 571622 464378 571654 464614
rect 571034 464294 571654 464378
rect 571034 464058 571066 464294
rect 571302 464058 571386 464294
rect 571622 464058 571654 464294
rect 571034 428614 571654 464058
rect 571034 428378 571066 428614
rect 571302 428378 571386 428614
rect 571622 428378 571654 428614
rect 571034 428294 571654 428378
rect 571034 428058 571066 428294
rect 571302 428058 571386 428294
rect 571622 428058 571654 428294
rect 571034 392614 571654 428058
rect 571034 392378 571066 392614
rect 571302 392378 571386 392614
rect 571622 392378 571654 392614
rect 571034 392294 571654 392378
rect 571034 392058 571066 392294
rect 571302 392058 571386 392294
rect 571622 392058 571654 392294
rect 571034 356614 571654 392058
rect 571034 356378 571066 356614
rect 571302 356378 571386 356614
rect 571622 356378 571654 356614
rect 571034 356294 571654 356378
rect 571034 356058 571066 356294
rect 571302 356058 571386 356294
rect 571622 356058 571654 356294
rect 571034 320614 571654 356058
rect 571034 320378 571066 320614
rect 571302 320378 571386 320614
rect 571622 320378 571654 320614
rect 571034 320294 571654 320378
rect 571034 320058 571066 320294
rect 571302 320058 571386 320294
rect 571622 320058 571654 320294
rect 571034 284614 571654 320058
rect 571034 284378 571066 284614
rect 571302 284378 571386 284614
rect 571622 284378 571654 284614
rect 571034 284294 571654 284378
rect 571034 284058 571066 284294
rect 571302 284058 571386 284294
rect 571622 284058 571654 284294
rect 571034 248614 571654 284058
rect 571034 248378 571066 248614
rect 571302 248378 571386 248614
rect 571622 248378 571654 248614
rect 571034 248294 571654 248378
rect 571034 248058 571066 248294
rect 571302 248058 571386 248294
rect 571622 248058 571654 248294
rect 571034 212614 571654 248058
rect 571034 212378 571066 212614
rect 571302 212378 571386 212614
rect 571622 212378 571654 212614
rect 571034 212294 571654 212378
rect 571034 212058 571066 212294
rect 571302 212058 571386 212294
rect 571622 212058 571654 212294
rect 571034 176614 571654 212058
rect 571034 176378 571066 176614
rect 571302 176378 571386 176614
rect 571622 176378 571654 176614
rect 571034 176294 571654 176378
rect 571034 176058 571066 176294
rect 571302 176058 571386 176294
rect 571622 176058 571654 176294
rect 571034 140614 571654 176058
rect 571034 140378 571066 140614
rect 571302 140378 571386 140614
rect 571622 140378 571654 140614
rect 571034 140294 571654 140378
rect 571034 140058 571066 140294
rect 571302 140058 571386 140294
rect 571622 140058 571654 140294
rect 571034 104614 571654 140058
rect 571034 104378 571066 104614
rect 571302 104378 571386 104614
rect 571622 104378 571654 104614
rect 571034 104294 571654 104378
rect 571034 104058 571066 104294
rect 571302 104058 571386 104294
rect 571622 104058 571654 104294
rect 571034 68614 571654 104058
rect 571034 68378 571066 68614
rect 571302 68378 571386 68614
rect 571622 68378 571654 68614
rect 571034 68294 571654 68378
rect 571034 68058 571066 68294
rect 571302 68058 571386 68294
rect 571622 68058 571654 68294
rect 571034 32614 571654 68058
rect 571034 32378 571066 32614
rect 571302 32378 571386 32614
rect 571622 32378 571654 32614
rect 571034 32294 571654 32378
rect 571034 32058 571066 32294
rect 571302 32058 571386 32294
rect 571622 32058 571654 32294
rect 568714 -2502 568746 -2266
rect 568982 -2502 569066 -2266
rect 569302 -2502 569334 -2266
rect 568714 -2586 569334 -2502
rect 568714 -2822 568746 -2586
rect 568982 -2822 569066 -2586
rect 569302 -2822 569334 -2586
rect 568714 -3814 569334 -2822
rect 567314 -5382 567346 -5146
rect 567582 -5382 567666 -5146
rect 567902 -5382 567934 -5146
rect 567314 -5466 567934 -5382
rect 567314 -5702 567346 -5466
rect 567582 -5702 567666 -5466
rect 567902 -5702 567934 -5466
rect 567314 -5734 567934 -5702
rect 565914 -6342 565946 -6106
rect 566182 -6342 566266 -6106
rect 566502 -6342 566534 -6106
rect 565914 -6426 566534 -6342
rect 565914 -6662 565946 -6426
rect 566182 -6662 566266 -6426
rect 566502 -6662 566534 -6426
rect 565914 -7654 566534 -6662
rect 571034 -7066 571654 32058
rect 572434 708678 573054 709670
rect 572434 708442 572466 708678
rect 572702 708442 572786 708678
rect 573022 708442 573054 708678
rect 572434 708358 573054 708442
rect 572434 708122 572466 708358
rect 572702 708122 572786 708358
rect 573022 708122 573054 708358
rect 572434 694894 573054 708122
rect 572434 694658 572466 694894
rect 572702 694658 572786 694894
rect 573022 694658 573054 694894
rect 572434 694574 573054 694658
rect 572434 694338 572466 694574
rect 572702 694338 572786 694574
rect 573022 694338 573054 694574
rect 572434 658894 573054 694338
rect 572434 658658 572466 658894
rect 572702 658658 572786 658894
rect 573022 658658 573054 658894
rect 572434 658574 573054 658658
rect 572434 658338 572466 658574
rect 572702 658338 572786 658574
rect 573022 658338 573054 658574
rect 572434 622894 573054 658338
rect 572434 622658 572466 622894
rect 572702 622658 572786 622894
rect 573022 622658 573054 622894
rect 572434 622574 573054 622658
rect 572434 622338 572466 622574
rect 572702 622338 572786 622574
rect 573022 622338 573054 622574
rect 572434 586894 573054 622338
rect 572434 586658 572466 586894
rect 572702 586658 572786 586894
rect 573022 586658 573054 586894
rect 572434 586574 573054 586658
rect 572434 586338 572466 586574
rect 572702 586338 572786 586574
rect 573022 586338 573054 586574
rect 572434 550894 573054 586338
rect 572434 550658 572466 550894
rect 572702 550658 572786 550894
rect 573022 550658 573054 550894
rect 572434 550574 573054 550658
rect 572434 550338 572466 550574
rect 572702 550338 572786 550574
rect 573022 550338 573054 550574
rect 572434 514894 573054 550338
rect 572434 514658 572466 514894
rect 572702 514658 572786 514894
rect 573022 514658 573054 514894
rect 572434 514574 573054 514658
rect 572434 514338 572466 514574
rect 572702 514338 572786 514574
rect 573022 514338 573054 514574
rect 572434 478894 573054 514338
rect 572434 478658 572466 478894
rect 572702 478658 572786 478894
rect 573022 478658 573054 478894
rect 572434 478574 573054 478658
rect 572434 478338 572466 478574
rect 572702 478338 572786 478574
rect 573022 478338 573054 478574
rect 572434 442894 573054 478338
rect 572434 442658 572466 442894
rect 572702 442658 572786 442894
rect 573022 442658 573054 442894
rect 572434 442574 573054 442658
rect 572434 442338 572466 442574
rect 572702 442338 572786 442574
rect 573022 442338 573054 442574
rect 572434 406894 573054 442338
rect 572434 406658 572466 406894
rect 572702 406658 572786 406894
rect 573022 406658 573054 406894
rect 572434 406574 573054 406658
rect 572434 406338 572466 406574
rect 572702 406338 572786 406574
rect 573022 406338 573054 406574
rect 572434 370894 573054 406338
rect 572434 370658 572466 370894
rect 572702 370658 572786 370894
rect 573022 370658 573054 370894
rect 572434 370574 573054 370658
rect 572434 370338 572466 370574
rect 572702 370338 572786 370574
rect 573022 370338 573054 370574
rect 572434 334894 573054 370338
rect 572434 334658 572466 334894
rect 572702 334658 572786 334894
rect 573022 334658 573054 334894
rect 572434 334574 573054 334658
rect 572434 334338 572466 334574
rect 572702 334338 572786 334574
rect 573022 334338 573054 334574
rect 572434 298894 573054 334338
rect 572434 298658 572466 298894
rect 572702 298658 572786 298894
rect 573022 298658 573054 298894
rect 572434 298574 573054 298658
rect 572434 298338 572466 298574
rect 572702 298338 572786 298574
rect 573022 298338 573054 298574
rect 572434 262894 573054 298338
rect 572434 262658 572466 262894
rect 572702 262658 572786 262894
rect 573022 262658 573054 262894
rect 572434 262574 573054 262658
rect 572434 262338 572466 262574
rect 572702 262338 572786 262574
rect 573022 262338 573054 262574
rect 572434 226894 573054 262338
rect 572434 226658 572466 226894
rect 572702 226658 572786 226894
rect 573022 226658 573054 226894
rect 572434 226574 573054 226658
rect 572434 226338 572466 226574
rect 572702 226338 572786 226574
rect 573022 226338 573054 226574
rect 572434 190894 573054 226338
rect 572434 190658 572466 190894
rect 572702 190658 572786 190894
rect 573022 190658 573054 190894
rect 572434 190574 573054 190658
rect 572434 190338 572466 190574
rect 572702 190338 572786 190574
rect 573022 190338 573054 190574
rect 572434 154894 573054 190338
rect 572434 154658 572466 154894
rect 572702 154658 572786 154894
rect 573022 154658 573054 154894
rect 572434 154574 573054 154658
rect 572434 154338 572466 154574
rect 572702 154338 572786 154574
rect 573022 154338 573054 154574
rect 572434 118894 573054 154338
rect 572434 118658 572466 118894
rect 572702 118658 572786 118894
rect 573022 118658 573054 118894
rect 572434 118574 573054 118658
rect 572434 118338 572466 118574
rect 572702 118338 572786 118574
rect 573022 118338 573054 118574
rect 572434 82894 573054 118338
rect 572434 82658 572466 82894
rect 572702 82658 572786 82894
rect 573022 82658 573054 82894
rect 572434 82574 573054 82658
rect 572434 82338 572466 82574
rect 572702 82338 572786 82574
rect 573022 82338 573054 82574
rect 572434 46894 573054 82338
rect 572434 46658 572466 46894
rect 572702 46658 572786 46894
rect 573022 46658 573054 46894
rect 572434 46574 573054 46658
rect 572434 46338 572466 46574
rect 572702 46338 572786 46574
rect 573022 46338 573054 46574
rect 572434 10894 573054 46338
rect 572434 10658 572466 10894
rect 572702 10658 572786 10894
rect 573022 10658 573054 10894
rect 572434 10574 573054 10658
rect 572434 10338 572466 10574
rect 572702 10338 572786 10574
rect 573022 10338 573054 10574
rect 572434 -4186 573054 10338
rect 573834 707718 574454 707750
rect 573834 707482 573866 707718
rect 574102 707482 574186 707718
rect 574422 707482 574454 707718
rect 573834 707398 574454 707482
rect 573834 707162 573866 707398
rect 574102 707162 574186 707398
rect 574422 707162 574454 707398
rect 573834 673174 574454 707162
rect 573834 672938 573866 673174
rect 574102 672938 574186 673174
rect 574422 672938 574454 673174
rect 573834 672854 574454 672938
rect 573834 672618 573866 672854
rect 574102 672618 574186 672854
rect 574422 672618 574454 672854
rect 573834 637174 574454 672618
rect 573834 636938 573866 637174
rect 574102 636938 574186 637174
rect 574422 636938 574454 637174
rect 573834 636854 574454 636938
rect 573834 636618 573866 636854
rect 574102 636618 574186 636854
rect 574422 636618 574454 636854
rect 573834 601174 574454 636618
rect 573834 600938 573866 601174
rect 574102 600938 574186 601174
rect 574422 600938 574454 601174
rect 573834 600854 574454 600938
rect 573834 600618 573866 600854
rect 574102 600618 574186 600854
rect 574422 600618 574454 600854
rect 573834 565174 574454 600618
rect 573834 564938 573866 565174
rect 574102 564938 574186 565174
rect 574422 564938 574454 565174
rect 573834 564854 574454 564938
rect 573834 564618 573866 564854
rect 574102 564618 574186 564854
rect 574422 564618 574454 564854
rect 573834 529174 574454 564618
rect 573834 528938 573866 529174
rect 574102 528938 574186 529174
rect 574422 528938 574454 529174
rect 573834 528854 574454 528938
rect 573834 528618 573866 528854
rect 574102 528618 574186 528854
rect 574422 528618 574454 528854
rect 573834 493174 574454 528618
rect 573834 492938 573866 493174
rect 574102 492938 574186 493174
rect 574422 492938 574454 493174
rect 573834 492854 574454 492938
rect 573834 492618 573866 492854
rect 574102 492618 574186 492854
rect 574422 492618 574454 492854
rect 573834 457174 574454 492618
rect 573834 456938 573866 457174
rect 574102 456938 574186 457174
rect 574422 456938 574454 457174
rect 573834 456854 574454 456938
rect 573834 456618 573866 456854
rect 574102 456618 574186 456854
rect 574422 456618 574454 456854
rect 573834 421174 574454 456618
rect 573834 420938 573866 421174
rect 574102 420938 574186 421174
rect 574422 420938 574454 421174
rect 573834 420854 574454 420938
rect 573834 420618 573866 420854
rect 574102 420618 574186 420854
rect 574422 420618 574454 420854
rect 573834 385174 574454 420618
rect 573834 384938 573866 385174
rect 574102 384938 574186 385174
rect 574422 384938 574454 385174
rect 573834 384854 574454 384938
rect 573834 384618 573866 384854
rect 574102 384618 574186 384854
rect 574422 384618 574454 384854
rect 573834 349174 574454 384618
rect 573834 348938 573866 349174
rect 574102 348938 574186 349174
rect 574422 348938 574454 349174
rect 573834 348854 574454 348938
rect 573834 348618 573866 348854
rect 574102 348618 574186 348854
rect 574422 348618 574454 348854
rect 573834 313174 574454 348618
rect 573834 312938 573866 313174
rect 574102 312938 574186 313174
rect 574422 312938 574454 313174
rect 573834 312854 574454 312938
rect 573834 312618 573866 312854
rect 574102 312618 574186 312854
rect 574422 312618 574454 312854
rect 573834 277174 574454 312618
rect 573834 276938 573866 277174
rect 574102 276938 574186 277174
rect 574422 276938 574454 277174
rect 573834 276854 574454 276938
rect 573834 276618 573866 276854
rect 574102 276618 574186 276854
rect 574422 276618 574454 276854
rect 573834 241174 574454 276618
rect 573834 240938 573866 241174
rect 574102 240938 574186 241174
rect 574422 240938 574454 241174
rect 573834 240854 574454 240938
rect 573834 240618 573866 240854
rect 574102 240618 574186 240854
rect 574422 240618 574454 240854
rect 573834 205174 574454 240618
rect 573834 204938 573866 205174
rect 574102 204938 574186 205174
rect 574422 204938 574454 205174
rect 573834 204854 574454 204938
rect 573834 204618 573866 204854
rect 574102 204618 574186 204854
rect 574422 204618 574454 204854
rect 573834 169174 574454 204618
rect 573834 168938 573866 169174
rect 574102 168938 574186 169174
rect 574422 168938 574454 169174
rect 573834 168854 574454 168938
rect 573834 168618 573866 168854
rect 574102 168618 574186 168854
rect 574422 168618 574454 168854
rect 573834 133174 574454 168618
rect 573834 132938 573866 133174
rect 574102 132938 574186 133174
rect 574422 132938 574454 133174
rect 573834 132854 574454 132938
rect 573834 132618 573866 132854
rect 574102 132618 574186 132854
rect 574422 132618 574454 132854
rect 573834 97174 574454 132618
rect 573834 96938 573866 97174
rect 574102 96938 574186 97174
rect 574422 96938 574454 97174
rect 573834 96854 574454 96938
rect 573834 96618 573866 96854
rect 574102 96618 574186 96854
rect 574422 96618 574454 96854
rect 573834 61174 574454 96618
rect 573834 60938 573866 61174
rect 574102 60938 574186 61174
rect 574422 60938 574454 61174
rect 573834 60854 574454 60938
rect 573834 60618 573866 60854
rect 574102 60618 574186 60854
rect 574422 60618 574454 60854
rect 573834 25174 574454 60618
rect 573834 24938 573866 25174
rect 574102 24938 574186 25174
rect 574422 24938 574454 25174
rect 573834 24854 574454 24938
rect 573834 24618 573866 24854
rect 574102 24618 574186 24854
rect 574422 24618 574454 24854
rect 573834 -3226 574454 24618
rect 575234 704838 575854 705830
rect 575234 704602 575266 704838
rect 575502 704602 575586 704838
rect 575822 704602 575854 704838
rect 575234 704518 575854 704602
rect 575234 704282 575266 704518
rect 575502 704282 575586 704518
rect 575822 704282 575854 704518
rect 575234 687454 575854 704282
rect 575234 687218 575266 687454
rect 575502 687218 575586 687454
rect 575822 687218 575854 687454
rect 575234 687134 575854 687218
rect 575234 686898 575266 687134
rect 575502 686898 575586 687134
rect 575822 686898 575854 687134
rect 575234 651454 575854 686898
rect 575234 651218 575266 651454
rect 575502 651218 575586 651454
rect 575822 651218 575854 651454
rect 575234 651134 575854 651218
rect 575234 650898 575266 651134
rect 575502 650898 575586 651134
rect 575822 650898 575854 651134
rect 575234 615454 575854 650898
rect 575234 615218 575266 615454
rect 575502 615218 575586 615454
rect 575822 615218 575854 615454
rect 575234 615134 575854 615218
rect 575234 614898 575266 615134
rect 575502 614898 575586 615134
rect 575822 614898 575854 615134
rect 575234 579454 575854 614898
rect 575234 579218 575266 579454
rect 575502 579218 575586 579454
rect 575822 579218 575854 579454
rect 575234 579134 575854 579218
rect 575234 578898 575266 579134
rect 575502 578898 575586 579134
rect 575822 578898 575854 579134
rect 575234 543454 575854 578898
rect 575234 543218 575266 543454
rect 575502 543218 575586 543454
rect 575822 543218 575854 543454
rect 575234 543134 575854 543218
rect 575234 542898 575266 543134
rect 575502 542898 575586 543134
rect 575822 542898 575854 543134
rect 575234 507454 575854 542898
rect 575234 507218 575266 507454
rect 575502 507218 575586 507454
rect 575822 507218 575854 507454
rect 575234 507134 575854 507218
rect 575234 506898 575266 507134
rect 575502 506898 575586 507134
rect 575822 506898 575854 507134
rect 575234 471454 575854 506898
rect 575234 471218 575266 471454
rect 575502 471218 575586 471454
rect 575822 471218 575854 471454
rect 575234 471134 575854 471218
rect 575234 470898 575266 471134
rect 575502 470898 575586 471134
rect 575822 470898 575854 471134
rect 575234 435454 575854 470898
rect 575234 435218 575266 435454
rect 575502 435218 575586 435454
rect 575822 435218 575854 435454
rect 575234 435134 575854 435218
rect 575234 434898 575266 435134
rect 575502 434898 575586 435134
rect 575822 434898 575854 435134
rect 575234 399454 575854 434898
rect 575234 399218 575266 399454
rect 575502 399218 575586 399454
rect 575822 399218 575854 399454
rect 575234 399134 575854 399218
rect 575234 398898 575266 399134
rect 575502 398898 575586 399134
rect 575822 398898 575854 399134
rect 575234 363454 575854 398898
rect 575234 363218 575266 363454
rect 575502 363218 575586 363454
rect 575822 363218 575854 363454
rect 575234 363134 575854 363218
rect 575234 362898 575266 363134
rect 575502 362898 575586 363134
rect 575822 362898 575854 363134
rect 575234 327454 575854 362898
rect 575234 327218 575266 327454
rect 575502 327218 575586 327454
rect 575822 327218 575854 327454
rect 575234 327134 575854 327218
rect 575234 326898 575266 327134
rect 575502 326898 575586 327134
rect 575822 326898 575854 327134
rect 575234 291454 575854 326898
rect 575234 291218 575266 291454
rect 575502 291218 575586 291454
rect 575822 291218 575854 291454
rect 575234 291134 575854 291218
rect 575234 290898 575266 291134
rect 575502 290898 575586 291134
rect 575822 290898 575854 291134
rect 575234 255454 575854 290898
rect 575234 255218 575266 255454
rect 575502 255218 575586 255454
rect 575822 255218 575854 255454
rect 575234 255134 575854 255218
rect 575234 254898 575266 255134
rect 575502 254898 575586 255134
rect 575822 254898 575854 255134
rect 575234 219454 575854 254898
rect 575234 219218 575266 219454
rect 575502 219218 575586 219454
rect 575822 219218 575854 219454
rect 575234 219134 575854 219218
rect 575234 218898 575266 219134
rect 575502 218898 575586 219134
rect 575822 218898 575854 219134
rect 575234 183454 575854 218898
rect 575234 183218 575266 183454
rect 575502 183218 575586 183454
rect 575822 183218 575854 183454
rect 575234 183134 575854 183218
rect 575234 182898 575266 183134
rect 575502 182898 575586 183134
rect 575822 182898 575854 183134
rect 575234 147454 575854 182898
rect 575234 147218 575266 147454
rect 575502 147218 575586 147454
rect 575822 147218 575854 147454
rect 575234 147134 575854 147218
rect 575234 146898 575266 147134
rect 575502 146898 575586 147134
rect 575822 146898 575854 147134
rect 575234 111454 575854 146898
rect 575234 111218 575266 111454
rect 575502 111218 575586 111454
rect 575822 111218 575854 111454
rect 575234 111134 575854 111218
rect 575234 110898 575266 111134
rect 575502 110898 575586 111134
rect 575822 110898 575854 111134
rect 575234 75454 575854 110898
rect 575234 75218 575266 75454
rect 575502 75218 575586 75454
rect 575822 75218 575854 75454
rect 575234 75134 575854 75218
rect 575234 74898 575266 75134
rect 575502 74898 575586 75134
rect 575822 74898 575854 75134
rect 575234 39454 575854 74898
rect 575234 39218 575266 39454
rect 575502 39218 575586 39454
rect 575822 39218 575854 39454
rect 575234 39134 575854 39218
rect 575234 38898 575266 39134
rect 575502 38898 575586 39134
rect 575822 38898 575854 39134
rect 575234 3454 575854 38898
rect 575234 3218 575266 3454
rect 575502 3218 575586 3454
rect 575822 3218 575854 3454
rect 575234 3134 575854 3218
rect 575234 2898 575266 3134
rect 575502 2898 575586 3134
rect 575822 2898 575854 3134
rect 575234 -346 575854 2898
rect 575234 -582 575266 -346
rect 575502 -582 575586 -346
rect 575822 -582 575854 -346
rect 575234 -666 575854 -582
rect 575234 -902 575266 -666
rect 575502 -902 575586 -666
rect 575822 -902 575854 -666
rect 575234 -1894 575854 -902
rect 576154 698614 576774 710042
rect 581274 711558 581894 711590
rect 581274 711322 581306 711558
rect 581542 711322 581626 711558
rect 581862 711322 581894 711558
rect 581274 711238 581894 711322
rect 581274 711002 581306 711238
rect 581542 711002 581626 711238
rect 581862 711002 581894 711238
rect 576154 698378 576186 698614
rect 576422 698378 576506 698614
rect 576742 698378 576774 698614
rect 576154 698294 576774 698378
rect 576154 698058 576186 698294
rect 576422 698058 576506 698294
rect 576742 698058 576774 698294
rect 576154 662614 576774 698058
rect 576154 662378 576186 662614
rect 576422 662378 576506 662614
rect 576742 662378 576774 662614
rect 576154 662294 576774 662378
rect 576154 662058 576186 662294
rect 576422 662058 576506 662294
rect 576742 662058 576774 662294
rect 576154 626614 576774 662058
rect 576154 626378 576186 626614
rect 576422 626378 576506 626614
rect 576742 626378 576774 626614
rect 576154 626294 576774 626378
rect 576154 626058 576186 626294
rect 576422 626058 576506 626294
rect 576742 626058 576774 626294
rect 576154 590614 576774 626058
rect 576154 590378 576186 590614
rect 576422 590378 576506 590614
rect 576742 590378 576774 590614
rect 576154 590294 576774 590378
rect 576154 590058 576186 590294
rect 576422 590058 576506 590294
rect 576742 590058 576774 590294
rect 576154 554614 576774 590058
rect 576154 554378 576186 554614
rect 576422 554378 576506 554614
rect 576742 554378 576774 554614
rect 576154 554294 576774 554378
rect 576154 554058 576186 554294
rect 576422 554058 576506 554294
rect 576742 554058 576774 554294
rect 576154 518614 576774 554058
rect 576154 518378 576186 518614
rect 576422 518378 576506 518614
rect 576742 518378 576774 518614
rect 576154 518294 576774 518378
rect 576154 518058 576186 518294
rect 576422 518058 576506 518294
rect 576742 518058 576774 518294
rect 576154 482614 576774 518058
rect 576154 482378 576186 482614
rect 576422 482378 576506 482614
rect 576742 482378 576774 482614
rect 576154 482294 576774 482378
rect 576154 482058 576186 482294
rect 576422 482058 576506 482294
rect 576742 482058 576774 482294
rect 576154 446614 576774 482058
rect 576154 446378 576186 446614
rect 576422 446378 576506 446614
rect 576742 446378 576774 446614
rect 576154 446294 576774 446378
rect 576154 446058 576186 446294
rect 576422 446058 576506 446294
rect 576742 446058 576774 446294
rect 576154 410614 576774 446058
rect 576154 410378 576186 410614
rect 576422 410378 576506 410614
rect 576742 410378 576774 410614
rect 576154 410294 576774 410378
rect 576154 410058 576186 410294
rect 576422 410058 576506 410294
rect 576742 410058 576774 410294
rect 576154 374614 576774 410058
rect 576154 374378 576186 374614
rect 576422 374378 576506 374614
rect 576742 374378 576774 374614
rect 576154 374294 576774 374378
rect 576154 374058 576186 374294
rect 576422 374058 576506 374294
rect 576742 374058 576774 374294
rect 576154 338614 576774 374058
rect 576154 338378 576186 338614
rect 576422 338378 576506 338614
rect 576742 338378 576774 338614
rect 576154 338294 576774 338378
rect 576154 338058 576186 338294
rect 576422 338058 576506 338294
rect 576742 338058 576774 338294
rect 576154 302614 576774 338058
rect 576154 302378 576186 302614
rect 576422 302378 576506 302614
rect 576742 302378 576774 302614
rect 576154 302294 576774 302378
rect 576154 302058 576186 302294
rect 576422 302058 576506 302294
rect 576742 302058 576774 302294
rect 576154 266614 576774 302058
rect 576154 266378 576186 266614
rect 576422 266378 576506 266614
rect 576742 266378 576774 266614
rect 576154 266294 576774 266378
rect 576154 266058 576186 266294
rect 576422 266058 576506 266294
rect 576742 266058 576774 266294
rect 576154 230614 576774 266058
rect 576154 230378 576186 230614
rect 576422 230378 576506 230614
rect 576742 230378 576774 230614
rect 576154 230294 576774 230378
rect 576154 230058 576186 230294
rect 576422 230058 576506 230294
rect 576742 230058 576774 230294
rect 576154 194614 576774 230058
rect 576154 194378 576186 194614
rect 576422 194378 576506 194614
rect 576742 194378 576774 194614
rect 576154 194294 576774 194378
rect 576154 194058 576186 194294
rect 576422 194058 576506 194294
rect 576742 194058 576774 194294
rect 576154 158614 576774 194058
rect 576154 158378 576186 158614
rect 576422 158378 576506 158614
rect 576742 158378 576774 158614
rect 576154 158294 576774 158378
rect 576154 158058 576186 158294
rect 576422 158058 576506 158294
rect 576742 158058 576774 158294
rect 576154 122614 576774 158058
rect 576154 122378 576186 122614
rect 576422 122378 576506 122614
rect 576742 122378 576774 122614
rect 576154 122294 576774 122378
rect 576154 122058 576186 122294
rect 576422 122058 576506 122294
rect 576742 122058 576774 122294
rect 576154 86614 576774 122058
rect 576154 86378 576186 86614
rect 576422 86378 576506 86614
rect 576742 86378 576774 86614
rect 576154 86294 576774 86378
rect 576154 86058 576186 86294
rect 576422 86058 576506 86294
rect 576742 86058 576774 86294
rect 576154 50614 576774 86058
rect 576154 50378 576186 50614
rect 576422 50378 576506 50614
rect 576742 50378 576774 50614
rect 576154 50294 576774 50378
rect 576154 50058 576186 50294
rect 576422 50058 576506 50294
rect 576742 50058 576774 50294
rect 576154 14614 576774 50058
rect 576154 14378 576186 14614
rect 576422 14378 576506 14614
rect 576742 14378 576774 14614
rect 576154 14294 576774 14378
rect 576154 14058 576186 14294
rect 576422 14058 576506 14294
rect 576742 14058 576774 14294
rect 573834 -3462 573866 -3226
rect 574102 -3462 574186 -3226
rect 574422 -3462 574454 -3226
rect 573834 -3546 574454 -3462
rect 573834 -3782 573866 -3546
rect 574102 -3782 574186 -3546
rect 574422 -3782 574454 -3546
rect 573834 -3814 574454 -3782
rect 572434 -4422 572466 -4186
rect 572702 -4422 572786 -4186
rect 573022 -4422 573054 -4186
rect 572434 -4506 573054 -4422
rect 572434 -4742 572466 -4506
rect 572702 -4742 572786 -4506
rect 573022 -4742 573054 -4506
rect 572434 -5734 573054 -4742
rect 571034 -7302 571066 -7066
rect 571302 -7302 571386 -7066
rect 571622 -7302 571654 -7066
rect 571034 -7386 571654 -7302
rect 571034 -7622 571066 -7386
rect 571302 -7622 571386 -7386
rect 571622 -7622 571654 -7386
rect 571034 -7654 571654 -7622
rect 576154 -6106 576774 14058
rect 577554 709638 578174 709670
rect 577554 709402 577586 709638
rect 577822 709402 577906 709638
rect 578142 709402 578174 709638
rect 577554 709318 578174 709402
rect 577554 709082 577586 709318
rect 577822 709082 577906 709318
rect 578142 709082 578174 709318
rect 577554 676894 578174 709082
rect 577554 676658 577586 676894
rect 577822 676658 577906 676894
rect 578142 676658 578174 676894
rect 577554 676574 578174 676658
rect 577554 676338 577586 676574
rect 577822 676338 577906 676574
rect 578142 676338 578174 676574
rect 577554 640894 578174 676338
rect 577554 640658 577586 640894
rect 577822 640658 577906 640894
rect 578142 640658 578174 640894
rect 577554 640574 578174 640658
rect 577554 640338 577586 640574
rect 577822 640338 577906 640574
rect 578142 640338 578174 640574
rect 577554 604894 578174 640338
rect 577554 604658 577586 604894
rect 577822 604658 577906 604894
rect 578142 604658 578174 604894
rect 577554 604574 578174 604658
rect 577554 604338 577586 604574
rect 577822 604338 577906 604574
rect 578142 604338 578174 604574
rect 577554 568894 578174 604338
rect 577554 568658 577586 568894
rect 577822 568658 577906 568894
rect 578142 568658 578174 568894
rect 577554 568574 578174 568658
rect 577554 568338 577586 568574
rect 577822 568338 577906 568574
rect 578142 568338 578174 568574
rect 577554 532894 578174 568338
rect 577554 532658 577586 532894
rect 577822 532658 577906 532894
rect 578142 532658 578174 532894
rect 577554 532574 578174 532658
rect 577554 532338 577586 532574
rect 577822 532338 577906 532574
rect 578142 532338 578174 532574
rect 577554 496894 578174 532338
rect 577554 496658 577586 496894
rect 577822 496658 577906 496894
rect 578142 496658 578174 496894
rect 577554 496574 578174 496658
rect 577554 496338 577586 496574
rect 577822 496338 577906 496574
rect 578142 496338 578174 496574
rect 577554 460894 578174 496338
rect 577554 460658 577586 460894
rect 577822 460658 577906 460894
rect 578142 460658 578174 460894
rect 577554 460574 578174 460658
rect 577554 460338 577586 460574
rect 577822 460338 577906 460574
rect 578142 460338 578174 460574
rect 577554 424894 578174 460338
rect 577554 424658 577586 424894
rect 577822 424658 577906 424894
rect 578142 424658 578174 424894
rect 577554 424574 578174 424658
rect 577554 424338 577586 424574
rect 577822 424338 577906 424574
rect 578142 424338 578174 424574
rect 577554 388894 578174 424338
rect 577554 388658 577586 388894
rect 577822 388658 577906 388894
rect 578142 388658 578174 388894
rect 577554 388574 578174 388658
rect 577554 388338 577586 388574
rect 577822 388338 577906 388574
rect 578142 388338 578174 388574
rect 577554 352894 578174 388338
rect 577554 352658 577586 352894
rect 577822 352658 577906 352894
rect 578142 352658 578174 352894
rect 577554 352574 578174 352658
rect 577554 352338 577586 352574
rect 577822 352338 577906 352574
rect 578142 352338 578174 352574
rect 577554 316894 578174 352338
rect 577554 316658 577586 316894
rect 577822 316658 577906 316894
rect 578142 316658 578174 316894
rect 577554 316574 578174 316658
rect 577554 316338 577586 316574
rect 577822 316338 577906 316574
rect 578142 316338 578174 316574
rect 577554 280894 578174 316338
rect 577554 280658 577586 280894
rect 577822 280658 577906 280894
rect 578142 280658 578174 280894
rect 577554 280574 578174 280658
rect 577554 280338 577586 280574
rect 577822 280338 577906 280574
rect 578142 280338 578174 280574
rect 577554 244894 578174 280338
rect 577554 244658 577586 244894
rect 577822 244658 577906 244894
rect 578142 244658 578174 244894
rect 577554 244574 578174 244658
rect 577554 244338 577586 244574
rect 577822 244338 577906 244574
rect 578142 244338 578174 244574
rect 577554 208894 578174 244338
rect 577554 208658 577586 208894
rect 577822 208658 577906 208894
rect 578142 208658 578174 208894
rect 577554 208574 578174 208658
rect 577554 208338 577586 208574
rect 577822 208338 577906 208574
rect 578142 208338 578174 208574
rect 577554 172894 578174 208338
rect 577554 172658 577586 172894
rect 577822 172658 577906 172894
rect 578142 172658 578174 172894
rect 577554 172574 578174 172658
rect 577554 172338 577586 172574
rect 577822 172338 577906 172574
rect 578142 172338 578174 172574
rect 577554 136894 578174 172338
rect 577554 136658 577586 136894
rect 577822 136658 577906 136894
rect 578142 136658 578174 136894
rect 577554 136574 578174 136658
rect 577554 136338 577586 136574
rect 577822 136338 577906 136574
rect 578142 136338 578174 136574
rect 577554 100894 578174 136338
rect 577554 100658 577586 100894
rect 577822 100658 577906 100894
rect 578142 100658 578174 100894
rect 577554 100574 578174 100658
rect 577554 100338 577586 100574
rect 577822 100338 577906 100574
rect 578142 100338 578174 100574
rect 577554 64894 578174 100338
rect 577554 64658 577586 64894
rect 577822 64658 577906 64894
rect 578142 64658 578174 64894
rect 577554 64574 578174 64658
rect 577554 64338 577586 64574
rect 577822 64338 577906 64574
rect 578142 64338 578174 64574
rect 577554 28894 578174 64338
rect 577554 28658 577586 28894
rect 577822 28658 577906 28894
rect 578142 28658 578174 28894
rect 577554 28574 578174 28658
rect 577554 28338 577586 28574
rect 577822 28338 577906 28574
rect 578142 28338 578174 28574
rect 577554 -5146 578174 28338
rect 578954 706758 579574 707750
rect 578954 706522 578986 706758
rect 579222 706522 579306 706758
rect 579542 706522 579574 706758
rect 578954 706438 579574 706522
rect 578954 706202 578986 706438
rect 579222 706202 579306 706438
rect 579542 706202 579574 706438
rect 578954 691174 579574 706202
rect 578954 690938 578986 691174
rect 579222 690938 579306 691174
rect 579542 690938 579574 691174
rect 578954 690854 579574 690938
rect 578954 690618 578986 690854
rect 579222 690618 579306 690854
rect 579542 690618 579574 690854
rect 578954 655174 579574 690618
rect 578954 654938 578986 655174
rect 579222 654938 579306 655174
rect 579542 654938 579574 655174
rect 578954 654854 579574 654938
rect 578954 654618 578986 654854
rect 579222 654618 579306 654854
rect 579542 654618 579574 654854
rect 578954 619174 579574 654618
rect 578954 618938 578986 619174
rect 579222 618938 579306 619174
rect 579542 618938 579574 619174
rect 578954 618854 579574 618938
rect 578954 618618 578986 618854
rect 579222 618618 579306 618854
rect 579542 618618 579574 618854
rect 578954 583174 579574 618618
rect 578954 582938 578986 583174
rect 579222 582938 579306 583174
rect 579542 582938 579574 583174
rect 578954 582854 579574 582938
rect 578954 582618 578986 582854
rect 579222 582618 579306 582854
rect 579542 582618 579574 582854
rect 578954 547174 579574 582618
rect 578954 546938 578986 547174
rect 579222 546938 579306 547174
rect 579542 546938 579574 547174
rect 578954 546854 579574 546938
rect 578954 546618 578986 546854
rect 579222 546618 579306 546854
rect 579542 546618 579574 546854
rect 578954 511174 579574 546618
rect 578954 510938 578986 511174
rect 579222 510938 579306 511174
rect 579542 510938 579574 511174
rect 578954 510854 579574 510938
rect 578954 510618 578986 510854
rect 579222 510618 579306 510854
rect 579542 510618 579574 510854
rect 578954 475174 579574 510618
rect 578954 474938 578986 475174
rect 579222 474938 579306 475174
rect 579542 474938 579574 475174
rect 578954 474854 579574 474938
rect 578954 474618 578986 474854
rect 579222 474618 579306 474854
rect 579542 474618 579574 474854
rect 578954 439174 579574 474618
rect 578954 438938 578986 439174
rect 579222 438938 579306 439174
rect 579542 438938 579574 439174
rect 578954 438854 579574 438938
rect 578954 438618 578986 438854
rect 579222 438618 579306 438854
rect 579542 438618 579574 438854
rect 578954 403174 579574 438618
rect 578954 402938 578986 403174
rect 579222 402938 579306 403174
rect 579542 402938 579574 403174
rect 578954 402854 579574 402938
rect 578954 402618 578986 402854
rect 579222 402618 579306 402854
rect 579542 402618 579574 402854
rect 578954 367174 579574 402618
rect 578954 366938 578986 367174
rect 579222 366938 579306 367174
rect 579542 366938 579574 367174
rect 578954 366854 579574 366938
rect 578954 366618 578986 366854
rect 579222 366618 579306 366854
rect 579542 366618 579574 366854
rect 578954 331174 579574 366618
rect 578954 330938 578986 331174
rect 579222 330938 579306 331174
rect 579542 330938 579574 331174
rect 578954 330854 579574 330938
rect 578954 330618 578986 330854
rect 579222 330618 579306 330854
rect 579542 330618 579574 330854
rect 578954 295174 579574 330618
rect 578954 294938 578986 295174
rect 579222 294938 579306 295174
rect 579542 294938 579574 295174
rect 578954 294854 579574 294938
rect 578954 294618 578986 294854
rect 579222 294618 579306 294854
rect 579542 294618 579574 294854
rect 578954 259174 579574 294618
rect 578954 258938 578986 259174
rect 579222 258938 579306 259174
rect 579542 258938 579574 259174
rect 578954 258854 579574 258938
rect 578954 258618 578986 258854
rect 579222 258618 579306 258854
rect 579542 258618 579574 258854
rect 578954 223174 579574 258618
rect 578954 222938 578986 223174
rect 579222 222938 579306 223174
rect 579542 222938 579574 223174
rect 578954 222854 579574 222938
rect 578954 222618 578986 222854
rect 579222 222618 579306 222854
rect 579542 222618 579574 222854
rect 578954 187174 579574 222618
rect 578954 186938 578986 187174
rect 579222 186938 579306 187174
rect 579542 186938 579574 187174
rect 578954 186854 579574 186938
rect 578954 186618 578986 186854
rect 579222 186618 579306 186854
rect 579542 186618 579574 186854
rect 578954 151174 579574 186618
rect 578954 150938 578986 151174
rect 579222 150938 579306 151174
rect 579542 150938 579574 151174
rect 578954 150854 579574 150938
rect 578954 150618 578986 150854
rect 579222 150618 579306 150854
rect 579542 150618 579574 150854
rect 578954 115174 579574 150618
rect 578954 114938 578986 115174
rect 579222 114938 579306 115174
rect 579542 114938 579574 115174
rect 578954 114854 579574 114938
rect 578954 114618 578986 114854
rect 579222 114618 579306 114854
rect 579542 114618 579574 114854
rect 578954 79174 579574 114618
rect 578954 78938 578986 79174
rect 579222 78938 579306 79174
rect 579542 78938 579574 79174
rect 578954 78854 579574 78938
rect 578954 78618 578986 78854
rect 579222 78618 579306 78854
rect 579542 78618 579574 78854
rect 578954 43174 579574 78618
rect 578954 42938 578986 43174
rect 579222 42938 579306 43174
rect 579542 42938 579574 43174
rect 578954 42854 579574 42938
rect 578954 42618 578986 42854
rect 579222 42618 579306 42854
rect 579542 42618 579574 42854
rect 578954 7174 579574 42618
rect 578954 6938 578986 7174
rect 579222 6938 579306 7174
rect 579542 6938 579574 7174
rect 578954 6854 579574 6938
rect 578954 6618 578986 6854
rect 579222 6618 579306 6854
rect 579542 6618 579574 6854
rect 578954 -2266 579574 6618
rect 580354 705798 580974 705830
rect 580354 705562 580386 705798
rect 580622 705562 580706 705798
rect 580942 705562 580974 705798
rect 580354 705478 580974 705562
rect 580354 705242 580386 705478
rect 580622 705242 580706 705478
rect 580942 705242 580974 705478
rect 580354 669454 580974 705242
rect 580354 669218 580386 669454
rect 580622 669218 580706 669454
rect 580942 669218 580974 669454
rect 580354 669134 580974 669218
rect 580354 668898 580386 669134
rect 580622 668898 580706 669134
rect 580942 668898 580974 669134
rect 580354 633454 580974 668898
rect 580354 633218 580386 633454
rect 580622 633218 580706 633454
rect 580942 633218 580974 633454
rect 580354 633134 580974 633218
rect 580354 632898 580386 633134
rect 580622 632898 580706 633134
rect 580942 632898 580974 633134
rect 580354 597454 580974 632898
rect 580354 597218 580386 597454
rect 580622 597218 580706 597454
rect 580942 597218 580974 597454
rect 580354 597134 580974 597218
rect 580354 596898 580386 597134
rect 580622 596898 580706 597134
rect 580942 596898 580974 597134
rect 580354 561454 580974 596898
rect 580354 561218 580386 561454
rect 580622 561218 580706 561454
rect 580942 561218 580974 561454
rect 580354 561134 580974 561218
rect 580354 560898 580386 561134
rect 580622 560898 580706 561134
rect 580942 560898 580974 561134
rect 580354 525454 580974 560898
rect 580354 525218 580386 525454
rect 580622 525218 580706 525454
rect 580942 525218 580974 525454
rect 580354 525134 580974 525218
rect 580354 524898 580386 525134
rect 580622 524898 580706 525134
rect 580942 524898 580974 525134
rect 580354 489454 580974 524898
rect 580354 489218 580386 489454
rect 580622 489218 580706 489454
rect 580942 489218 580974 489454
rect 580354 489134 580974 489218
rect 580354 488898 580386 489134
rect 580622 488898 580706 489134
rect 580942 488898 580974 489134
rect 580354 453454 580974 488898
rect 580354 453218 580386 453454
rect 580622 453218 580706 453454
rect 580942 453218 580974 453454
rect 580354 453134 580974 453218
rect 580354 452898 580386 453134
rect 580622 452898 580706 453134
rect 580942 452898 580974 453134
rect 580354 417454 580974 452898
rect 580354 417218 580386 417454
rect 580622 417218 580706 417454
rect 580942 417218 580974 417454
rect 580354 417134 580974 417218
rect 580354 416898 580386 417134
rect 580622 416898 580706 417134
rect 580942 416898 580974 417134
rect 580354 381454 580974 416898
rect 580354 381218 580386 381454
rect 580622 381218 580706 381454
rect 580942 381218 580974 381454
rect 580354 381134 580974 381218
rect 580354 380898 580386 381134
rect 580622 380898 580706 381134
rect 580942 380898 580974 381134
rect 580354 345454 580974 380898
rect 580354 345218 580386 345454
rect 580622 345218 580706 345454
rect 580942 345218 580974 345454
rect 580354 345134 580974 345218
rect 580354 344898 580386 345134
rect 580622 344898 580706 345134
rect 580942 344898 580974 345134
rect 580354 309454 580974 344898
rect 580354 309218 580386 309454
rect 580622 309218 580706 309454
rect 580942 309218 580974 309454
rect 580354 309134 580974 309218
rect 580354 308898 580386 309134
rect 580622 308898 580706 309134
rect 580942 308898 580974 309134
rect 580354 273454 580974 308898
rect 580354 273218 580386 273454
rect 580622 273218 580706 273454
rect 580942 273218 580974 273454
rect 580354 273134 580974 273218
rect 580354 272898 580386 273134
rect 580622 272898 580706 273134
rect 580942 272898 580974 273134
rect 580354 237454 580974 272898
rect 580354 237218 580386 237454
rect 580622 237218 580706 237454
rect 580942 237218 580974 237454
rect 580354 237134 580974 237218
rect 580354 236898 580386 237134
rect 580622 236898 580706 237134
rect 580942 236898 580974 237134
rect 580354 201454 580974 236898
rect 580354 201218 580386 201454
rect 580622 201218 580706 201454
rect 580942 201218 580974 201454
rect 580354 201134 580974 201218
rect 580354 200898 580386 201134
rect 580622 200898 580706 201134
rect 580942 200898 580974 201134
rect 580354 165454 580974 200898
rect 580354 165218 580386 165454
rect 580622 165218 580706 165454
rect 580942 165218 580974 165454
rect 580354 165134 580974 165218
rect 580354 164898 580386 165134
rect 580622 164898 580706 165134
rect 580942 164898 580974 165134
rect 580354 129454 580974 164898
rect 580354 129218 580386 129454
rect 580622 129218 580706 129454
rect 580942 129218 580974 129454
rect 580354 129134 580974 129218
rect 580354 128898 580386 129134
rect 580622 128898 580706 129134
rect 580942 128898 580974 129134
rect 580354 93454 580974 128898
rect 580354 93218 580386 93454
rect 580622 93218 580706 93454
rect 580942 93218 580974 93454
rect 580354 93134 580974 93218
rect 580354 92898 580386 93134
rect 580622 92898 580706 93134
rect 580942 92898 580974 93134
rect 580354 57454 580974 92898
rect 580354 57218 580386 57454
rect 580622 57218 580706 57454
rect 580942 57218 580974 57454
rect 580354 57134 580974 57218
rect 580354 56898 580386 57134
rect 580622 56898 580706 57134
rect 580942 56898 580974 57134
rect 580354 21454 580974 56898
rect 580354 21218 580386 21454
rect 580622 21218 580706 21454
rect 580942 21218 580974 21454
rect 580354 21134 580974 21218
rect 580354 20898 580386 21134
rect 580622 20898 580706 21134
rect 580942 20898 580974 21134
rect 580354 -1306 580974 20898
rect 580354 -1542 580386 -1306
rect 580622 -1542 580706 -1306
rect 580942 -1542 580974 -1306
rect 580354 -1626 580974 -1542
rect 580354 -1862 580386 -1626
rect 580622 -1862 580706 -1626
rect 580942 -1862 580974 -1626
rect 580354 -1894 580974 -1862
rect 581274 680614 581894 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581274 680378 581306 680614
rect 581542 680378 581626 680614
rect 581862 680378 581894 680614
rect 581274 680294 581894 680378
rect 581274 680058 581306 680294
rect 581542 680058 581626 680294
rect 581862 680058 581894 680294
rect 581274 644614 581894 680058
rect 581274 644378 581306 644614
rect 581542 644378 581626 644614
rect 581862 644378 581894 644614
rect 581274 644294 581894 644378
rect 581274 644058 581306 644294
rect 581542 644058 581626 644294
rect 581862 644058 581894 644294
rect 581274 608614 581894 644058
rect 581274 608378 581306 608614
rect 581542 608378 581626 608614
rect 581862 608378 581894 608614
rect 581274 608294 581894 608378
rect 581274 608058 581306 608294
rect 581542 608058 581626 608294
rect 581862 608058 581894 608294
rect 581274 572614 581894 608058
rect 581274 572378 581306 572614
rect 581542 572378 581626 572614
rect 581862 572378 581894 572614
rect 581274 572294 581894 572378
rect 581274 572058 581306 572294
rect 581542 572058 581626 572294
rect 581862 572058 581894 572294
rect 581274 536614 581894 572058
rect 581274 536378 581306 536614
rect 581542 536378 581626 536614
rect 581862 536378 581894 536614
rect 581274 536294 581894 536378
rect 581274 536058 581306 536294
rect 581542 536058 581626 536294
rect 581862 536058 581894 536294
rect 581274 500614 581894 536058
rect 581274 500378 581306 500614
rect 581542 500378 581626 500614
rect 581862 500378 581894 500614
rect 581274 500294 581894 500378
rect 581274 500058 581306 500294
rect 581542 500058 581626 500294
rect 581862 500058 581894 500294
rect 581274 464614 581894 500058
rect 581274 464378 581306 464614
rect 581542 464378 581626 464614
rect 581862 464378 581894 464614
rect 581274 464294 581894 464378
rect 581274 464058 581306 464294
rect 581542 464058 581626 464294
rect 581862 464058 581894 464294
rect 581274 428614 581894 464058
rect 581274 428378 581306 428614
rect 581542 428378 581626 428614
rect 581862 428378 581894 428614
rect 581274 428294 581894 428378
rect 581274 428058 581306 428294
rect 581542 428058 581626 428294
rect 581862 428058 581894 428294
rect 581274 392614 581894 428058
rect 581274 392378 581306 392614
rect 581542 392378 581626 392614
rect 581862 392378 581894 392614
rect 581274 392294 581894 392378
rect 581274 392058 581306 392294
rect 581542 392058 581626 392294
rect 581862 392058 581894 392294
rect 581274 356614 581894 392058
rect 581274 356378 581306 356614
rect 581542 356378 581626 356614
rect 581862 356378 581894 356614
rect 581274 356294 581894 356378
rect 581274 356058 581306 356294
rect 581542 356058 581626 356294
rect 581862 356058 581894 356294
rect 581274 320614 581894 356058
rect 581274 320378 581306 320614
rect 581542 320378 581626 320614
rect 581862 320378 581894 320614
rect 581274 320294 581894 320378
rect 581274 320058 581306 320294
rect 581542 320058 581626 320294
rect 581862 320058 581894 320294
rect 581274 284614 581894 320058
rect 581274 284378 581306 284614
rect 581542 284378 581626 284614
rect 581862 284378 581894 284614
rect 581274 284294 581894 284378
rect 581274 284058 581306 284294
rect 581542 284058 581626 284294
rect 581862 284058 581894 284294
rect 581274 248614 581894 284058
rect 581274 248378 581306 248614
rect 581542 248378 581626 248614
rect 581862 248378 581894 248614
rect 581274 248294 581894 248378
rect 581274 248058 581306 248294
rect 581542 248058 581626 248294
rect 581862 248058 581894 248294
rect 581274 212614 581894 248058
rect 581274 212378 581306 212614
rect 581542 212378 581626 212614
rect 581862 212378 581894 212614
rect 581274 212294 581894 212378
rect 581274 212058 581306 212294
rect 581542 212058 581626 212294
rect 581862 212058 581894 212294
rect 581274 176614 581894 212058
rect 581274 176378 581306 176614
rect 581542 176378 581626 176614
rect 581862 176378 581894 176614
rect 581274 176294 581894 176378
rect 581274 176058 581306 176294
rect 581542 176058 581626 176294
rect 581862 176058 581894 176294
rect 581274 140614 581894 176058
rect 581274 140378 581306 140614
rect 581542 140378 581626 140614
rect 581862 140378 581894 140614
rect 581274 140294 581894 140378
rect 581274 140058 581306 140294
rect 581542 140058 581626 140294
rect 581862 140058 581894 140294
rect 581274 104614 581894 140058
rect 581274 104378 581306 104614
rect 581542 104378 581626 104614
rect 581862 104378 581894 104614
rect 581274 104294 581894 104378
rect 581274 104058 581306 104294
rect 581542 104058 581626 104294
rect 581862 104058 581894 104294
rect 581274 68614 581894 104058
rect 581274 68378 581306 68614
rect 581542 68378 581626 68614
rect 581862 68378 581894 68614
rect 581274 68294 581894 68378
rect 581274 68058 581306 68294
rect 581542 68058 581626 68294
rect 581862 68058 581894 68294
rect 581274 32614 581894 68058
rect 581274 32378 581306 32614
rect 581542 32378 581626 32614
rect 581862 32378 581894 32614
rect 581274 32294 581894 32378
rect 581274 32058 581306 32294
rect 581542 32058 581626 32294
rect 581862 32058 581894 32294
rect 578954 -2502 578986 -2266
rect 579222 -2502 579306 -2266
rect 579542 -2502 579574 -2266
rect 578954 -2586 579574 -2502
rect 578954 -2822 578986 -2586
rect 579222 -2822 579306 -2586
rect 579542 -2822 579574 -2586
rect 578954 -3814 579574 -2822
rect 577554 -5382 577586 -5146
rect 577822 -5382 577906 -5146
rect 578142 -5382 578174 -5146
rect 577554 -5466 578174 -5382
rect 577554 -5702 577586 -5466
rect 577822 -5702 577906 -5466
rect 578142 -5702 578174 -5466
rect 577554 -5734 578174 -5702
rect 576154 -6342 576186 -6106
rect 576422 -6342 576506 -6106
rect 576742 -6342 576774 -6106
rect 576154 -6426 576774 -6342
rect 576154 -6662 576186 -6426
rect 576422 -6662 576506 -6426
rect 576742 -6662 576774 -6426
rect 576154 -7654 576774 -6662
rect 581274 -7066 581894 32058
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 581274 -7302 581306 -7066
rect 581542 -7302 581626 -7066
rect 581862 -7302 581894 -7066
rect 581274 -7386 581894 -7302
rect 581274 -7622 581306 -7386
rect 581542 -7622 581626 -7386
rect 581862 -7622 581894 -7386
rect 581274 -7654 581894 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 6946 705562 7182 705798
rect 7266 705562 7502 705798
rect 6946 705242 7182 705478
rect 7266 705242 7502 705478
rect 6946 669218 7182 669454
rect 7266 669218 7502 669454
rect 6946 668898 7182 669134
rect 7266 668898 7502 669134
rect 6946 633218 7182 633454
rect 7266 633218 7502 633454
rect 6946 632898 7182 633134
rect 7266 632898 7502 633134
rect 6946 597218 7182 597454
rect 7266 597218 7502 597454
rect 6946 596898 7182 597134
rect 7266 596898 7502 597134
rect 6946 561218 7182 561454
rect 7266 561218 7502 561454
rect 6946 560898 7182 561134
rect 7266 560898 7502 561134
rect 6946 525218 7182 525454
rect 7266 525218 7502 525454
rect 6946 524898 7182 525134
rect 7266 524898 7502 525134
rect 6946 489218 7182 489454
rect 7266 489218 7502 489454
rect 6946 488898 7182 489134
rect 7266 488898 7502 489134
rect 6946 453218 7182 453454
rect 7266 453218 7502 453454
rect 6946 452898 7182 453134
rect 7266 452898 7502 453134
rect 6946 417218 7182 417454
rect 7266 417218 7502 417454
rect 6946 416898 7182 417134
rect 7266 416898 7502 417134
rect 6946 381218 7182 381454
rect 7266 381218 7502 381454
rect 6946 380898 7182 381134
rect 7266 380898 7502 381134
rect 6946 345218 7182 345454
rect 7266 345218 7502 345454
rect 6946 344898 7182 345134
rect 7266 344898 7502 345134
rect 6946 309218 7182 309454
rect 7266 309218 7502 309454
rect 6946 308898 7182 309134
rect 7266 308898 7502 309134
rect 6946 273218 7182 273454
rect 7266 273218 7502 273454
rect 6946 272898 7182 273134
rect 7266 272898 7502 273134
rect 6946 237218 7182 237454
rect 7266 237218 7502 237454
rect 6946 236898 7182 237134
rect 7266 236898 7502 237134
rect 6946 201218 7182 201454
rect 7266 201218 7502 201454
rect 6946 200898 7182 201134
rect 7266 200898 7502 201134
rect 6946 165218 7182 165454
rect 7266 165218 7502 165454
rect 6946 164898 7182 165134
rect 7266 164898 7502 165134
rect 6946 129218 7182 129454
rect 7266 129218 7502 129454
rect 6946 128898 7182 129134
rect 7266 128898 7502 129134
rect 6946 93218 7182 93454
rect 7266 93218 7502 93454
rect 6946 92898 7182 93134
rect 7266 92898 7502 93134
rect 6946 57218 7182 57454
rect 7266 57218 7502 57454
rect 6946 56898 7182 57134
rect 7266 56898 7502 57134
rect 6946 21218 7182 21454
rect 7266 21218 7502 21454
rect 6946 20898 7182 21134
rect 7266 20898 7502 21134
rect 6946 -1542 7182 -1306
rect 7266 -1542 7502 -1306
rect 6946 -1862 7182 -1626
rect 7266 -1862 7502 -1626
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 10666 707482 10902 707718
rect 10986 707482 11222 707718
rect 10666 707162 10902 707398
rect 10986 707162 11222 707398
rect 10666 672938 10902 673174
rect 10986 672938 11222 673174
rect 10666 672618 10902 672854
rect 10986 672618 11222 672854
rect 10666 636938 10902 637174
rect 10986 636938 11222 637174
rect 10666 636618 10902 636854
rect 10986 636618 11222 636854
rect 10666 600938 10902 601174
rect 10986 600938 11222 601174
rect 10666 600618 10902 600854
rect 10986 600618 11222 600854
rect 10666 564938 10902 565174
rect 10986 564938 11222 565174
rect 10666 564618 10902 564854
rect 10986 564618 11222 564854
rect 10666 528938 10902 529174
rect 10986 528938 11222 529174
rect 10666 528618 10902 528854
rect 10986 528618 11222 528854
rect 10666 492938 10902 493174
rect 10986 492938 11222 493174
rect 10666 492618 10902 492854
rect 10986 492618 11222 492854
rect 10666 456938 10902 457174
rect 10986 456938 11222 457174
rect 10666 456618 10902 456854
rect 10986 456618 11222 456854
rect 10666 420938 10902 421174
rect 10986 420938 11222 421174
rect 10666 420618 10902 420854
rect 10986 420618 11222 420854
rect 10666 384938 10902 385174
rect 10986 384938 11222 385174
rect 10666 384618 10902 384854
rect 10986 384618 11222 384854
rect 10666 348938 10902 349174
rect 10986 348938 11222 349174
rect 10666 348618 10902 348854
rect 10986 348618 11222 348854
rect 10666 312938 10902 313174
rect 10986 312938 11222 313174
rect 10666 312618 10902 312854
rect 10986 312618 11222 312854
rect 10666 276938 10902 277174
rect 10986 276938 11222 277174
rect 10666 276618 10902 276854
rect 10986 276618 11222 276854
rect 10666 240938 10902 241174
rect 10986 240938 11222 241174
rect 10666 240618 10902 240854
rect 10986 240618 11222 240854
rect 10666 204938 10902 205174
rect 10986 204938 11222 205174
rect 10666 204618 10902 204854
rect 10986 204618 11222 204854
rect 10666 168938 10902 169174
rect 10986 168938 11222 169174
rect 10666 168618 10902 168854
rect 10986 168618 11222 168854
rect 10666 132938 10902 133174
rect 10986 132938 11222 133174
rect 10666 132618 10902 132854
rect 10986 132618 11222 132854
rect 10666 96938 10902 97174
rect 10986 96938 11222 97174
rect 10666 96618 10902 96854
rect 10986 96618 11222 96854
rect 10666 60938 10902 61174
rect 10986 60938 11222 61174
rect 10666 60618 10902 60854
rect 10986 60618 11222 60854
rect 10666 24938 10902 25174
rect 10986 24938 11222 25174
rect 10666 24618 10902 24854
rect 10986 24618 11222 24854
rect 12066 704602 12302 704838
rect 12386 704602 12622 704838
rect 12066 704282 12302 704518
rect 12386 704282 12622 704518
rect 12066 687218 12302 687454
rect 12386 687218 12622 687454
rect 12066 686898 12302 687134
rect 12386 686898 12622 687134
rect 12066 651218 12302 651454
rect 12386 651218 12622 651454
rect 12066 650898 12302 651134
rect 12386 650898 12622 651134
rect 12066 615218 12302 615454
rect 12386 615218 12622 615454
rect 12066 614898 12302 615134
rect 12386 614898 12622 615134
rect 12066 579218 12302 579454
rect 12386 579218 12622 579454
rect 12066 578898 12302 579134
rect 12386 578898 12622 579134
rect 12066 543218 12302 543454
rect 12386 543218 12622 543454
rect 12066 542898 12302 543134
rect 12386 542898 12622 543134
rect 12066 507218 12302 507454
rect 12386 507218 12622 507454
rect 12066 506898 12302 507134
rect 12386 506898 12622 507134
rect 12066 471218 12302 471454
rect 12386 471218 12622 471454
rect 12066 470898 12302 471134
rect 12386 470898 12622 471134
rect 12066 435218 12302 435454
rect 12386 435218 12622 435454
rect 12066 434898 12302 435134
rect 12386 434898 12622 435134
rect 12066 399218 12302 399454
rect 12386 399218 12622 399454
rect 12066 398898 12302 399134
rect 12386 398898 12622 399134
rect 12066 363218 12302 363454
rect 12386 363218 12622 363454
rect 12066 362898 12302 363134
rect 12386 362898 12622 363134
rect 12066 327218 12302 327454
rect 12386 327218 12622 327454
rect 12066 326898 12302 327134
rect 12386 326898 12622 327134
rect 12066 291218 12302 291454
rect 12386 291218 12622 291454
rect 12066 290898 12302 291134
rect 12386 290898 12622 291134
rect 12066 255218 12302 255454
rect 12386 255218 12622 255454
rect 12066 254898 12302 255134
rect 12386 254898 12622 255134
rect 12066 219218 12302 219454
rect 12386 219218 12622 219454
rect 12066 218898 12302 219134
rect 12386 218898 12622 219134
rect 12066 183218 12302 183454
rect 12386 183218 12622 183454
rect 12066 182898 12302 183134
rect 12386 182898 12622 183134
rect 12066 147218 12302 147454
rect 12386 147218 12622 147454
rect 12066 146898 12302 147134
rect 12386 146898 12622 147134
rect 12066 111218 12302 111454
rect 12386 111218 12622 111454
rect 12066 110898 12302 111134
rect 12386 110898 12622 111134
rect 12066 75218 12302 75454
rect 12386 75218 12622 75454
rect 12066 74898 12302 75134
rect 12386 74898 12622 75134
rect 12066 39218 12302 39454
rect 12386 39218 12622 39454
rect 12066 38898 12302 39134
rect 12386 38898 12622 39134
rect 12066 3218 12302 3454
rect 12386 3218 12622 3454
rect 12066 2898 12302 3134
rect 12386 2898 12622 3134
rect 12066 -582 12302 -346
rect 12386 -582 12622 -346
rect 12066 -902 12302 -666
rect 12386 -902 12622 -666
rect 18106 711322 18342 711558
rect 18426 711322 18662 711558
rect 18106 711002 18342 711238
rect 18426 711002 18662 711238
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 10666 -3462 10902 -3226
rect 10986 -3462 11222 -3226
rect 10666 -3782 10902 -3546
rect 10986 -3782 11222 -3546
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 14386 709402 14622 709638
rect 14706 709402 14942 709638
rect 14386 709082 14622 709318
rect 14706 709082 14942 709318
rect 14386 676658 14622 676894
rect 14706 676658 14942 676894
rect 14386 676338 14622 676574
rect 14706 676338 14942 676574
rect 14386 640658 14622 640894
rect 14706 640658 14942 640894
rect 14386 640338 14622 640574
rect 14706 640338 14942 640574
rect 14386 604658 14622 604894
rect 14706 604658 14942 604894
rect 14386 604338 14622 604574
rect 14706 604338 14942 604574
rect 14386 568658 14622 568894
rect 14706 568658 14942 568894
rect 14386 568338 14622 568574
rect 14706 568338 14942 568574
rect 14386 532658 14622 532894
rect 14706 532658 14942 532894
rect 14386 532338 14622 532574
rect 14706 532338 14942 532574
rect 14386 496658 14622 496894
rect 14706 496658 14942 496894
rect 14386 496338 14622 496574
rect 14706 496338 14942 496574
rect 14386 460658 14622 460894
rect 14706 460658 14942 460894
rect 14386 460338 14622 460574
rect 14706 460338 14942 460574
rect 14386 424658 14622 424894
rect 14706 424658 14942 424894
rect 14386 424338 14622 424574
rect 14706 424338 14942 424574
rect 14386 388658 14622 388894
rect 14706 388658 14942 388894
rect 14386 388338 14622 388574
rect 14706 388338 14942 388574
rect 14386 352658 14622 352894
rect 14706 352658 14942 352894
rect 14386 352338 14622 352574
rect 14706 352338 14942 352574
rect 14386 316658 14622 316894
rect 14706 316658 14942 316894
rect 14386 316338 14622 316574
rect 14706 316338 14942 316574
rect 14386 280658 14622 280894
rect 14706 280658 14942 280894
rect 14386 280338 14622 280574
rect 14706 280338 14942 280574
rect 14386 244658 14622 244894
rect 14706 244658 14942 244894
rect 14386 244338 14622 244574
rect 14706 244338 14942 244574
rect 14386 208658 14622 208894
rect 14706 208658 14942 208894
rect 14386 208338 14622 208574
rect 14706 208338 14942 208574
rect 14386 172658 14622 172894
rect 14706 172658 14942 172894
rect 14386 172338 14622 172574
rect 14706 172338 14942 172574
rect 14386 136658 14622 136894
rect 14706 136658 14942 136894
rect 14386 136338 14622 136574
rect 14706 136338 14942 136574
rect 14386 100658 14622 100894
rect 14706 100658 14942 100894
rect 14386 100338 14622 100574
rect 14706 100338 14942 100574
rect 14386 64658 14622 64894
rect 14706 64658 14942 64894
rect 14386 64338 14622 64574
rect 14706 64338 14942 64574
rect 14386 28658 14622 28894
rect 14706 28658 14942 28894
rect 14386 28338 14622 28574
rect 14706 28338 14942 28574
rect 15786 706522 16022 706758
rect 16106 706522 16342 706758
rect 15786 706202 16022 706438
rect 16106 706202 16342 706438
rect 15786 690938 16022 691174
rect 16106 690938 16342 691174
rect 15786 690618 16022 690854
rect 16106 690618 16342 690854
rect 17186 705562 17422 705798
rect 17506 705562 17742 705798
rect 17186 705242 17422 705478
rect 17506 705242 17742 705478
rect 17186 669218 17422 669454
rect 17506 669218 17742 669454
rect 17186 668898 17422 669134
rect 17506 668898 17742 669134
rect 23226 710362 23462 710598
rect 23546 710362 23782 710598
rect 23226 710042 23462 710278
rect 23546 710042 23782 710278
rect 18106 680378 18342 680614
rect 18426 680378 18662 680614
rect 18106 680058 18342 680294
rect 18426 680058 18662 680294
rect 19506 708442 19742 708678
rect 19826 708442 20062 708678
rect 19506 708122 19742 708358
rect 19826 708122 20062 708358
rect 19506 694658 19742 694894
rect 19826 694658 20062 694894
rect 19506 694338 19742 694574
rect 19826 694338 20062 694574
rect 19506 658658 19742 658894
rect 19826 658658 20062 658894
rect 19506 658338 19742 658574
rect 19826 658338 20062 658574
rect 20906 707482 21142 707718
rect 21226 707482 21462 707718
rect 20906 707162 21142 707398
rect 21226 707162 21462 707398
rect 20906 672938 21142 673174
rect 21226 672938 21462 673174
rect 20906 672618 21142 672854
rect 21226 672618 21462 672854
rect 22306 704602 22542 704838
rect 22626 704602 22862 704838
rect 22306 704282 22542 704518
rect 22626 704282 22862 704518
rect 22306 687218 22542 687454
rect 22626 687218 22862 687454
rect 22306 686898 22542 687134
rect 22626 686898 22862 687134
rect 28346 711322 28582 711558
rect 28666 711322 28902 711558
rect 28346 711002 28582 711238
rect 28666 711002 28902 711238
rect 23226 698378 23462 698614
rect 23546 698378 23782 698614
rect 23226 698058 23462 698294
rect 23546 698058 23782 698294
rect 23226 662378 23462 662614
rect 23546 662378 23782 662614
rect 23226 662058 23462 662294
rect 23546 662058 23782 662294
rect 24626 709402 24862 709638
rect 24946 709402 25182 709638
rect 24626 709082 24862 709318
rect 24946 709082 25182 709318
rect 24626 676658 24862 676894
rect 24946 676658 25182 676894
rect 24626 676338 24862 676574
rect 24946 676338 25182 676574
rect 26026 706522 26262 706758
rect 26346 706522 26582 706758
rect 26026 706202 26262 706438
rect 26346 706202 26582 706438
rect 26026 690938 26262 691174
rect 26346 690938 26582 691174
rect 26026 690618 26262 690854
rect 26346 690618 26582 690854
rect 27426 705562 27662 705798
rect 27746 705562 27982 705798
rect 27426 705242 27662 705478
rect 27746 705242 27982 705478
rect 27426 669218 27662 669454
rect 27746 669218 27982 669454
rect 27426 668898 27662 669134
rect 27746 668898 27982 669134
rect 33466 710362 33702 710598
rect 33786 710362 34022 710598
rect 33466 710042 33702 710278
rect 33786 710042 34022 710278
rect 28346 680378 28582 680614
rect 28666 680378 28902 680614
rect 28346 680058 28582 680294
rect 28666 680058 28902 680294
rect 29746 708442 29982 708678
rect 30066 708442 30302 708678
rect 29746 708122 29982 708358
rect 30066 708122 30302 708358
rect 29746 694658 29982 694894
rect 30066 694658 30302 694894
rect 29746 694338 29982 694574
rect 30066 694338 30302 694574
rect 29746 658658 29982 658894
rect 30066 658658 30302 658894
rect 29746 658338 29982 658574
rect 30066 658338 30302 658574
rect 31146 707482 31382 707718
rect 31466 707482 31702 707718
rect 31146 707162 31382 707398
rect 31466 707162 31702 707398
rect 31146 672938 31382 673174
rect 31466 672938 31702 673174
rect 31146 672618 31382 672854
rect 31466 672618 31702 672854
rect 32546 704602 32782 704838
rect 32866 704602 33102 704838
rect 32546 704282 32782 704518
rect 32866 704282 33102 704518
rect 32546 687218 32782 687454
rect 32866 687218 33102 687454
rect 32546 686898 32782 687134
rect 32866 686898 33102 687134
rect 38586 711322 38822 711558
rect 38906 711322 39142 711558
rect 38586 711002 38822 711238
rect 38906 711002 39142 711238
rect 33466 698378 33702 698614
rect 33786 698378 34022 698614
rect 33466 698058 33702 698294
rect 33786 698058 34022 698294
rect 33466 662378 33702 662614
rect 33786 662378 34022 662614
rect 33466 662058 33702 662294
rect 33786 662058 34022 662294
rect 34866 709402 35102 709638
rect 35186 709402 35422 709638
rect 34866 709082 35102 709318
rect 35186 709082 35422 709318
rect 34866 676658 35102 676894
rect 35186 676658 35422 676894
rect 34866 676338 35102 676574
rect 35186 676338 35422 676574
rect 36266 706522 36502 706758
rect 36586 706522 36822 706758
rect 36266 706202 36502 706438
rect 36586 706202 36822 706438
rect 36266 690938 36502 691174
rect 36586 690938 36822 691174
rect 36266 690618 36502 690854
rect 36586 690618 36822 690854
rect 37666 705562 37902 705798
rect 37986 705562 38222 705798
rect 37666 705242 37902 705478
rect 37986 705242 38222 705478
rect 37666 669218 37902 669454
rect 37986 669218 38222 669454
rect 37666 668898 37902 669134
rect 37986 668898 38222 669134
rect 43706 710362 43942 710598
rect 44026 710362 44262 710598
rect 43706 710042 43942 710278
rect 44026 710042 44262 710278
rect 38586 680378 38822 680614
rect 38906 680378 39142 680614
rect 38586 680058 38822 680294
rect 38906 680058 39142 680294
rect 39986 708442 40222 708678
rect 40306 708442 40542 708678
rect 39986 708122 40222 708358
rect 40306 708122 40542 708358
rect 39986 694658 40222 694894
rect 40306 694658 40542 694894
rect 39986 694338 40222 694574
rect 40306 694338 40542 694574
rect 39986 658658 40222 658894
rect 40306 658658 40542 658894
rect 39986 658338 40222 658574
rect 40306 658338 40542 658574
rect 41386 707482 41622 707718
rect 41706 707482 41942 707718
rect 41386 707162 41622 707398
rect 41706 707162 41942 707398
rect 41386 672938 41622 673174
rect 41706 672938 41942 673174
rect 41386 672618 41622 672854
rect 41706 672618 41942 672854
rect 42786 704602 43022 704838
rect 43106 704602 43342 704838
rect 42786 704282 43022 704518
rect 43106 704282 43342 704518
rect 42786 687218 43022 687454
rect 43106 687218 43342 687454
rect 42786 686898 43022 687134
rect 43106 686898 43342 687134
rect 48826 711322 49062 711558
rect 49146 711322 49382 711558
rect 48826 711002 49062 711238
rect 49146 711002 49382 711238
rect 43706 698378 43942 698614
rect 44026 698378 44262 698614
rect 43706 698058 43942 698294
rect 44026 698058 44262 698294
rect 43706 662378 43942 662614
rect 44026 662378 44262 662614
rect 43706 662058 43942 662294
rect 44026 662058 44262 662294
rect 45106 709402 45342 709638
rect 45426 709402 45662 709638
rect 45106 709082 45342 709318
rect 45426 709082 45662 709318
rect 45106 676658 45342 676894
rect 45426 676658 45662 676894
rect 45106 676338 45342 676574
rect 45426 676338 45662 676574
rect 46506 706522 46742 706758
rect 46826 706522 47062 706758
rect 46506 706202 46742 706438
rect 46826 706202 47062 706438
rect 46506 690938 46742 691174
rect 46826 690938 47062 691174
rect 46506 690618 46742 690854
rect 46826 690618 47062 690854
rect 47906 705562 48142 705798
rect 48226 705562 48462 705798
rect 47906 705242 48142 705478
rect 48226 705242 48462 705478
rect 47906 669218 48142 669454
rect 48226 669218 48462 669454
rect 47906 668898 48142 669134
rect 48226 668898 48462 669134
rect 53946 710362 54182 710598
rect 54266 710362 54502 710598
rect 53946 710042 54182 710278
rect 54266 710042 54502 710278
rect 48826 680378 49062 680614
rect 49146 680378 49382 680614
rect 48826 680058 49062 680294
rect 49146 680058 49382 680294
rect 50226 708442 50462 708678
rect 50546 708442 50782 708678
rect 50226 708122 50462 708358
rect 50546 708122 50782 708358
rect 50226 694658 50462 694894
rect 50546 694658 50782 694894
rect 50226 694338 50462 694574
rect 50546 694338 50782 694574
rect 50226 658658 50462 658894
rect 50546 658658 50782 658894
rect 50226 658338 50462 658574
rect 50546 658338 50782 658574
rect 51626 707482 51862 707718
rect 51946 707482 52182 707718
rect 51626 707162 51862 707398
rect 51946 707162 52182 707398
rect 51626 672938 51862 673174
rect 51946 672938 52182 673174
rect 51626 672618 51862 672854
rect 51946 672618 52182 672854
rect 53026 704602 53262 704838
rect 53346 704602 53582 704838
rect 53026 704282 53262 704518
rect 53346 704282 53582 704518
rect 53026 687218 53262 687454
rect 53346 687218 53582 687454
rect 53026 686898 53262 687134
rect 53346 686898 53582 687134
rect 59066 711322 59302 711558
rect 59386 711322 59622 711558
rect 59066 711002 59302 711238
rect 59386 711002 59622 711238
rect 53946 698378 54182 698614
rect 54266 698378 54502 698614
rect 53946 698058 54182 698294
rect 54266 698058 54502 698294
rect 53946 662378 54182 662614
rect 54266 662378 54502 662614
rect 53946 662058 54182 662294
rect 54266 662058 54502 662294
rect 55346 709402 55582 709638
rect 55666 709402 55902 709638
rect 55346 709082 55582 709318
rect 55666 709082 55902 709318
rect 55346 676658 55582 676894
rect 55666 676658 55902 676894
rect 55346 676338 55582 676574
rect 55666 676338 55902 676574
rect 56746 706522 56982 706758
rect 57066 706522 57302 706758
rect 56746 706202 56982 706438
rect 57066 706202 57302 706438
rect 56746 690938 56982 691174
rect 57066 690938 57302 691174
rect 56746 690618 56982 690854
rect 57066 690618 57302 690854
rect 58146 705562 58382 705798
rect 58466 705562 58702 705798
rect 58146 705242 58382 705478
rect 58466 705242 58702 705478
rect 58146 669218 58382 669454
rect 58466 669218 58702 669454
rect 58146 668898 58382 669134
rect 58466 668898 58702 669134
rect 64186 710362 64422 710598
rect 64506 710362 64742 710598
rect 64186 710042 64422 710278
rect 64506 710042 64742 710278
rect 59066 680378 59302 680614
rect 59386 680378 59622 680614
rect 59066 680058 59302 680294
rect 59386 680058 59622 680294
rect 60466 708442 60702 708678
rect 60786 708442 61022 708678
rect 60466 708122 60702 708358
rect 60786 708122 61022 708358
rect 60466 694658 60702 694894
rect 60786 694658 61022 694894
rect 60466 694338 60702 694574
rect 60786 694338 61022 694574
rect 60466 658658 60702 658894
rect 60786 658658 61022 658894
rect 60466 658338 60702 658574
rect 60786 658338 61022 658574
rect 61866 707482 62102 707718
rect 62186 707482 62422 707718
rect 61866 707162 62102 707398
rect 62186 707162 62422 707398
rect 61866 672938 62102 673174
rect 62186 672938 62422 673174
rect 61866 672618 62102 672854
rect 62186 672618 62422 672854
rect 63266 704602 63502 704838
rect 63586 704602 63822 704838
rect 63266 704282 63502 704518
rect 63586 704282 63822 704518
rect 63266 687218 63502 687454
rect 63586 687218 63822 687454
rect 63266 686898 63502 687134
rect 63586 686898 63822 687134
rect 69306 711322 69542 711558
rect 69626 711322 69862 711558
rect 69306 711002 69542 711238
rect 69626 711002 69862 711238
rect 64186 698378 64422 698614
rect 64506 698378 64742 698614
rect 64186 698058 64422 698294
rect 64506 698058 64742 698294
rect 64186 662378 64422 662614
rect 64506 662378 64742 662614
rect 64186 662058 64422 662294
rect 64506 662058 64742 662294
rect 65586 709402 65822 709638
rect 65906 709402 66142 709638
rect 65586 709082 65822 709318
rect 65906 709082 66142 709318
rect 65586 676658 65822 676894
rect 65906 676658 66142 676894
rect 65586 676338 65822 676574
rect 65906 676338 66142 676574
rect 66986 706522 67222 706758
rect 67306 706522 67542 706758
rect 66986 706202 67222 706438
rect 67306 706202 67542 706438
rect 66986 690938 67222 691174
rect 67306 690938 67542 691174
rect 66986 690618 67222 690854
rect 67306 690618 67542 690854
rect 68386 705562 68622 705798
rect 68706 705562 68942 705798
rect 68386 705242 68622 705478
rect 68706 705242 68942 705478
rect 68386 669218 68622 669454
rect 68706 669218 68942 669454
rect 68386 668898 68622 669134
rect 68706 668898 68942 669134
rect 74426 710362 74662 710598
rect 74746 710362 74982 710598
rect 74426 710042 74662 710278
rect 74746 710042 74982 710278
rect 69306 680378 69542 680614
rect 69626 680378 69862 680614
rect 69306 680058 69542 680294
rect 69626 680058 69862 680294
rect 70706 708442 70942 708678
rect 71026 708442 71262 708678
rect 70706 708122 70942 708358
rect 71026 708122 71262 708358
rect 70706 694658 70942 694894
rect 71026 694658 71262 694894
rect 70706 694338 70942 694574
rect 71026 694338 71262 694574
rect 70706 658658 70942 658894
rect 71026 658658 71262 658894
rect 70706 658338 70942 658574
rect 71026 658338 71262 658574
rect 72106 707482 72342 707718
rect 72426 707482 72662 707718
rect 72106 707162 72342 707398
rect 72426 707162 72662 707398
rect 72106 672938 72342 673174
rect 72426 672938 72662 673174
rect 72106 672618 72342 672854
rect 72426 672618 72662 672854
rect 73506 704602 73742 704838
rect 73826 704602 74062 704838
rect 73506 704282 73742 704518
rect 73826 704282 74062 704518
rect 73506 687218 73742 687454
rect 73826 687218 74062 687454
rect 73506 686898 73742 687134
rect 73826 686898 74062 687134
rect 79546 711322 79782 711558
rect 79866 711322 80102 711558
rect 79546 711002 79782 711238
rect 79866 711002 80102 711238
rect 74426 698378 74662 698614
rect 74746 698378 74982 698614
rect 74426 698058 74662 698294
rect 74746 698058 74982 698294
rect 74426 662378 74662 662614
rect 74746 662378 74982 662614
rect 74426 662058 74662 662294
rect 74746 662058 74982 662294
rect 75826 709402 76062 709638
rect 76146 709402 76382 709638
rect 75826 709082 76062 709318
rect 76146 709082 76382 709318
rect 75826 676658 76062 676894
rect 76146 676658 76382 676894
rect 75826 676338 76062 676574
rect 76146 676338 76382 676574
rect 77226 706522 77462 706758
rect 77546 706522 77782 706758
rect 77226 706202 77462 706438
rect 77546 706202 77782 706438
rect 77226 690938 77462 691174
rect 77546 690938 77782 691174
rect 77226 690618 77462 690854
rect 77546 690618 77782 690854
rect 78626 705562 78862 705798
rect 78946 705562 79182 705798
rect 78626 705242 78862 705478
rect 78946 705242 79182 705478
rect 78626 669218 78862 669454
rect 78946 669218 79182 669454
rect 78626 668898 78862 669134
rect 78946 668898 79182 669134
rect 84666 710362 84902 710598
rect 84986 710362 85222 710598
rect 84666 710042 84902 710278
rect 84986 710042 85222 710278
rect 79546 680378 79782 680614
rect 79866 680378 80102 680614
rect 79546 680058 79782 680294
rect 79866 680058 80102 680294
rect 80946 708442 81182 708678
rect 81266 708442 81502 708678
rect 80946 708122 81182 708358
rect 81266 708122 81502 708358
rect 80946 694658 81182 694894
rect 81266 694658 81502 694894
rect 80946 694338 81182 694574
rect 81266 694338 81502 694574
rect 80946 658658 81182 658894
rect 81266 658658 81502 658894
rect 80946 658338 81182 658574
rect 81266 658338 81502 658574
rect 82346 707482 82582 707718
rect 82666 707482 82902 707718
rect 82346 707162 82582 707398
rect 82666 707162 82902 707398
rect 82346 672938 82582 673174
rect 82666 672938 82902 673174
rect 82346 672618 82582 672854
rect 82666 672618 82902 672854
rect 83746 704602 83982 704838
rect 84066 704602 84302 704838
rect 83746 704282 83982 704518
rect 84066 704282 84302 704518
rect 83746 687218 83982 687454
rect 84066 687218 84302 687454
rect 83746 686898 83982 687134
rect 84066 686898 84302 687134
rect 89786 711322 90022 711558
rect 90106 711322 90342 711558
rect 89786 711002 90022 711238
rect 90106 711002 90342 711238
rect 84666 698378 84902 698614
rect 84986 698378 85222 698614
rect 84666 698058 84902 698294
rect 84986 698058 85222 698294
rect 84666 662378 84902 662614
rect 84986 662378 85222 662614
rect 84666 662058 84902 662294
rect 84986 662058 85222 662294
rect 86066 709402 86302 709638
rect 86386 709402 86622 709638
rect 86066 709082 86302 709318
rect 86386 709082 86622 709318
rect 86066 676658 86302 676894
rect 86386 676658 86622 676894
rect 86066 676338 86302 676574
rect 86386 676338 86622 676574
rect 87466 706522 87702 706758
rect 87786 706522 88022 706758
rect 87466 706202 87702 706438
rect 87786 706202 88022 706438
rect 87466 690938 87702 691174
rect 87786 690938 88022 691174
rect 87466 690618 87702 690854
rect 87786 690618 88022 690854
rect 88866 705562 89102 705798
rect 89186 705562 89422 705798
rect 88866 705242 89102 705478
rect 89186 705242 89422 705478
rect 88866 669218 89102 669454
rect 89186 669218 89422 669454
rect 88866 668898 89102 669134
rect 89186 668898 89422 669134
rect 94906 710362 95142 710598
rect 95226 710362 95462 710598
rect 94906 710042 95142 710278
rect 95226 710042 95462 710278
rect 89786 680378 90022 680614
rect 90106 680378 90342 680614
rect 89786 680058 90022 680294
rect 90106 680058 90342 680294
rect 91186 708442 91422 708678
rect 91506 708442 91742 708678
rect 91186 708122 91422 708358
rect 91506 708122 91742 708358
rect 91186 694658 91422 694894
rect 91506 694658 91742 694894
rect 91186 694338 91422 694574
rect 91506 694338 91742 694574
rect 91186 658658 91422 658894
rect 91506 658658 91742 658894
rect 91186 658338 91422 658574
rect 91506 658338 91742 658574
rect 92586 707482 92822 707718
rect 92906 707482 93142 707718
rect 92586 707162 92822 707398
rect 92906 707162 93142 707398
rect 92586 672938 92822 673174
rect 92906 672938 93142 673174
rect 92586 672618 92822 672854
rect 92906 672618 93142 672854
rect 93986 704602 94222 704838
rect 94306 704602 94542 704838
rect 93986 704282 94222 704518
rect 94306 704282 94542 704518
rect 93986 687218 94222 687454
rect 94306 687218 94542 687454
rect 93986 686898 94222 687134
rect 94306 686898 94542 687134
rect 100026 711322 100262 711558
rect 100346 711322 100582 711558
rect 100026 711002 100262 711238
rect 100346 711002 100582 711238
rect 94906 698378 95142 698614
rect 95226 698378 95462 698614
rect 94906 698058 95142 698294
rect 95226 698058 95462 698294
rect 94906 662378 95142 662614
rect 95226 662378 95462 662614
rect 94906 662058 95142 662294
rect 95226 662058 95462 662294
rect 96306 709402 96542 709638
rect 96626 709402 96862 709638
rect 96306 709082 96542 709318
rect 96626 709082 96862 709318
rect 96306 676658 96542 676894
rect 96626 676658 96862 676894
rect 96306 676338 96542 676574
rect 96626 676338 96862 676574
rect 97706 706522 97942 706758
rect 98026 706522 98262 706758
rect 97706 706202 97942 706438
rect 98026 706202 98262 706438
rect 97706 690938 97942 691174
rect 98026 690938 98262 691174
rect 97706 690618 97942 690854
rect 98026 690618 98262 690854
rect 99106 705562 99342 705798
rect 99426 705562 99662 705798
rect 99106 705242 99342 705478
rect 99426 705242 99662 705478
rect 99106 669218 99342 669454
rect 99426 669218 99662 669454
rect 99106 668898 99342 669134
rect 99426 668898 99662 669134
rect 105146 710362 105382 710598
rect 105466 710362 105702 710598
rect 105146 710042 105382 710278
rect 105466 710042 105702 710278
rect 100026 680378 100262 680614
rect 100346 680378 100582 680614
rect 100026 680058 100262 680294
rect 100346 680058 100582 680294
rect 101426 708442 101662 708678
rect 101746 708442 101982 708678
rect 101426 708122 101662 708358
rect 101746 708122 101982 708358
rect 101426 694658 101662 694894
rect 101746 694658 101982 694894
rect 101426 694338 101662 694574
rect 101746 694338 101982 694574
rect 101426 658658 101662 658894
rect 101746 658658 101982 658894
rect 101426 658338 101662 658574
rect 101746 658338 101982 658574
rect 102826 707482 103062 707718
rect 103146 707482 103382 707718
rect 102826 707162 103062 707398
rect 103146 707162 103382 707398
rect 102826 672938 103062 673174
rect 103146 672938 103382 673174
rect 102826 672618 103062 672854
rect 103146 672618 103382 672854
rect 104226 704602 104462 704838
rect 104546 704602 104782 704838
rect 104226 704282 104462 704518
rect 104546 704282 104782 704518
rect 104226 687218 104462 687454
rect 104546 687218 104782 687454
rect 104226 686898 104462 687134
rect 104546 686898 104782 687134
rect 110266 711322 110502 711558
rect 110586 711322 110822 711558
rect 110266 711002 110502 711238
rect 110586 711002 110822 711238
rect 105146 698378 105382 698614
rect 105466 698378 105702 698614
rect 105146 698058 105382 698294
rect 105466 698058 105702 698294
rect 105146 662378 105382 662614
rect 105466 662378 105702 662614
rect 105146 662058 105382 662294
rect 105466 662058 105702 662294
rect 106546 709402 106782 709638
rect 106866 709402 107102 709638
rect 106546 709082 106782 709318
rect 106866 709082 107102 709318
rect 106546 676658 106782 676894
rect 106866 676658 107102 676894
rect 106546 676338 106782 676574
rect 106866 676338 107102 676574
rect 107946 706522 108182 706758
rect 108266 706522 108502 706758
rect 107946 706202 108182 706438
rect 108266 706202 108502 706438
rect 107946 690938 108182 691174
rect 108266 690938 108502 691174
rect 107946 690618 108182 690854
rect 108266 690618 108502 690854
rect 109346 705562 109582 705798
rect 109666 705562 109902 705798
rect 109346 705242 109582 705478
rect 109666 705242 109902 705478
rect 109346 669218 109582 669454
rect 109666 669218 109902 669454
rect 109346 668898 109582 669134
rect 109666 668898 109902 669134
rect 115386 710362 115622 710598
rect 115706 710362 115942 710598
rect 115386 710042 115622 710278
rect 115706 710042 115942 710278
rect 110266 680378 110502 680614
rect 110586 680378 110822 680614
rect 110266 680058 110502 680294
rect 110586 680058 110822 680294
rect 111666 708442 111902 708678
rect 111986 708442 112222 708678
rect 111666 708122 111902 708358
rect 111986 708122 112222 708358
rect 111666 694658 111902 694894
rect 111986 694658 112222 694894
rect 111666 694338 111902 694574
rect 111986 694338 112222 694574
rect 111666 658658 111902 658894
rect 111986 658658 112222 658894
rect 111666 658338 111902 658574
rect 111986 658338 112222 658574
rect 113066 707482 113302 707718
rect 113386 707482 113622 707718
rect 113066 707162 113302 707398
rect 113386 707162 113622 707398
rect 113066 672938 113302 673174
rect 113386 672938 113622 673174
rect 113066 672618 113302 672854
rect 113386 672618 113622 672854
rect 114466 704602 114702 704838
rect 114786 704602 115022 704838
rect 114466 704282 114702 704518
rect 114786 704282 115022 704518
rect 114466 687218 114702 687454
rect 114786 687218 115022 687454
rect 114466 686898 114702 687134
rect 114786 686898 115022 687134
rect 120506 711322 120742 711558
rect 120826 711322 121062 711558
rect 120506 711002 120742 711238
rect 120826 711002 121062 711238
rect 115386 698378 115622 698614
rect 115706 698378 115942 698614
rect 115386 698058 115622 698294
rect 115706 698058 115942 698294
rect 115386 662378 115622 662614
rect 115706 662378 115942 662614
rect 115386 662058 115622 662294
rect 115706 662058 115942 662294
rect 116786 709402 117022 709638
rect 117106 709402 117342 709638
rect 116786 709082 117022 709318
rect 117106 709082 117342 709318
rect 116786 676658 117022 676894
rect 117106 676658 117342 676894
rect 116786 676338 117022 676574
rect 117106 676338 117342 676574
rect 118186 706522 118422 706758
rect 118506 706522 118742 706758
rect 118186 706202 118422 706438
rect 118506 706202 118742 706438
rect 118186 690938 118422 691174
rect 118506 690938 118742 691174
rect 118186 690618 118422 690854
rect 118506 690618 118742 690854
rect 119586 705562 119822 705798
rect 119906 705562 120142 705798
rect 119586 705242 119822 705478
rect 119906 705242 120142 705478
rect 119586 669218 119822 669454
rect 119906 669218 120142 669454
rect 119586 668898 119822 669134
rect 119906 668898 120142 669134
rect 125626 710362 125862 710598
rect 125946 710362 126182 710598
rect 125626 710042 125862 710278
rect 125946 710042 126182 710278
rect 120506 680378 120742 680614
rect 120826 680378 121062 680614
rect 120506 680058 120742 680294
rect 120826 680058 121062 680294
rect 121906 708442 122142 708678
rect 122226 708442 122462 708678
rect 121906 708122 122142 708358
rect 122226 708122 122462 708358
rect 121906 694658 122142 694894
rect 122226 694658 122462 694894
rect 121906 694338 122142 694574
rect 122226 694338 122462 694574
rect 121906 658658 122142 658894
rect 122226 658658 122462 658894
rect 121906 658338 122142 658574
rect 122226 658338 122462 658574
rect 123306 707482 123542 707718
rect 123626 707482 123862 707718
rect 123306 707162 123542 707398
rect 123626 707162 123862 707398
rect 123306 672938 123542 673174
rect 123626 672938 123862 673174
rect 123306 672618 123542 672854
rect 123626 672618 123862 672854
rect 124706 704602 124942 704838
rect 125026 704602 125262 704838
rect 124706 704282 124942 704518
rect 125026 704282 125262 704518
rect 124706 687218 124942 687454
rect 125026 687218 125262 687454
rect 124706 686898 124942 687134
rect 125026 686898 125262 687134
rect 130746 711322 130982 711558
rect 131066 711322 131302 711558
rect 130746 711002 130982 711238
rect 131066 711002 131302 711238
rect 125626 698378 125862 698614
rect 125946 698378 126182 698614
rect 125626 698058 125862 698294
rect 125946 698058 126182 698294
rect 125626 662378 125862 662614
rect 125946 662378 126182 662614
rect 125626 662058 125862 662294
rect 125946 662058 126182 662294
rect 127026 709402 127262 709638
rect 127346 709402 127582 709638
rect 127026 709082 127262 709318
rect 127346 709082 127582 709318
rect 127026 676658 127262 676894
rect 127346 676658 127582 676894
rect 127026 676338 127262 676574
rect 127346 676338 127582 676574
rect 128426 706522 128662 706758
rect 128746 706522 128982 706758
rect 128426 706202 128662 706438
rect 128746 706202 128982 706438
rect 128426 690938 128662 691174
rect 128746 690938 128982 691174
rect 128426 690618 128662 690854
rect 128746 690618 128982 690854
rect 129826 705562 130062 705798
rect 130146 705562 130382 705798
rect 129826 705242 130062 705478
rect 130146 705242 130382 705478
rect 129826 669218 130062 669454
rect 130146 669218 130382 669454
rect 129826 668898 130062 669134
rect 130146 668898 130382 669134
rect 135866 710362 136102 710598
rect 136186 710362 136422 710598
rect 135866 710042 136102 710278
rect 136186 710042 136422 710278
rect 130746 680378 130982 680614
rect 131066 680378 131302 680614
rect 130746 680058 130982 680294
rect 131066 680058 131302 680294
rect 132146 708442 132382 708678
rect 132466 708442 132702 708678
rect 132146 708122 132382 708358
rect 132466 708122 132702 708358
rect 132146 694658 132382 694894
rect 132466 694658 132702 694894
rect 132146 694338 132382 694574
rect 132466 694338 132702 694574
rect 132146 658658 132382 658894
rect 132466 658658 132702 658894
rect 132146 658338 132382 658574
rect 132466 658338 132702 658574
rect 133546 707482 133782 707718
rect 133866 707482 134102 707718
rect 133546 707162 133782 707398
rect 133866 707162 134102 707398
rect 133546 672938 133782 673174
rect 133866 672938 134102 673174
rect 133546 672618 133782 672854
rect 133866 672618 134102 672854
rect 134946 704602 135182 704838
rect 135266 704602 135502 704838
rect 134946 704282 135182 704518
rect 135266 704282 135502 704518
rect 134946 687218 135182 687454
rect 135266 687218 135502 687454
rect 134946 686898 135182 687134
rect 135266 686898 135502 687134
rect 140986 711322 141222 711558
rect 141306 711322 141542 711558
rect 140986 711002 141222 711238
rect 141306 711002 141542 711238
rect 135866 698378 136102 698614
rect 136186 698378 136422 698614
rect 135866 698058 136102 698294
rect 136186 698058 136422 698294
rect 135866 662378 136102 662614
rect 136186 662378 136422 662614
rect 135866 662058 136102 662294
rect 136186 662058 136422 662294
rect 137266 709402 137502 709638
rect 137586 709402 137822 709638
rect 137266 709082 137502 709318
rect 137586 709082 137822 709318
rect 137266 676658 137502 676894
rect 137586 676658 137822 676894
rect 137266 676338 137502 676574
rect 137586 676338 137822 676574
rect 138666 706522 138902 706758
rect 138986 706522 139222 706758
rect 138666 706202 138902 706438
rect 138986 706202 139222 706438
rect 138666 690938 138902 691174
rect 138986 690938 139222 691174
rect 138666 690618 138902 690854
rect 138986 690618 139222 690854
rect 140066 705562 140302 705798
rect 140386 705562 140622 705798
rect 140066 705242 140302 705478
rect 140386 705242 140622 705478
rect 140066 669218 140302 669454
rect 140386 669218 140622 669454
rect 140066 668898 140302 669134
rect 140386 668898 140622 669134
rect 146106 710362 146342 710598
rect 146426 710362 146662 710598
rect 146106 710042 146342 710278
rect 146426 710042 146662 710278
rect 140986 680378 141222 680614
rect 141306 680378 141542 680614
rect 140986 680058 141222 680294
rect 141306 680058 141542 680294
rect 142386 708442 142622 708678
rect 142706 708442 142942 708678
rect 142386 708122 142622 708358
rect 142706 708122 142942 708358
rect 142386 694658 142622 694894
rect 142706 694658 142942 694894
rect 142386 694338 142622 694574
rect 142706 694338 142942 694574
rect 142386 658658 142622 658894
rect 142706 658658 142942 658894
rect 142386 658338 142622 658574
rect 142706 658338 142942 658574
rect 143786 707482 144022 707718
rect 144106 707482 144342 707718
rect 143786 707162 144022 707398
rect 144106 707162 144342 707398
rect 143786 672938 144022 673174
rect 144106 672938 144342 673174
rect 143786 672618 144022 672854
rect 144106 672618 144342 672854
rect 145186 704602 145422 704838
rect 145506 704602 145742 704838
rect 145186 704282 145422 704518
rect 145506 704282 145742 704518
rect 145186 687218 145422 687454
rect 145506 687218 145742 687454
rect 145186 686898 145422 687134
rect 145506 686898 145742 687134
rect 151226 711322 151462 711558
rect 151546 711322 151782 711558
rect 151226 711002 151462 711238
rect 151546 711002 151782 711238
rect 146106 698378 146342 698614
rect 146426 698378 146662 698614
rect 146106 698058 146342 698294
rect 146426 698058 146662 698294
rect 146106 662378 146342 662614
rect 146426 662378 146662 662614
rect 146106 662058 146342 662294
rect 146426 662058 146662 662294
rect 147506 709402 147742 709638
rect 147826 709402 148062 709638
rect 147506 709082 147742 709318
rect 147826 709082 148062 709318
rect 147506 676658 147742 676894
rect 147826 676658 148062 676894
rect 147506 676338 147742 676574
rect 147826 676338 148062 676574
rect 148906 706522 149142 706758
rect 149226 706522 149462 706758
rect 148906 706202 149142 706438
rect 149226 706202 149462 706438
rect 148906 690938 149142 691174
rect 149226 690938 149462 691174
rect 148906 690618 149142 690854
rect 149226 690618 149462 690854
rect 150306 705562 150542 705798
rect 150626 705562 150862 705798
rect 150306 705242 150542 705478
rect 150626 705242 150862 705478
rect 150306 669218 150542 669454
rect 150626 669218 150862 669454
rect 150306 668898 150542 669134
rect 150626 668898 150862 669134
rect 156346 710362 156582 710598
rect 156666 710362 156902 710598
rect 156346 710042 156582 710278
rect 156666 710042 156902 710278
rect 151226 680378 151462 680614
rect 151546 680378 151782 680614
rect 151226 680058 151462 680294
rect 151546 680058 151782 680294
rect 152626 708442 152862 708678
rect 152946 708442 153182 708678
rect 152626 708122 152862 708358
rect 152946 708122 153182 708358
rect 152626 694658 152862 694894
rect 152946 694658 153182 694894
rect 152626 694338 152862 694574
rect 152946 694338 153182 694574
rect 152626 658658 152862 658894
rect 152946 658658 153182 658894
rect 152626 658338 152862 658574
rect 152946 658338 153182 658574
rect 154026 707482 154262 707718
rect 154346 707482 154582 707718
rect 154026 707162 154262 707398
rect 154346 707162 154582 707398
rect 154026 672938 154262 673174
rect 154346 672938 154582 673174
rect 154026 672618 154262 672854
rect 154346 672618 154582 672854
rect 155426 704602 155662 704838
rect 155746 704602 155982 704838
rect 155426 704282 155662 704518
rect 155746 704282 155982 704518
rect 155426 687218 155662 687454
rect 155746 687218 155982 687454
rect 155426 686898 155662 687134
rect 155746 686898 155982 687134
rect 161466 711322 161702 711558
rect 161786 711322 162022 711558
rect 161466 711002 161702 711238
rect 161786 711002 162022 711238
rect 156346 698378 156582 698614
rect 156666 698378 156902 698614
rect 156346 698058 156582 698294
rect 156666 698058 156902 698294
rect 156346 662378 156582 662614
rect 156666 662378 156902 662614
rect 156346 662058 156582 662294
rect 156666 662058 156902 662294
rect 157746 709402 157982 709638
rect 158066 709402 158302 709638
rect 157746 709082 157982 709318
rect 158066 709082 158302 709318
rect 157746 676658 157982 676894
rect 158066 676658 158302 676894
rect 157746 676338 157982 676574
rect 158066 676338 158302 676574
rect 159146 706522 159382 706758
rect 159466 706522 159702 706758
rect 159146 706202 159382 706438
rect 159466 706202 159702 706438
rect 159146 690938 159382 691174
rect 159466 690938 159702 691174
rect 159146 690618 159382 690854
rect 159466 690618 159702 690854
rect 160546 705562 160782 705798
rect 160866 705562 161102 705798
rect 160546 705242 160782 705478
rect 160866 705242 161102 705478
rect 160546 669218 160782 669454
rect 160866 669218 161102 669454
rect 160546 668898 160782 669134
rect 160866 668898 161102 669134
rect 166586 710362 166822 710598
rect 166906 710362 167142 710598
rect 166586 710042 166822 710278
rect 166906 710042 167142 710278
rect 161466 680378 161702 680614
rect 161786 680378 162022 680614
rect 161466 680058 161702 680294
rect 161786 680058 162022 680294
rect 162866 708442 163102 708678
rect 163186 708442 163422 708678
rect 162866 708122 163102 708358
rect 163186 708122 163422 708358
rect 162866 694658 163102 694894
rect 163186 694658 163422 694894
rect 162866 694338 163102 694574
rect 163186 694338 163422 694574
rect 162866 658658 163102 658894
rect 163186 658658 163422 658894
rect 162866 658338 163102 658574
rect 163186 658338 163422 658574
rect 164266 707482 164502 707718
rect 164586 707482 164822 707718
rect 164266 707162 164502 707398
rect 164586 707162 164822 707398
rect 164266 672938 164502 673174
rect 164586 672938 164822 673174
rect 164266 672618 164502 672854
rect 164586 672618 164822 672854
rect 165666 704602 165902 704838
rect 165986 704602 166222 704838
rect 165666 704282 165902 704518
rect 165986 704282 166222 704518
rect 165666 687218 165902 687454
rect 165986 687218 166222 687454
rect 165666 686898 165902 687134
rect 165986 686898 166222 687134
rect 171706 711322 171942 711558
rect 172026 711322 172262 711558
rect 171706 711002 171942 711238
rect 172026 711002 172262 711238
rect 166586 698378 166822 698614
rect 166906 698378 167142 698614
rect 166586 698058 166822 698294
rect 166906 698058 167142 698294
rect 166586 662378 166822 662614
rect 166906 662378 167142 662614
rect 166586 662058 166822 662294
rect 166906 662058 167142 662294
rect 167986 709402 168222 709638
rect 168306 709402 168542 709638
rect 167986 709082 168222 709318
rect 168306 709082 168542 709318
rect 167986 676658 168222 676894
rect 168306 676658 168542 676894
rect 167986 676338 168222 676574
rect 168306 676338 168542 676574
rect 169386 706522 169622 706758
rect 169706 706522 169942 706758
rect 169386 706202 169622 706438
rect 169706 706202 169942 706438
rect 169386 690938 169622 691174
rect 169706 690938 169942 691174
rect 169386 690618 169622 690854
rect 169706 690618 169942 690854
rect 170786 705562 171022 705798
rect 171106 705562 171342 705798
rect 170786 705242 171022 705478
rect 171106 705242 171342 705478
rect 170786 669218 171022 669454
rect 171106 669218 171342 669454
rect 170786 668898 171022 669134
rect 171106 668898 171342 669134
rect 176826 710362 177062 710598
rect 177146 710362 177382 710598
rect 176826 710042 177062 710278
rect 177146 710042 177382 710278
rect 171706 680378 171942 680614
rect 172026 680378 172262 680614
rect 171706 680058 171942 680294
rect 172026 680058 172262 680294
rect 173106 708442 173342 708678
rect 173426 708442 173662 708678
rect 173106 708122 173342 708358
rect 173426 708122 173662 708358
rect 173106 694658 173342 694894
rect 173426 694658 173662 694894
rect 173106 694338 173342 694574
rect 173426 694338 173662 694574
rect 173106 658658 173342 658894
rect 173426 658658 173662 658894
rect 173106 658338 173342 658574
rect 173426 658338 173662 658574
rect 174506 707482 174742 707718
rect 174826 707482 175062 707718
rect 174506 707162 174742 707398
rect 174826 707162 175062 707398
rect 174506 672938 174742 673174
rect 174826 672938 175062 673174
rect 174506 672618 174742 672854
rect 174826 672618 175062 672854
rect 175906 704602 176142 704838
rect 176226 704602 176462 704838
rect 175906 704282 176142 704518
rect 176226 704282 176462 704518
rect 175906 687218 176142 687454
rect 176226 687218 176462 687454
rect 175906 686898 176142 687134
rect 176226 686898 176462 687134
rect 181946 711322 182182 711558
rect 182266 711322 182502 711558
rect 181946 711002 182182 711238
rect 182266 711002 182502 711238
rect 176826 698378 177062 698614
rect 177146 698378 177382 698614
rect 176826 698058 177062 698294
rect 177146 698058 177382 698294
rect 176826 662378 177062 662614
rect 177146 662378 177382 662614
rect 176826 662058 177062 662294
rect 177146 662058 177382 662294
rect 178226 709402 178462 709638
rect 178546 709402 178782 709638
rect 178226 709082 178462 709318
rect 178546 709082 178782 709318
rect 178226 676658 178462 676894
rect 178546 676658 178782 676894
rect 178226 676338 178462 676574
rect 178546 676338 178782 676574
rect 179626 706522 179862 706758
rect 179946 706522 180182 706758
rect 179626 706202 179862 706438
rect 179946 706202 180182 706438
rect 179626 690938 179862 691174
rect 179946 690938 180182 691174
rect 179626 690618 179862 690854
rect 179946 690618 180182 690854
rect 181026 705562 181262 705798
rect 181346 705562 181582 705798
rect 181026 705242 181262 705478
rect 181346 705242 181582 705478
rect 181026 669218 181262 669454
rect 181346 669218 181582 669454
rect 181026 668898 181262 669134
rect 181346 668898 181582 669134
rect 187066 710362 187302 710598
rect 187386 710362 187622 710598
rect 187066 710042 187302 710278
rect 187386 710042 187622 710278
rect 181946 680378 182182 680614
rect 182266 680378 182502 680614
rect 181946 680058 182182 680294
rect 182266 680058 182502 680294
rect 183346 708442 183582 708678
rect 183666 708442 183902 708678
rect 183346 708122 183582 708358
rect 183666 708122 183902 708358
rect 183346 694658 183582 694894
rect 183666 694658 183902 694894
rect 183346 694338 183582 694574
rect 183666 694338 183902 694574
rect 183346 658658 183582 658894
rect 183666 658658 183902 658894
rect 183346 658338 183582 658574
rect 183666 658338 183902 658574
rect 184746 707482 184982 707718
rect 185066 707482 185302 707718
rect 184746 707162 184982 707398
rect 185066 707162 185302 707398
rect 184746 672938 184982 673174
rect 185066 672938 185302 673174
rect 184746 672618 184982 672854
rect 185066 672618 185302 672854
rect 186146 704602 186382 704838
rect 186466 704602 186702 704838
rect 186146 704282 186382 704518
rect 186466 704282 186702 704518
rect 186146 687218 186382 687454
rect 186466 687218 186702 687454
rect 186146 686898 186382 687134
rect 186466 686898 186702 687134
rect 192186 711322 192422 711558
rect 192506 711322 192742 711558
rect 192186 711002 192422 711238
rect 192506 711002 192742 711238
rect 187066 698378 187302 698614
rect 187386 698378 187622 698614
rect 187066 698058 187302 698294
rect 187386 698058 187622 698294
rect 187066 662378 187302 662614
rect 187386 662378 187622 662614
rect 187066 662058 187302 662294
rect 187386 662058 187622 662294
rect 188466 709402 188702 709638
rect 188786 709402 189022 709638
rect 188466 709082 188702 709318
rect 188786 709082 189022 709318
rect 188466 676658 188702 676894
rect 188786 676658 189022 676894
rect 188466 676338 188702 676574
rect 188786 676338 189022 676574
rect 189866 706522 190102 706758
rect 190186 706522 190422 706758
rect 189866 706202 190102 706438
rect 190186 706202 190422 706438
rect 189866 690938 190102 691174
rect 190186 690938 190422 691174
rect 189866 690618 190102 690854
rect 190186 690618 190422 690854
rect 191266 705562 191502 705798
rect 191586 705562 191822 705798
rect 191266 705242 191502 705478
rect 191586 705242 191822 705478
rect 191266 669218 191502 669454
rect 191586 669218 191822 669454
rect 191266 668898 191502 669134
rect 191586 668898 191822 669134
rect 197306 710362 197542 710598
rect 197626 710362 197862 710598
rect 197306 710042 197542 710278
rect 197626 710042 197862 710278
rect 192186 680378 192422 680614
rect 192506 680378 192742 680614
rect 192186 680058 192422 680294
rect 192506 680058 192742 680294
rect 193586 708442 193822 708678
rect 193906 708442 194142 708678
rect 193586 708122 193822 708358
rect 193906 708122 194142 708358
rect 193586 694658 193822 694894
rect 193906 694658 194142 694894
rect 193586 694338 193822 694574
rect 193906 694338 194142 694574
rect 193586 658658 193822 658894
rect 193906 658658 194142 658894
rect 193586 658338 193822 658574
rect 193906 658338 194142 658574
rect 194986 707482 195222 707718
rect 195306 707482 195542 707718
rect 194986 707162 195222 707398
rect 195306 707162 195542 707398
rect 194986 672938 195222 673174
rect 195306 672938 195542 673174
rect 194986 672618 195222 672854
rect 195306 672618 195542 672854
rect 196386 704602 196622 704838
rect 196706 704602 196942 704838
rect 196386 704282 196622 704518
rect 196706 704282 196942 704518
rect 196386 687218 196622 687454
rect 196706 687218 196942 687454
rect 196386 686898 196622 687134
rect 196706 686898 196942 687134
rect 202426 711322 202662 711558
rect 202746 711322 202982 711558
rect 202426 711002 202662 711238
rect 202746 711002 202982 711238
rect 197306 698378 197542 698614
rect 197626 698378 197862 698614
rect 197306 698058 197542 698294
rect 197626 698058 197862 698294
rect 197306 662378 197542 662614
rect 197626 662378 197862 662614
rect 197306 662058 197542 662294
rect 197626 662058 197862 662294
rect 198706 709402 198942 709638
rect 199026 709402 199262 709638
rect 198706 709082 198942 709318
rect 199026 709082 199262 709318
rect 198706 676658 198942 676894
rect 199026 676658 199262 676894
rect 198706 676338 198942 676574
rect 199026 676338 199262 676574
rect 200106 706522 200342 706758
rect 200426 706522 200662 706758
rect 200106 706202 200342 706438
rect 200426 706202 200662 706438
rect 200106 690938 200342 691174
rect 200426 690938 200662 691174
rect 200106 690618 200342 690854
rect 200426 690618 200662 690854
rect 201506 705562 201742 705798
rect 201826 705562 202062 705798
rect 201506 705242 201742 705478
rect 201826 705242 202062 705478
rect 201506 669218 201742 669454
rect 201826 669218 202062 669454
rect 201506 668898 201742 669134
rect 201826 668898 202062 669134
rect 207546 710362 207782 710598
rect 207866 710362 208102 710598
rect 207546 710042 207782 710278
rect 207866 710042 208102 710278
rect 202426 680378 202662 680614
rect 202746 680378 202982 680614
rect 202426 680058 202662 680294
rect 202746 680058 202982 680294
rect 203826 708442 204062 708678
rect 204146 708442 204382 708678
rect 203826 708122 204062 708358
rect 204146 708122 204382 708358
rect 203826 694658 204062 694894
rect 204146 694658 204382 694894
rect 203826 694338 204062 694574
rect 204146 694338 204382 694574
rect 203826 658658 204062 658894
rect 204146 658658 204382 658894
rect 203826 658338 204062 658574
rect 204146 658338 204382 658574
rect 205226 707482 205462 707718
rect 205546 707482 205782 707718
rect 205226 707162 205462 707398
rect 205546 707162 205782 707398
rect 205226 672938 205462 673174
rect 205546 672938 205782 673174
rect 205226 672618 205462 672854
rect 205546 672618 205782 672854
rect 206626 704602 206862 704838
rect 206946 704602 207182 704838
rect 206626 704282 206862 704518
rect 206946 704282 207182 704518
rect 206626 687218 206862 687454
rect 206946 687218 207182 687454
rect 206626 686898 206862 687134
rect 206946 686898 207182 687134
rect 212666 711322 212902 711558
rect 212986 711322 213222 711558
rect 212666 711002 212902 711238
rect 212986 711002 213222 711238
rect 207546 698378 207782 698614
rect 207866 698378 208102 698614
rect 207546 698058 207782 698294
rect 207866 698058 208102 698294
rect 207546 662378 207782 662614
rect 207866 662378 208102 662614
rect 207546 662058 207782 662294
rect 207866 662058 208102 662294
rect 208946 709402 209182 709638
rect 209266 709402 209502 709638
rect 208946 709082 209182 709318
rect 209266 709082 209502 709318
rect 208946 676658 209182 676894
rect 209266 676658 209502 676894
rect 208946 676338 209182 676574
rect 209266 676338 209502 676574
rect 210346 706522 210582 706758
rect 210666 706522 210902 706758
rect 210346 706202 210582 706438
rect 210666 706202 210902 706438
rect 210346 690938 210582 691174
rect 210666 690938 210902 691174
rect 210346 690618 210582 690854
rect 210666 690618 210902 690854
rect 211746 705562 211982 705798
rect 212066 705562 212302 705798
rect 211746 705242 211982 705478
rect 212066 705242 212302 705478
rect 211746 669218 211982 669454
rect 212066 669218 212302 669454
rect 211746 668898 211982 669134
rect 212066 668898 212302 669134
rect 217786 710362 218022 710598
rect 218106 710362 218342 710598
rect 217786 710042 218022 710278
rect 218106 710042 218342 710278
rect 212666 680378 212902 680614
rect 212986 680378 213222 680614
rect 212666 680058 212902 680294
rect 212986 680058 213222 680294
rect 214066 708442 214302 708678
rect 214386 708442 214622 708678
rect 214066 708122 214302 708358
rect 214386 708122 214622 708358
rect 214066 694658 214302 694894
rect 214386 694658 214622 694894
rect 214066 694338 214302 694574
rect 214386 694338 214622 694574
rect 214066 658658 214302 658894
rect 214386 658658 214622 658894
rect 214066 658338 214302 658574
rect 214386 658338 214622 658574
rect 215466 707482 215702 707718
rect 215786 707482 216022 707718
rect 215466 707162 215702 707398
rect 215786 707162 216022 707398
rect 215466 672938 215702 673174
rect 215786 672938 216022 673174
rect 215466 672618 215702 672854
rect 215786 672618 216022 672854
rect 216866 704602 217102 704838
rect 217186 704602 217422 704838
rect 216866 704282 217102 704518
rect 217186 704282 217422 704518
rect 216866 687218 217102 687454
rect 217186 687218 217422 687454
rect 216866 686898 217102 687134
rect 217186 686898 217422 687134
rect 222906 711322 223142 711558
rect 223226 711322 223462 711558
rect 222906 711002 223142 711238
rect 223226 711002 223462 711238
rect 217786 698378 218022 698614
rect 218106 698378 218342 698614
rect 217786 698058 218022 698294
rect 218106 698058 218342 698294
rect 217786 662378 218022 662614
rect 218106 662378 218342 662614
rect 217786 662058 218022 662294
rect 218106 662058 218342 662294
rect 219186 709402 219422 709638
rect 219506 709402 219742 709638
rect 219186 709082 219422 709318
rect 219506 709082 219742 709318
rect 219186 676658 219422 676894
rect 219506 676658 219742 676894
rect 219186 676338 219422 676574
rect 219506 676338 219742 676574
rect 220586 706522 220822 706758
rect 220906 706522 221142 706758
rect 220586 706202 220822 706438
rect 220906 706202 221142 706438
rect 220586 690938 220822 691174
rect 220906 690938 221142 691174
rect 220586 690618 220822 690854
rect 220906 690618 221142 690854
rect 221986 705562 222222 705798
rect 222306 705562 222542 705798
rect 221986 705242 222222 705478
rect 222306 705242 222542 705478
rect 221986 669218 222222 669454
rect 222306 669218 222542 669454
rect 221986 668898 222222 669134
rect 222306 668898 222542 669134
rect 228026 710362 228262 710598
rect 228346 710362 228582 710598
rect 228026 710042 228262 710278
rect 228346 710042 228582 710278
rect 222906 680378 223142 680614
rect 223226 680378 223462 680614
rect 222906 680058 223142 680294
rect 223226 680058 223462 680294
rect 224306 708442 224542 708678
rect 224626 708442 224862 708678
rect 224306 708122 224542 708358
rect 224626 708122 224862 708358
rect 224306 694658 224542 694894
rect 224626 694658 224862 694894
rect 224306 694338 224542 694574
rect 224626 694338 224862 694574
rect 224306 658658 224542 658894
rect 224626 658658 224862 658894
rect 224306 658338 224542 658574
rect 224626 658338 224862 658574
rect 225706 707482 225942 707718
rect 226026 707482 226262 707718
rect 225706 707162 225942 707398
rect 226026 707162 226262 707398
rect 225706 672938 225942 673174
rect 226026 672938 226262 673174
rect 225706 672618 225942 672854
rect 226026 672618 226262 672854
rect 227106 704602 227342 704838
rect 227426 704602 227662 704838
rect 227106 704282 227342 704518
rect 227426 704282 227662 704518
rect 227106 687218 227342 687454
rect 227426 687218 227662 687454
rect 227106 686898 227342 687134
rect 227426 686898 227662 687134
rect 233146 711322 233382 711558
rect 233466 711322 233702 711558
rect 233146 711002 233382 711238
rect 233466 711002 233702 711238
rect 228026 698378 228262 698614
rect 228346 698378 228582 698614
rect 228026 698058 228262 698294
rect 228346 698058 228582 698294
rect 228026 662378 228262 662614
rect 228346 662378 228582 662614
rect 228026 662058 228262 662294
rect 228346 662058 228582 662294
rect 229426 709402 229662 709638
rect 229746 709402 229982 709638
rect 229426 709082 229662 709318
rect 229746 709082 229982 709318
rect 229426 676658 229662 676894
rect 229746 676658 229982 676894
rect 229426 676338 229662 676574
rect 229746 676338 229982 676574
rect 230826 706522 231062 706758
rect 231146 706522 231382 706758
rect 230826 706202 231062 706438
rect 231146 706202 231382 706438
rect 230826 690938 231062 691174
rect 231146 690938 231382 691174
rect 230826 690618 231062 690854
rect 231146 690618 231382 690854
rect 232226 705562 232462 705798
rect 232546 705562 232782 705798
rect 232226 705242 232462 705478
rect 232546 705242 232782 705478
rect 232226 669218 232462 669454
rect 232546 669218 232782 669454
rect 232226 668898 232462 669134
rect 232546 668898 232782 669134
rect 238266 710362 238502 710598
rect 238586 710362 238822 710598
rect 238266 710042 238502 710278
rect 238586 710042 238822 710278
rect 233146 680378 233382 680614
rect 233466 680378 233702 680614
rect 233146 680058 233382 680294
rect 233466 680058 233702 680294
rect 234546 708442 234782 708678
rect 234866 708442 235102 708678
rect 234546 708122 234782 708358
rect 234866 708122 235102 708358
rect 234546 694658 234782 694894
rect 234866 694658 235102 694894
rect 234546 694338 234782 694574
rect 234866 694338 235102 694574
rect 234546 658658 234782 658894
rect 234866 658658 235102 658894
rect 234546 658338 234782 658574
rect 234866 658338 235102 658574
rect 235946 707482 236182 707718
rect 236266 707482 236502 707718
rect 235946 707162 236182 707398
rect 236266 707162 236502 707398
rect 235946 672938 236182 673174
rect 236266 672938 236502 673174
rect 235946 672618 236182 672854
rect 236266 672618 236502 672854
rect 237346 704602 237582 704838
rect 237666 704602 237902 704838
rect 237346 704282 237582 704518
rect 237666 704282 237902 704518
rect 237346 687218 237582 687454
rect 237666 687218 237902 687454
rect 237346 686898 237582 687134
rect 237666 686898 237902 687134
rect 243386 711322 243622 711558
rect 243706 711322 243942 711558
rect 243386 711002 243622 711238
rect 243706 711002 243942 711238
rect 238266 698378 238502 698614
rect 238586 698378 238822 698614
rect 238266 698058 238502 698294
rect 238586 698058 238822 698294
rect 238266 662378 238502 662614
rect 238586 662378 238822 662614
rect 238266 662058 238502 662294
rect 238586 662058 238822 662294
rect 239666 709402 239902 709638
rect 239986 709402 240222 709638
rect 239666 709082 239902 709318
rect 239986 709082 240222 709318
rect 239666 676658 239902 676894
rect 239986 676658 240222 676894
rect 239666 676338 239902 676574
rect 239986 676338 240222 676574
rect 241066 706522 241302 706758
rect 241386 706522 241622 706758
rect 241066 706202 241302 706438
rect 241386 706202 241622 706438
rect 241066 690938 241302 691174
rect 241386 690938 241622 691174
rect 241066 690618 241302 690854
rect 241386 690618 241622 690854
rect 242466 705562 242702 705798
rect 242786 705562 243022 705798
rect 242466 705242 242702 705478
rect 242786 705242 243022 705478
rect 242466 669218 242702 669454
rect 242786 669218 243022 669454
rect 242466 668898 242702 669134
rect 242786 668898 243022 669134
rect 248506 710362 248742 710598
rect 248826 710362 249062 710598
rect 248506 710042 248742 710278
rect 248826 710042 249062 710278
rect 243386 680378 243622 680614
rect 243706 680378 243942 680614
rect 243386 680058 243622 680294
rect 243706 680058 243942 680294
rect 244786 708442 245022 708678
rect 245106 708442 245342 708678
rect 244786 708122 245022 708358
rect 245106 708122 245342 708358
rect 244786 694658 245022 694894
rect 245106 694658 245342 694894
rect 244786 694338 245022 694574
rect 245106 694338 245342 694574
rect 244786 658658 245022 658894
rect 245106 658658 245342 658894
rect 244786 658338 245022 658574
rect 245106 658338 245342 658574
rect 246186 707482 246422 707718
rect 246506 707482 246742 707718
rect 246186 707162 246422 707398
rect 246506 707162 246742 707398
rect 246186 672938 246422 673174
rect 246506 672938 246742 673174
rect 246186 672618 246422 672854
rect 246506 672618 246742 672854
rect 247586 704602 247822 704838
rect 247906 704602 248142 704838
rect 247586 704282 247822 704518
rect 247906 704282 248142 704518
rect 247586 687218 247822 687454
rect 247906 687218 248142 687454
rect 247586 686898 247822 687134
rect 247906 686898 248142 687134
rect 253626 711322 253862 711558
rect 253946 711322 254182 711558
rect 253626 711002 253862 711238
rect 253946 711002 254182 711238
rect 248506 698378 248742 698614
rect 248826 698378 249062 698614
rect 248506 698058 248742 698294
rect 248826 698058 249062 698294
rect 248506 662378 248742 662614
rect 248826 662378 249062 662614
rect 248506 662058 248742 662294
rect 248826 662058 249062 662294
rect 249906 709402 250142 709638
rect 250226 709402 250462 709638
rect 249906 709082 250142 709318
rect 250226 709082 250462 709318
rect 249906 676658 250142 676894
rect 250226 676658 250462 676894
rect 249906 676338 250142 676574
rect 250226 676338 250462 676574
rect 251306 706522 251542 706758
rect 251626 706522 251862 706758
rect 251306 706202 251542 706438
rect 251626 706202 251862 706438
rect 251306 690938 251542 691174
rect 251626 690938 251862 691174
rect 251306 690618 251542 690854
rect 251626 690618 251862 690854
rect 252706 705562 252942 705798
rect 253026 705562 253262 705798
rect 252706 705242 252942 705478
rect 253026 705242 253262 705478
rect 252706 669218 252942 669454
rect 253026 669218 253262 669454
rect 252706 668898 252942 669134
rect 253026 668898 253262 669134
rect 258746 710362 258982 710598
rect 259066 710362 259302 710598
rect 258746 710042 258982 710278
rect 259066 710042 259302 710278
rect 253626 680378 253862 680614
rect 253946 680378 254182 680614
rect 253626 680058 253862 680294
rect 253946 680058 254182 680294
rect 255026 708442 255262 708678
rect 255346 708442 255582 708678
rect 255026 708122 255262 708358
rect 255346 708122 255582 708358
rect 255026 694658 255262 694894
rect 255346 694658 255582 694894
rect 255026 694338 255262 694574
rect 255346 694338 255582 694574
rect 255026 658658 255262 658894
rect 255346 658658 255582 658894
rect 255026 658338 255262 658574
rect 255346 658338 255582 658574
rect 256426 707482 256662 707718
rect 256746 707482 256982 707718
rect 256426 707162 256662 707398
rect 256746 707162 256982 707398
rect 256426 672938 256662 673174
rect 256746 672938 256982 673174
rect 256426 672618 256662 672854
rect 256746 672618 256982 672854
rect 257826 704602 258062 704838
rect 258146 704602 258382 704838
rect 257826 704282 258062 704518
rect 258146 704282 258382 704518
rect 257826 687218 258062 687454
rect 258146 687218 258382 687454
rect 257826 686898 258062 687134
rect 258146 686898 258382 687134
rect 263866 711322 264102 711558
rect 264186 711322 264422 711558
rect 263866 711002 264102 711238
rect 264186 711002 264422 711238
rect 258746 698378 258982 698614
rect 259066 698378 259302 698614
rect 258746 698058 258982 698294
rect 259066 698058 259302 698294
rect 258746 662378 258982 662614
rect 259066 662378 259302 662614
rect 258746 662058 258982 662294
rect 259066 662058 259302 662294
rect 260146 709402 260382 709638
rect 260466 709402 260702 709638
rect 260146 709082 260382 709318
rect 260466 709082 260702 709318
rect 260146 676658 260382 676894
rect 260466 676658 260702 676894
rect 260146 676338 260382 676574
rect 260466 676338 260702 676574
rect 261546 706522 261782 706758
rect 261866 706522 262102 706758
rect 261546 706202 261782 706438
rect 261866 706202 262102 706438
rect 261546 690938 261782 691174
rect 261866 690938 262102 691174
rect 261546 690618 261782 690854
rect 261866 690618 262102 690854
rect 262946 705562 263182 705798
rect 263266 705562 263502 705798
rect 262946 705242 263182 705478
rect 263266 705242 263502 705478
rect 262946 669218 263182 669454
rect 263266 669218 263502 669454
rect 262946 668898 263182 669134
rect 263266 668898 263502 669134
rect 268986 710362 269222 710598
rect 269306 710362 269542 710598
rect 268986 710042 269222 710278
rect 269306 710042 269542 710278
rect 263866 680378 264102 680614
rect 264186 680378 264422 680614
rect 263866 680058 264102 680294
rect 264186 680058 264422 680294
rect 265266 708442 265502 708678
rect 265586 708442 265822 708678
rect 265266 708122 265502 708358
rect 265586 708122 265822 708358
rect 265266 694658 265502 694894
rect 265586 694658 265822 694894
rect 265266 694338 265502 694574
rect 265586 694338 265822 694574
rect 265266 658658 265502 658894
rect 265586 658658 265822 658894
rect 265266 658338 265502 658574
rect 265586 658338 265822 658574
rect 266666 707482 266902 707718
rect 266986 707482 267222 707718
rect 266666 707162 266902 707398
rect 266986 707162 267222 707398
rect 266666 672938 266902 673174
rect 266986 672938 267222 673174
rect 266666 672618 266902 672854
rect 266986 672618 267222 672854
rect 268066 704602 268302 704838
rect 268386 704602 268622 704838
rect 268066 704282 268302 704518
rect 268386 704282 268622 704518
rect 268066 687218 268302 687454
rect 268386 687218 268622 687454
rect 268066 686898 268302 687134
rect 268386 686898 268622 687134
rect 274106 711322 274342 711558
rect 274426 711322 274662 711558
rect 274106 711002 274342 711238
rect 274426 711002 274662 711238
rect 268986 698378 269222 698614
rect 269306 698378 269542 698614
rect 268986 698058 269222 698294
rect 269306 698058 269542 698294
rect 268986 662378 269222 662614
rect 269306 662378 269542 662614
rect 268986 662058 269222 662294
rect 269306 662058 269542 662294
rect 270386 709402 270622 709638
rect 270706 709402 270942 709638
rect 270386 709082 270622 709318
rect 270706 709082 270942 709318
rect 270386 676658 270622 676894
rect 270706 676658 270942 676894
rect 270386 676338 270622 676574
rect 270706 676338 270942 676574
rect 271786 706522 272022 706758
rect 272106 706522 272342 706758
rect 271786 706202 272022 706438
rect 272106 706202 272342 706438
rect 271786 690938 272022 691174
rect 272106 690938 272342 691174
rect 271786 690618 272022 690854
rect 272106 690618 272342 690854
rect 273186 705562 273422 705798
rect 273506 705562 273742 705798
rect 273186 705242 273422 705478
rect 273506 705242 273742 705478
rect 273186 669218 273422 669454
rect 273506 669218 273742 669454
rect 273186 668898 273422 669134
rect 273506 668898 273742 669134
rect 279226 710362 279462 710598
rect 279546 710362 279782 710598
rect 279226 710042 279462 710278
rect 279546 710042 279782 710278
rect 274106 680378 274342 680614
rect 274426 680378 274662 680614
rect 274106 680058 274342 680294
rect 274426 680058 274662 680294
rect 275506 708442 275742 708678
rect 275826 708442 276062 708678
rect 275506 708122 275742 708358
rect 275826 708122 276062 708358
rect 275506 694658 275742 694894
rect 275826 694658 276062 694894
rect 275506 694338 275742 694574
rect 275826 694338 276062 694574
rect 275506 658658 275742 658894
rect 275826 658658 276062 658894
rect 275506 658338 275742 658574
rect 275826 658338 276062 658574
rect 276906 707482 277142 707718
rect 277226 707482 277462 707718
rect 276906 707162 277142 707398
rect 277226 707162 277462 707398
rect 276906 672938 277142 673174
rect 277226 672938 277462 673174
rect 276906 672618 277142 672854
rect 277226 672618 277462 672854
rect 278306 704602 278542 704838
rect 278626 704602 278862 704838
rect 278306 704282 278542 704518
rect 278626 704282 278862 704518
rect 278306 687218 278542 687454
rect 278626 687218 278862 687454
rect 278306 686898 278542 687134
rect 278626 686898 278862 687134
rect 284346 711322 284582 711558
rect 284666 711322 284902 711558
rect 284346 711002 284582 711238
rect 284666 711002 284902 711238
rect 279226 698378 279462 698614
rect 279546 698378 279782 698614
rect 279226 698058 279462 698294
rect 279546 698058 279782 698294
rect 279226 662378 279462 662614
rect 279546 662378 279782 662614
rect 279226 662058 279462 662294
rect 279546 662058 279782 662294
rect 280626 709402 280862 709638
rect 280946 709402 281182 709638
rect 280626 709082 280862 709318
rect 280946 709082 281182 709318
rect 280626 676658 280862 676894
rect 280946 676658 281182 676894
rect 280626 676338 280862 676574
rect 280946 676338 281182 676574
rect 282026 706522 282262 706758
rect 282346 706522 282582 706758
rect 282026 706202 282262 706438
rect 282346 706202 282582 706438
rect 282026 690938 282262 691174
rect 282346 690938 282582 691174
rect 282026 690618 282262 690854
rect 282346 690618 282582 690854
rect 283426 705562 283662 705798
rect 283746 705562 283982 705798
rect 283426 705242 283662 705478
rect 283746 705242 283982 705478
rect 283426 669218 283662 669454
rect 283746 669218 283982 669454
rect 283426 668898 283662 669134
rect 283746 668898 283982 669134
rect 289466 710362 289702 710598
rect 289786 710362 290022 710598
rect 289466 710042 289702 710278
rect 289786 710042 290022 710278
rect 284346 680378 284582 680614
rect 284666 680378 284902 680614
rect 284346 680058 284582 680294
rect 284666 680058 284902 680294
rect 285746 708442 285982 708678
rect 286066 708442 286302 708678
rect 285746 708122 285982 708358
rect 286066 708122 286302 708358
rect 285746 694658 285982 694894
rect 286066 694658 286302 694894
rect 285746 694338 285982 694574
rect 286066 694338 286302 694574
rect 285746 658658 285982 658894
rect 286066 658658 286302 658894
rect 285746 658338 285982 658574
rect 286066 658338 286302 658574
rect 287146 707482 287382 707718
rect 287466 707482 287702 707718
rect 287146 707162 287382 707398
rect 287466 707162 287702 707398
rect 287146 672938 287382 673174
rect 287466 672938 287702 673174
rect 287146 672618 287382 672854
rect 287466 672618 287702 672854
rect 288546 704602 288782 704838
rect 288866 704602 289102 704838
rect 288546 704282 288782 704518
rect 288866 704282 289102 704518
rect 288546 687218 288782 687454
rect 288866 687218 289102 687454
rect 288546 686898 288782 687134
rect 288866 686898 289102 687134
rect 294586 711322 294822 711558
rect 294906 711322 295142 711558
rect 294586 711002 294822 711238
rect 294906 711002 295142 711238
rect 289466 698378 289702 698614
rect 289786 698378 290022 698614
rect 289466 698058 289702 698294
rect 289786 698058 290022 698294
rect 289466 662378 289702 662614
rect 289786 662378 290022 662614
rect 289466 662058 289702 662294
rect 289786 662058 290022 662294
rect 290866 709402 291102 709638
rect 291186 709402 291422 709638
rect 290866 709082 291102 709318
rect 291186 709082 291422 709318
rect 290866 676658 291102 676894
rect 291186 676658 291422 676894
rect 290866 676338 291102 676574
rect 291186 676338 291422 676574
rect 292266 706522 292502 706758
rect 292586 706522 292822 706758
rect 292266 706202 292502 706438
rect 292586 706202 292822 706438
rect 292266 690938 292502 691174
rect 292586 690938 292822 691174
rect 292266 690618 292502 690854
rect 292586 690618 292822 690854
rect 293666 705562 293902 705798
rect 293986 705562 294222 705798
rect 293666 705242 293902 705478
rect 293986 705242 294222 705478
rect 293666 669218 293902 669454
rect 293986 669218 294222 669454
rect 293666 668898 293902 669134
rect 293986 668898 294222 669134
rect 299706 710362 299942 710598
rect 300026 710362 300262 710598
rect 299706 710042 299942 710278
rect 300026 710042 300262 710278
rect 294586 680378 294822 680614
rect 294906 680378 295142 680614
rect 294586 680058 294822 680294
rect 294906 680058 295142 680294
rect 295986 708442 296222 708678
rect 296306 708442 296542 708678
rect 295986 708122 296222 708358
rect 296306 708122 296542 708358
rect 295986 694658 296222 694894
rect 296306 694658 296542 694894
rect 295986 694338 296222 694574
rect 296306 694338 296542 694574
rect 295986 658658 296222 658894
rect 296306 658658 296542 658894
rect 295986 658338 296222 658574
rect 296306 658338 296542 658574
rect 297386 707482 297622 707718
rect 297706 707482 297942 707718
rect 297386 707162 297622 707398
rect 297706 707162 297942 707398
rect 297386 672938 297622 673174
rect 297706 672938 297942 673174
rect 297386 672618 297622 672854
rect 297706 672618 297942 672854
rect 298786 704602 299022 704838
rect 299106 704602 299342 704838
rect 298786 704282 299022 704518
rect 299106 704282 299342 704518
rect 298786 687218 299022 687454
rect 299106 687218 299342 687454
rect 298786 686898 299022 687134
rect 299106 686898 299342 687134
rect 304826 711322 305062 711558
rect 305146 711322 305382 711558
rect 304826 711002 305062 711238
rect 305146 711002 305382 711238
rect 299706 698378 299942 698614
rect 300026 698378 300262 698614
rect 299706 698058 299942 698294
rect 300026 698058 300262 698294
rect 299706 662378 299942 662614
rect 300026 662378 300262 662614
rect 299706 662058 299942 662294
rect 300026 662058 300262 662294
rect 301106 709402 301342 709638
rect 301426 709402 301662 709638
rect 301106 709082 301342 709318
rect 301426 709082 301662 709318
rect 301106 676658 301342 676894
rect 301426 676658 301662 676894
rect 301106 676338 301342 676574
rect 301426 676338 301662 676574
rect 302506 706522 302742 706758
rect 302826 706522 303062 706758
rect 302506 706202 302742 706438
rect 302826 706202 303062 706438
rect 302506 690938 302742 691174
rect 302826 690938 303062 691174
rect 302506 690618 302742 690854
rect 302826 690618 303062 690854
rect 303906 705562 304142 705798
rect 304226 705562 304462 705798
rect 303906 705242 304142 705478
rect 304226 705242 304462 705478
rect 303906 669218 304142 669454
rect 304226 669218 304462 669454
rect 303906 668898 304142 669134
rect 304226 668898 304462 669134
rect 309946 710362 310182 710598
rect 310266 710362 310502 710598
rect 309946 710042 310182 710278
rect 310266 710042 310502 710278
rect 304826 680378 305062 680614
rect 305146 680378 305382 680614
rect 304826 680058 305062 680294
rect 305146 680058 305382 680294
rect 306226 708442 306462 708678
rect 306546 708442 306782 708678
rect 306226 708122 306462 708358
rect 306546 708122 306782 708358
rect 306226 694658 306462 694894
rect 306546 694658 306782 694894
rect 306226 694338 306462 694574
rect 306546 694338 306782 694574
rect 306226 658658 306462 658894
rect 306546 658658 306782 658894
rect 306226 658338 306462 658574
rect 306546 658338 306782 658574
rect 307626 707482 307862 707718
rect 307946 707482 308182 707718
rect 307626 707162 307862 707398
rect 307946 707162 308182 707398
rect 307626 672938 307862 673174
rect 307946 672938 308182 673174
rect 307626 672618 307862 672854
rect 307946 672618 308182 672854
rect 309026 704602 309262 704838
rect 309346 704602 309582 704838
rect 309026 704282 309262 704518
rect 309346 704282 309582 704518
rect 309026 687218 309262 687454
rect 309346 687218 309582 687454
rect 309026 686898 309262 687134
rect 309346 686898 309582 687134
rect 315066 711322 315302 711558
rect 315386 711322 315622 711558
rect 315066 711002 315302 711238
rect 315386 711002 315622 711238
rect 309946 698378 310182 698614
rect 310266 698378 310502 698614
rect 309946 698058 310182 698294
rect 310266 698058 310502 698294
rect 309946 662378 310182 662614
rect 310266 662378 310502 662614
rect 309946 662058 310182 662294
rect 310266 662058 310502 662294
rect 311346 709402 311582 709638
rect 311666 709402 311902 709638
rect 311346 709082 311582 709318
rect 311666 709082 311902 709318
rect 311346 676658 311582 676894
rect 311666 676658 311902 676894
rect 311346 676338 311582 676574
rect 311666 676338 311902 676574
rect 312746 706522 312982 706758
rect 313066 706522 313302 706758
rect 312746 706202 312982 706438
rect 313066 706202 313302 706438
rect 312746 690938 312982 691174
rect 313066 690938 313302 691174
rect 312746 690618 312982 690854
rect 313066 690618 313302 690854
rect 314146 705562 314382 705798
rect 314466 705562 314702 705798
rect 314146 705242 314382 705478
rect 314466 705242 314702 705478
rect 314146 669218 314382 669454
rect 314466 669218 314702 669454
rect 314146 668898 314382 669134
rect 314466 668898 314702 669134
rect 320186 710362 320422 710598
rect 320506 710362 320742 710598
rect 320186 710042 320422 710278
rect 320506 710042 320742 710278
rect 315066 680378 315302 680614
rect 315386 680378 315622 680614
rect 315066 680058 315302 680294
rect 315386 680058 315622 680294
rect 316466 708442 316702 708678
rect 316786 708442 317022 708678
rect 316466 708122 316702 708358
rect 316786 708122 317022 708358
rect 316466 694658 316702 694894
rect 316786 694658 317022 694894
rect 316466 694338 316702 694574
rect 316786 694338 317022 694574
rect 316466 658658 316702 658894
rect 316786 658658 317022 658894
rect 316466 658338 316702 658574
rect 316786 658338 317022 658574
rect 317866 707482 318102 707718
rect 318186 707482 318422 707718
rect 317866 707162 318102 707398
rect 318186 707162 318422 707398
rect 317866 672938 318102 673174
rect 318186 672938 318422 673174
rect 317866 672618 318102 672854
rect 318186 672618 318422 672854
rect 319266 704602 319502 704838
rect 319586 704602 319822 704838
rect 319266 704282 319502 704518
rect 319586 704282 319822 704518
rect 319266 687218 319502 687454
rect 319586 687218 319822 687454
rect 319266 686898 319502 687134
rect 319586 686898 319822 687134
rect 325306 711322 325542 711558
rect 325626 711322 325862 711558
rect 325306 711002 325542 711238
rect 325626 711002 325862 711238
rect 320186 698378 320422 698614
rect 320506 698378 320742 698614
rect 320186 698058 320422 698294
rect 320506 698058 320742 698294
rect 320186 662378 320422 662614
rect 320506 662378 320742 662614
rect 320186 662058 320422 662294
rect 320506 662058 320742 662294
rect 321586 709402 321822 709638
rect 321906 709402 322142 709638
rect 321586 709082 321822 709318
rect 321906 709082 322142 709318
rect 321586 676658 321822 676894
rect 321906 676658 322142 676894
rect 321586 676338 321822 676574
rect 321906 676338 322142 676574
rect 322986 706522 323222 706758
rect 323306 706522 323542 706758
rect 322986 706202 323222 706438
rect 323306 706202 323542 706438
rect 322986 690938 323222 691174
rect 323306 690938 323542 691174
rect 322986 690618 323222 690854
rect 323306 690618 323542 690854
rect 324386 705562 324622 705798
rect 324706 705562 324942 705798
rect 324386 705242 324622 705478
rect 324706 705242 324942 705478
rect 324386 669218 324622 669454
rect 324706 669218 324942 669454
rect 324386 668898 324622 669134
rect 324706 668898 324942 669134
rect 330426 710362 330662 710598
rect 330746 710362 330982 710598
rect 330426 710042 330662 710278
rect 330746 710042 330982 710278
rect 325306 680378 325542 680614
rect 325626 680378 325862 680614
rect 325306 680058 325542 680294
rect 325626 680058 325862 680294
rect 326706 708442 326942 708678
rect 327026 708442 327262 708678
rect 326706 708122 326942 708358
rect 327026 708122 327262 708358
rect 326706 694658 326942 694894
rect 327026 694658 327262 694894
rect 326706 694338 326942 694574
rect 327026 694338 327262 694574
rect 326706 658658 326942 658894
rect 327026 658658 327262 658894
rect 326706 658338 326942 658574
rect 327026 658338 327262 658574
rect 328106 707482 328342 707718
rect 328426 707482 328662 707718
rect 328106 707162 328342 707398
rect 328426 707162 328662 707398
rect 328106 672938 328342 673174
rect 328426 672938 328662 673174
rect 328106 672618 328342 672854
rect 328426 672618 328662 672854
rect 329506 704602 329742 704838
rect 329826 704602 330062 704838
rect 329506 704282 329742 704518
rect 329826 704282 330062 704518
rect 329506 687218 329742 687454
rect 329826 687218 330062 687454
rect 329506 686898 329742 687134
rect 329826 686898 330062 687134
rect 335546 711322 335782 711558
rect 335866 711322 336102 711558
rect 335546 711002 335782 711238
rect 335866 711002 336102 711238
rect 330426 698378 330662 698614
rect 330746 698378 330982 698614
rect 330426 698058 330662 698294
rect 330746 698058 330982 698294
rect 330426 662378 330662 662614
rect 330746 662378 330982 662614
rect 330426 662058 330662 662294
rect 330746 662058 330982 662294
rect 331826 709402 332062 709638
rect 332146 709402 332382 709638
rect 331826 709082 332062 709318
rect 332146 709082 332382 709318
rect 331826 676658 332062 676894
rect 332146 676658 332382 676894
rect 331826 676338 332062 676574
rect 332146 676338 332382 676574
rect 333226 706522 333462 706758
rect 333546 706522 333782 706758
rect 333226 706202 333462 706438
rect 333546 706202 333782 706438
rect 333226 690938 333462 691174
rect 333546 690938 333782 691174
rect 333226 690618 333462 690854
rect 333546 690618 333782 690854
rect 334626 705562 334862 705798
rect 334946 705562 335182 705798
rect 334626 705242 334862 705478
rect 334946 705242 335182 705478
rect 334626 669218 334862 669454
rect 334946 669218 335182 669454
rect 334626 668898 334862 669134
rect 334946 668898 335182 669134
rect 340666 710362 340902 710598
rect 340986 710362 341222 710598
rect 340666 710042 340902 710278
rect 340986 710042 341222 710278
rect 335546 680378 335782 680614
rect 335866 680378 336102 680614
rect 335546 680058 335782 680294
rect 335866 680058 336102 680294
rect 336946 708442 337182 708678
rect 337266 708442 337502 708678
rect 336946 708122 337182 708358
rect 337266 708122 337502 708358
rect 336946 694658 337182 694894
rect 337266 694658 337502 694894
rect 336946 694338 337182 694574
rect 337266 694338 337502 694574
rect 336946 658658 337182 658894
rect 337266 658658 337502 658894
rect 336946 658338 337182 658574
rect 337266 658338 337502 658574
rect 338346 707482 338582 707718
rect 338666 707482 338902 707718
rect 338346 707162 338582 707398
rect 338666 707162 338902 707398
rect 338346 672938 338582 673174
rect 338666 672938 338902 673174
rect 338346 672618 338582 672854
rect 338666 672618 338902 672854
rect 339746 704602 339982 704838
rect 340066 704602 340302 704838
rect 339746 704282 339982 704518
rect 340066 704282 340302 704518
rect 339746 687218 339982 687454
rect 340066 687218 340302 687454
rect 339746 686898 339982 687134
rect 340066 686898 340302 687134
rect 345786 711322 346022 711558
rect 346106 711322 346342 711558
rect 345786 711002 346022 711238
rect 346106 711002 346342 711238
rect 340666 698378 340902 698614
rect 340986 698378 341222 698614
rect 340666 698058 340902 698294
rect 340986 698058 341222 698294
rect 340666 662378 340902 662614
rect 340986 662378 341222 662614
rect 340666 662058 340902 662294
rect 340986 662058 341222 662294
rect 342066 709402 342302 709638
rect 342386 709402 342622 709638
rect 342066 709082 342302 709318
rect 342386 709082 342622 709318
rect 342066 676658 342302 676894
rect 342386 676658 342622 676894
rect 342066 676338 342302 676574
rect 342386 676338 342622 676574
rect 343466 706522 343702 706758
rect 343786 706522 344022 706758
rect 343466 706202 343702 706438
rect 343786 706202 344022 706438
rect 343466 690938 343702 691174
rect 343786 690938 344022 691174
rect 343466 690618 343702 690854
rect 343786 690618 344022 690854
rect 344866 705562 345102 705798
rect 345186 705562 345422 705798
rect 344866 705242 345102 705478
rect 345186 705242 345422 705478
rect 344866 669218 345102 669454
rect 345186 669218 345422 669454
rect 344866 668898 345102 669134
rect 345186 668898 345422 669134
rect 350906 710362 351142 710598
rect 351226 710362 351462 710598
rect 350906 710042 351142 710278
rect 351226 710042 351462 710278
rect 345786 680378 346022 680614
rect 346106 680378 346342 680614
rect 345786 680058 346022 680294
rect 346106 680058 346342 680294
rect 347186 708442 347422 708678
rect 347506 708442 347742 708678
rect 347186 708122 347422 708358
rect 347506 708122 347742 708358
rect 347186 694658 347422 694894
rect 347506 694658 347742 694894
rect 347186 694338 347422 694574
rect 347506 694338 347742 694574
rect 347186 658658 347422 658894
rect 347506 658658 347742 658894
rect 347186 658338 347422 658574
rect 347506 658338 347742 658574
rect 348586 707482 348822 707718
rect 348906 707482 349142 707718
rect 348586 707162 348822 707398
rect 348906 707162 349142 707398
rect 348586 672938 348822 673174
rect 348906 672938 349142 673174
rect 348586 672618 348822 672854
rect 348906 672618 349142 672854
rect 349986 704602 350222 704838
rect 350306 704602 350542 704838
rect 349986 704282 350222 704518
rect 350306 704282 350542 704518
rect 349986 687218 350222 687454
rect 350306 687218 350542 687454
rect 349986 686898 350222 687134
rect 350306 686898 350542 687134
rect 356026 711322 356262 711558
rect 356346 711322 356582 711558
rect 356026 711002 356262 711238
rect 356346 711002 356582 711238
rect 350906 698378 351142 698614
rect 351226 698378 351462 698614
rect 350906 698058 351142 698294
rect 351226 698058 351462 698294
rect 350906 662378 351142 662614
rect 351226 662378 351462 662614
rect 350906 662058 351142 662294
rect 351226 662058 351462 662294
rect 352306 709402 352542 709638
rect 352626 709402 352862 709638
rect 352306 709082 352542 709318
rect 352626 709082 352862 709318
rect 352306 676658 352542 676894
rect 352626 676658 352862 676894
rect 352306 676338 352542 676574
rect 352626 676338 352862 676574
rect 353706 706522 353942 706758
rect 354026 706522 354262 706758
rect 353706 706202 353942 706438
rect 354026 706202 354262 706438
rect 353706 690938 353942 691174
rect 354026 690938 354262 691174
rect 353706 690618 353942 690854
rect 354026 690618 354262 690854
rect 355106 705562 355342 705798
rect 355426 705562 355662 705798
rect 355106 705242 355342 705478
rect 355426 705242 355662 705478
rect 355106 669218 355342 669454
rect 355426 669218 355662 669454
rect 355106 668898 355342 669134
rect 355426 668898 355662 669134
rect 361146 710362 361382 710598
rect 361466 710362 361702 710598
rect 361146 710042 361382 710278
rect 361466 710042 361702 710278
rect 356026 680378 356262 680614
rect 356346 680378 356582 680614
rect 356026 680058 356262 680294
rect 356346 680058 356582 680294
rect 357426 708442 357662 708678
rect 357746 708442 357982 708678
rect 357426 708122 357662 708358
rect 357746 708122 357982 708358
rect 357426 694658 357662 694894
rect 357746 694658 357982 694894
rect 357426 694338 357662 694574
rect 357746 694338 357982 694574
rect 357426 658658 357662 658894
rect 357746 658658 357982 658894
rect 357426 658338 357662 658574
rect 357746 658338 357982 658574
rect 358826 707482 359062 707718
rect 359146 707482 359382 707718
rect 358826 707162 359062 707398
rect 359146 707162 359382 707398
rect 358826 672938 359062 673174
rect 359146 672938 359382 673174
rect 358826 672618 359062 672854
rect 359146 672618 359382 672854
rect 360226 704602 360462 704838
rect 360546 704602 360782 704838
rect 360226 704282 360462 704518
rect 360546 704282 360782 704518
rect 360226 687218 360462 687454
rect 360546 687218 360782 687454
rect 360226 686898 360462 687134
rect 360546 686898 360782 687134
rect 366266 711322 366502 711558
rect 366586 711322 366822 711558
rect 366266 711002 366502 711238
rect 366586 711002 366822 711238
rect 361146 698378 361382 698614
rect 361466 698378 361702 698614
rect 361146 698058 361382 698294
rect 361466 698058 361702 698294
rect 361146 662378 361382 662614
rect 361466 662378 361702 662614
rect 361146 662058 361382 662294
rect 361466 662058 361702 662294
rect 362546 709402 362782 709638
rect 362866 709402 363102 709638
rect 362546 709082 362782 709318
rect 362866 709082 363102 709318
rect 362546 676658 362782 676894
rect 362866 676658 363102 676894
rect 362546 676338 362782 676574
rect 362866 676338 363102 676574
rect 363946 706522 364182 706758
rect 364266 706522 364502 706758
rect 363946 706202 364182 706438
rect 364266 706202 364502 706438
rect 363946 690938 364182 691174
rect 364266 690938 364502 691174
rect 363946 690618 364182 690854
rect 364266 690618 364502 690854
rect 365346 705562 365582 705798
rect 365666 705562 365902 705798
rect 365346 705242 365582 705478
rect 365666 705242 365902 705478
rect 365346 669218 365582 669454
rect 365666 669218 365902 669454
rect 365346 668898 365582 669134
rect 365666 668898 365902 669134
rect 371386 710362 371622 710598
rect 371706 710362 371942 710598
rect 371386 710042 371622 710278
rect 371706 710042 371942 710278
rect 366266 680378 366502 680614
rect 366586 680378 366822 680614
rect 366266 680058 366502 680294
rect 366586 680058 366822 680294
rect 367666 708442 367902 708678
rect 367986 708442 368222 708678
rect 367666 708122 367902 708358
rect 367986 708122 368222 708358
rect 367666 694658 367902 694894
rect 367986 694658 368222 694894
rect 367666 694338 367902 694574
rect 367986 694338 368222 694574
rect 367666 658658 367902 658894
rect 367986 658658 368222 658894
rect 367666 658338 367902 658574
rect 367986 658338 368222 658574
rect 369066 707482 369302 707718
rect 369386 707482 369622 707718
rect 369066 707162 369302 707398
rect 369386 707162 369622 707398
rect 369066 672938 369302 673174
rect 369386 672938 369622 673174
rect 369066 672618 369302 672854
rect 369386 672618 369622 672854
rect 370466 704602 370702 704838
rect 370786 704602 371022 704838
rect 370466 704282 370702 704518
rect 370786 704282 371022 704518
rect 370466 687218 370702 687454
rect 370786 687218 371022 687454
rect 370466 686898 370702 687134
rect 370786 686898 371022 687134
rect 376506 711322 376742 711558
rect 376826 711322 377062 711558
rect 376506 711002 376742 711238
rect 376826 711002 377062 711238
rect 371386 698378 371622 698614
rect 371706 698378 371942 698614
rect 371386 698058 371622 698294
rect 371706 698058 371942 698294
rect 371386 662378 371622 662614
rect 371706 662378 371942 662614
rect 371386 662058 371622 662294
rect 371706 662058 371942 662294
rect 372786 709402 373022 709638
rect 373106 709402 373342 709638
rect 372786 709082 373022 709318
rect 373106 709082 373342 709318
rect 372786 676658 373022 676894
rect 373106 676658 373342 676894
rect 372786 676338 373022 676574
rect 373106 676338 373342 676574
rect 374186 706522 374422 706758
rect 374506 706522 374742 706758
rect 374186 706202 374422 706438
rect 374506 706202 374742 706438
rect 374186 690938 374422 691174
rect 374506 690938 374742 691174
rect 374186 690618 374422 690854
rect 374506 690618 374742 690854
rect 375586 705562 375822 705798
rect 375906 705562 376142 705798
rect 375586 705242 375822 705478
rect 375906 705242 376142 705478
rect 375586 669218 375822 669454
rect 375906 669218 376142 669454
rect 375586 668898 375822 669134
rect 375906 668898 376142 669134
rect 381626 710362 381862 710598
rect 381946 710362 382182 710598
rect 381626 710042 381862 710278
rect 381946 710042 382182 710278
rect 376506 680378 376742 680614
rect 376826 680378 377062 680614
rect 376506 680058 376742 680294
rect 376826 680058 377062 680294
rect 377906 708442 378142 708678
rect 378226 708442 378462 708678
rect 377906 708122 378142 708358
rect 378226 708122 378462 708358
rect 377906 694658 378142 694894
rect 378226 694658 378462 694894
rect 377906 694338 378142 694574
rect 378226 694338 378462 694574
rect 377906 658658 378142 658894
rect 378226 658658 378462 658894
rect 377906 658338 378142 658574
rect 378226 658338 378462 658574
rect 379306 707482 379542 707718
rect 379626 707482 379862 707718
rect 379306 707162 379542 707398
rect 379626 707162 379862 707398
rect 379306 672938 379542 673174
rect 379626 672938 379862 673174
rect 379306 672618 379542 672854
rect 379626 672618 379862 672854
rect 380706 704602 380942 704838
rect 381026 704602 381262 704838
rect 380706 704282 380942 704518
rect 381026 704282 381262 704518
rect 380706 687218 380942 687454
rect 381026 687218 381262 687454
rect 380706 686898 380942 687134
rect 381026 686898 381262 687134
rect 386746 711322 386982 711558
rect 387066 711322 387302 711558
rect 386746 711002 386982 711238
rect 387066 711002 387302 711238
rect 381626 698378 381862 698614
rect 381946 698378 382182 698614
rect 381626 698058 381862 698294
rect 381946 698058 382182 698294
rect 381626 662378 381862 662614
rect 381946 662378 382182 662614
rect 381626 662058 381862 662294
rect 381946 662058 382182 662294
rect 383026 709402 383262 709638
rect 383346 709402 383582 709638
rect 383026 709082 383262 709318
rect 383346 709082 383582 709318
rect 383026 676658 383262 676894
rect 383346 676658 383582 676894
rect 383026 676338 383262 676574
rect 383346 676338 383582 676574
rect 384426 706522 384662 706758
rect 384746 706522 384982 706758
rect 384426 706202 384662 706438
rect 384746 706202 384982 706438
rect 384426 690938 384662 691174
rect 384746 690938 384982 691174
rect 384426 690618 384662 690854
rect 384746 690618 384982 690854
rect 385826 705562 386062 705798
rect 386146 705562 386382 705798
rect 385826 705242 386062 705478
rect 386146 705242 386382 705478
rect 385826 669218 386062 669454
rect 386146 669218 386382 669454
rect 385826 668898 386062 669134
rect 386146 668898 386382 669134
rect 391866 710362 392102 710598
rect 392186 710362 392422 710598
rect 391866 710042 392102 710278
rect 392186 710042 392422 710278
rect 386746 680378 386982 680614
rect 387066 680378 387302 680614
rect 386746 680058 386982 680294
rect 387066 680058 387302 680294
rect 388146 708442 388382 708678
rect 388466 708442 388702 708678
rect 388146 708122 388382 708358
rect 388466 708122 388702 708358
rect 388146 694658 388382 694894
rect 388466 694658 388702 694894
rect 388146 694338 388382 694574
rect 388466 694338 388702 694574
rect 388146 658658 388382 658894
rect 388466 658658 388702 658894
rect 388146 658338 388382 658574
rect 388466 658338 388702 658574
rect 389546 707482 389782 707718
rect 389866 707482 390102 707718
rect 389546 707162 389782 707398
rect 389866 707162 390102 707398
rect 389546 672938 389782 673174
rect 389866 672938 390102 673174
rect 389546 672618 389782 672854
rect 389866 672618 390102 672854
rect 390946 704602 391182 704838
rect 391266 704602 391502 704838
rect 390946 704282 391182 704518
rect 391266 704282 391502 704518
rect 390946 687218 391182 687454
rect 391266 687218 391502 687454
rect 390946 686898 391182 687134
rect 391266 686898 391502 687134
rect 396986 711322 397222 711558
rect 397306 711322 397542 711558
rect 396986 711002 397222 711238
rect 397306 711002 397542 711238
rect 391866 698378 392102 698614
rect 392186 698378 392422 698614
rect 391866 698058 392102 698294
rect 392186 698058 392422 698294
rect 391866 662378 392102 662614
rect 392186 662378 392422 662614
rect 391866 662058 392102 662294
rect 392186 662058 392422 662294
rect 393266 709402 393502 709638
rect 393586 709402 393822 709638
rect 393266 709082 393502 709318
rect 393586 709082 393822 709318
rect 393266 676658 393502 676894
rect 393586 676658 393822 676894
rect 393266 676338 393502 676574
rect 393586 676338 393822 676574
rect 394666 706522 394902 706758
rect 394986 706522 395222 706758
rect 394666 706202 394902 706438
rect 394986 706202 395222 706438
rect 394666 690938 394902 691174
rect 394986 690938 395222 691174
rect 394666 690618 394902 690854
rect 394986 690618 395222 690854
rect 396066 705562 396302 705798
rect 396386 705562 396622 705798
rect 396066 705242 396302 705478
rect 396386 705242 396622 705478
rect 396066 669218 396302 669454
rect 396386 669218 396622 669454
rect 396066 668898 396302 669134
rect 396386 668898 396622 669134
rect 402106 710362 402342 710598
rect 402426 710362 402662 710598
rect 402106 710042 402342 710278
rect 402426 710042 402662 710278
rect 396986 680378 397222 680614
rect 397306 680378 397542 680614
rect 396986 680058 397222 680294
rect 397306 680058 397542 680294
rect 398386 708442 398622 708678
rect 398706 708442 398942 708678
rect 398386 708122 398622 708358
rect 398706 708122 398942 708358
rect 398386 694658 398622 694894
rect 398706 694658 398942 694894
rect 398386 694338 398622 694574
rect 398706 694338 398942 694574
rect 398386 658658 398622 658894
rect 398706 658658 398942 658894
rect 398386 658338 398622 658574
rect 398706 658338 398942 658574
rect 399786 707482 400022 707718
rect 400106 707482 400342 707718
rect 399786 707162 400022 707398
rect 400106 707162 400342 707398
rect 399786 672938 400022 673174
rect 400106 672938 400342 673174
rect 399786 672618 400022 672854
rect 400106 672618 400342 672854
rect 401186 704602 401422 704838
rect 401506 704602 401742 704838
rect 401186 704282 401422 704518
rect 401506 704282 401742 704518
rect 401186 687218 401422 687454
rect 401506 687218 401742 687454
rect 401186 686898 401422 687134
rect 401506 686898 401742 687134
rect 407226 711322 407462 711558
rect 407546 711322 407782 711558
rect 407226 711002 407462 711238
rect 407546 711002 407782 711238
rect 402106 698378 402342 698614
rect 402426 698378 402662 698614
rect 402106 698058 402342 698294
rect 402426 698058 402662 698294
rect 402106 662378 402342 662614
rect 402426 662378 402662 662614
rect 402106 662058 402342 662294
rect 402426 662058 402662 662294
rect 403506 709402 403742 709638
rect 403826 709402 404062 709638
rect 403506 709082 403742 709318
rect 403826 709082 404062 709318
rect 403506 676658 403742 676894
rect 403826 676658 404062 676894
rect 403506 676338 403742 676574
rect 403826 676338 404062 676574
rect 404906 706522 405142 706758
rect 405226 706522 405462 706758
rect 404906 706202 405142 706438
rect 405226 706202 405462 706438
rect 404906 690938 405142 691174
rect 405226 690938 405462 691174
rect 404906 690618 405142 690854
rect 405226 690618 405462 690854
rect 406306 705562 406542 705798
rect 406626 705562 406862 705798
rect 406306 705242 406542 705478
rect 406626 705242 406862 705478
rect 406306 669218 406542 669454
rect 406626 669218 406862 669454
rect 406306 668898 406542 669134
rect 406626 668898 406862 669134
rect 412346 710362 412582 710598
rect 412666 710362 412902 710598
rect 412346 710042 412582 710278
rect 412666 710042 412902 710278
rect 407226 680378 407462 680614
rect 407546 680378 407782 680614
rect 407226 680058 407462 680294
rect 407546 680058 407782 680294
rect 408626 708442 408862 708678
rect 408946 708442 409182 708678
rect 408626 708122 408862 708358
rect 408946 708122 409182 708358
rect 408626 694658 408862 694894
rect 408946 694658 409182 694894
rect 408626 694338 408862 694574
rect 408946 694338 409182 694574
rect 408626 658658 408862 658894
rect 408946 658658 409182 658894
rect 408626 658338 408862 658574
rect 408946 658338 409182 658574
rect 410026 707482 410262 707718
rect 410346 707482 410582 707718
rect 410026 707162 410262 707398
rect 410346 707162 410582 707398
rect 410026 672938 410262 673174
rect 410346 672938 410582 673174
rect 410026 672618 410262 672854
rect 410346 672618 410582 672854
rect 411426 704602 411662 704838
rect 411746 704602 411982 704838
rect 411426 704282 411662 704518
rect 411746 704282 411982 704518
rect 411426 687218 411662 687454
rect 411746 687218 411982 687454
rect 411426 686898 411662 687134
rect 411746 686898 411982 687134
rect 417466 711322 417702 711558
rect 417786 711322 418022 711558
rect 417466 711002 417702 711238
rect 417786 711002 418022 711238
rect 412346 698378 412582 698614
rect 412666 698378 412902 698614
rect 412346 698058 412582 698294
rect 412666 698058 412902 698294
rect 412346 662378 412582 662614
rect 412666 662378 412902 662614
rect 412346 662058 412582 662294
rect 412666 662058 412902 662294
rect 413746 709402 413982 709638
rect 414066 709402 414302 709638
rect 413746 709082 413982 709318
rect 414066 709082 414302 709318
rect 413746 676658 413982 676894
rect 414066 676658 414302 676894
rect 413746 676338 413982 676574
rect 414066 676338 414302 676574
rect 415146 706522 415382 706758
rect 415466 706522 415702 706758
rect 415146 706202 415382 706438
rect 415466 706202 415702 706438
rect 415146 690938 415382 691174
rect 415466 690938 415702 691174
rect 415146 690618 415382 690854
rect 415466 690618 415702 690854
rect 416546 705562 416782 705798
rect 416866 705562 417102 705798
rect 416546 705242 416782 705478
rect 416866 705242 417102 705478
rect 416546 669218 416782 669454
rect 416866 669218 417102 669454
rect 416546 668898 416782 669134
rect 416866 668898 417102 669134
rect 422586 710362 422822 710598
rect 422906 710362 423142 710598
rect 422586 710042 422822 710278
rect 422906 710042 423142 710278
rect 417466 680378 417702 680614
rect 417786 680378 418022 680614
rect 417466 680058 417702 680294
rect 417786 680058 418022 680294
rect 418866 708442 419102 708678
rect 419186 708442 419422 708678
rect 418866 708122 419102 708358
rect 419186 708122 419422 708358
rect 418866 694658 419102 694894
rect 419186 694658 419422 694894
rect 418866 694338 419102 694574
rect 419186 694338 419422 694574
rect 418866 658658 419102 658894
rect 419186 658658 419422 658894
rect 418866 658338 419102 658574
rect 419186 658338 419422 658574
rect 420266 707482 420502 707718
rect 420586 707482 420822 707718
rect 420266 707162 420502 707398
rect 420586 707162 420822 707398
rect 420266 672938 420502 673174
rect 420586 672938 420822 673174
rect 420266 672618 420502 672854
rect 420586 672618 420822 672854
rect 421666 704602 421902 704838
rect 421986 704602 422222 704838
rect 421666 704282 421902 704518
rect 421986 704282 422222 704518
rect 421666 687218 421902 687454
rect 421986 687218 422222 687454
rect 421666 686898 421902 687134
rect 421986 686898 422222 687134
rect 427706 711322 427942 711558
rect 428026 711322 428262 711558
rect 427706 711002 427942 711238
rect 428026 711002 428262 711238
rect 422586 698378 422822 698614
rect 422906 698378 423142 698614
rect 422586 698058 422822 698294
rect 422906 698058 423142 698294
rect 422586 662378 422822 662614
rect 422906 662378 423142 662614
rect 422586 662058 422822 662294
rect 422906 662058 423142 662294
rect 423986 709402 424222 709638
rect 424306 709402 424542 709638
rect 423986 709082 424222 709318
rect 424306 709082 424542 709318
rect 423986 676658 424222 676894
rect 424306 676658 424542 676894
rect 423986 676338 424222 676574
rect 424306 676338 424542 676574
rect 425386 706522 425622 706758
rect 425706 706522 425942 706758
rect 425386 706202 425622 706438
rect 425706 706202 425942 706438
rect 425386 690938 425622 691174
rect 425706 690938 425942 691174
rect 425386 690618 425622 690854
rect 425706 690618 425942 690854
rect 426786 705562 427022 705798
rect 427106 705562 427342 705798
rect 426786 705242 427022 705478
rect 427106 705242 427342 705478
rect 426786 669218 427022 669454
rect 427106 669218 427342 669454
rect 426786 668898 427022 669134
rect 427106 668898 427342 669134
rect 432826 710362 433062 710598
rect 433146 710362 433382 710598
rect 432826 710042 433062 710278
rect 433146 710042 433382 710278
rect 427706 680378 427942 680614
rect 428026 680378 428262 680614
rect 427706 680058 427942 680294
rect 428026 680058 428262 680294
rect 429106 708442 429342 708678
rect 429426 708442 429662 708678
rect 429106 708122 429342 708358
rect 429426 708122 429662 708358
rect 429106 694658 429342 694894
rect 429426 694658 429662 694894
rect 429106 694338 429342 694574
rect 429426 694338 429662 694574
rect 429106 658658 429342 658894
rect 429426 658658 429662 658894
rect 429106 658338 429342 658574
rect 429426 658338 429662 658574
rect 430506 707482 430742 707718
rect 430826 707482 431062 707718
rect 430506 707162 430742 707398
rect 430826 707162 431062 707398
rect 430506 672938 430742 673174
rect 430826 672938 431062 673174
rect 430506 672618 430742 672854
rect 430826 672618 431062 672854
rect 431906 704602 432142 704838
rect 432226 704602 432462 704838
rect 431906 704282 432142 704518
rect 432226 704282 432462 704518
rect 431906 687218 432142 687454
rect 432226 687218 432462 687454
rect 431906 686898 432142 687134
rect 432226 686898 432462 687134
rect 437946 711322 438182 711558
rect 438266 711322 438502 711558
rect 437946 711002 438182 711238
rect 438266 711002 438502 711238
rect 432826 698378 433062 698614
rect 433146 698378 433382 698614
rect 432826 698058 433062 698294
rect 433146 698058 433382 698294
rect 432826 662378 433062 662614
rect 433146 662378 433382 662614
rect 432826 662058 433062 662294
rect 433146 662058 433382 662294
rect 434226 709402 434462 709638
rect 434546 709402 434782 709638
rect 434226 709082 434462 709318
rect 434546 709082 434782 709318
rect 434226 676658 434462 676894
rect 434546 676658 434782 676894
rect 434226 676338 434462 676574
rect 434546 676338 434782 676574
rect 435626 706522 435862 706758
rect 435946 706522 436182 706758
rect 435626 706202 435862 706438
rect 435946 706202 436182 706438
rect 435626 690938 435862 691174
rect 435946 690938 436182 691174
rect 435626 690618 435862 690854
rect 435946 690618 436182 690854
rect 437026 705562 437262 705798
rect 437346 705562 437582 705798
rect 437026 705242 437262 705478
rect 437346 705242 437582 705478
rect 437026 669218 437262 669454
rect 437346 669218 437582 669454
rect 437026 668898 437262 669134
rect 437346 668898 437582 669134
rect 443066 710362 443302 710598
rect 443386 710362 443622 710598
rect 443066 710042 443302 710278
rect 443386 710042 443622 710278
rect 437946 680378 438182 680614
rect 438266 680378 438502 680614
rect 437946 680058 438182 680294
rect 438266 680058 438502 680294
rect 439346 708442 439582 708678
rect 439666 708442 439902 708678
rect 439346 708122 439582 708358
rect 439666 708122 439902 708358
rect 439346 694658 439582 694894
rect 439666 694658 439902 694894
rect 439346 694338 439582 694574
rect 439666 694338 439902 694574
rect 439346 658658 439582 658894
rect 439666 658658 439902 658894
rect 439346 658338 439582 658574
rect 439666 658338 439902 658574
rect 440746 707482 440982 707718
rect 441066 707482 441302 707718
rect 440746 707162 440982 707398
rect 441066 707162 441302 707398
rect 440746 672938 440982 673174
rect 441066 672938 441302 673174
rect 440746 672618 440982 672854
rect 441066 672618 441302 672854
rect 442146 704602 442382 704838
rect 442466 704602 442702 704838
rect 442146 704282 442382 704518
rect 442466 704282 442702 704518
rect 442146 687218 442382 687454
rect 442466 687218 442702 687454
rect 442146 686898 442382 687134
rect 442466 686898 442702 687134
rect 448186 711322 448422 711558
rect 448506 711322 448742 711558
rect 448186 711002 448422 711238
rect 448506 711002 448742 711238
rect 443066 698378 443302 698614
rect 443386 698378 443622 698614
rect 443066 698058 443302 698294
rect 443386 698058 443622 698294
rect 443066 662378 443302 662614
rect 443386 662378 443622 662614
rect 443066 662058 443302 662294
rect 443386 662058 443622 662294
rect 444466 709402 444702 709638
rect 444786 709402 445022 709638
rect 444466 709082 444702 709318
rect 444786 709082 445022 709318
rect 444466 676658 444702 676894
rect 444786 676658 445022 676894
rect 444466 676338 444702 676574
rect 444786 676338 445022 676574
rect 445866 706522 446102 706758
rect 446186 706522 446422 706758
rect 445866 706202 446102 706438
rect 446186 706202 446422 706438
rect 445866 690938 446102 691174
rect 446186 690938 446422 691174
rect 445866 690618 446102 690854
rect 446186 690618 446422 690854
rect 447266 705562 447502 705798
rect 447586 705562 447822 705798
rect 447266 705242 447502 705478
rect 447586 705242 447822 705478
rect 447266 669218 447502 669454
rect 447586 669218 447822 669454
rect 447266 668898 447502 669134
rect 447586 668898 447822 669134
rect 453306 710362 453542 710598
rect 453626 710362 453862 710598
rect 453306 710042 453542 710278
rect 453626 710042 453862 710278
rect 448186 680378 448422 680614
rect 448506 680378 448742 680614
rect 448186 680058 448422 680294
rect 448506 680058 448742 680294
rect 449586 708442 449822 708678
rect 449906 708442 450142 708678
rect 449586 708122 449822 708358
rect 449906 708122 450142 708358
rect 449586 694658 449822 694894
rect 449906 694658 450142 694894
rect 449586 694338 449822 694574
rect 449906 694338 450142 694574
rect 449586 658658 449822 658894
rect 449906 658658 450142 658894
rect 449586 658338 449822 658574
rect 449906 658338 450142 658574
rect 450986 707482 451222 707718
rect 451306 707482 451542 707718
rect 450986 707162 451222 707398
rect 451306 707162 451542 707398
rect 450986 672938 451222 673174
rect 451306 672938 451542 673174
rect 450986 672618 451222 672854
rect 451306 672618 451542 672854
rect 452386 704602 452622 704838
rect 452706 704602 452942 704838
rect 452386 704282 452622 704518
rect 452706 704282 452942 704518
rect 452386 687218 452622 687454
rect 452706 687218 452942 687454
rect 452386 686898 452622 687134
rect 452706 686898 452942 687134
rect 458426 711322 458662 711558
rect 458746 711322 458982 711558
rect 458426 711002 458662 711238
rect 458746 711002 458982 711238
rect 453306 698378 453542 698614
rect 453626 698378 453862 698614
rect 453306 698058 453542 698294
rect 453626 698058 453862 698294
rect 453306 662378 453542 662614
rect 453626 662378 453862 662614
rect 453306 662058 453542 662294
rect 453626 662058 453862 662294
rect 454706 709402 454942 709638
rect 455026 709402 455262 709638
rect 454706 709082 454942 709318
rect 455026 709082 455262 709318
rect 454706 676658 454942 676894
rect 455026 676658 455262 676894
rect 454706 676338 454942 676574
rect 455026 676338 455262 676574
rect 456106 706522 456342 706758
rect 456426 706522 456662 706758
rect 456106 706202 456342 706438
rect 456426 706202 456662 706438
rect 456106 690938 456342 691174
rect 456426 690938 456662 691174
rect 456106 690618 456342 690854
rect 456426 690618 456662 690854
rect 457506 705562 457742 705798
rect 457826 705562 458062 705798
rect 457506 705242 457742 705478
rect 457826 705242 458062 705478
rect 457506 669218 457742 669454
rect 457826 669218 458062 669454
rect 457506 668898 457742 669134
rect 457826 668898 458062 669134
rect 463546 710362 463782 710598
rect 463866 710362 464102 710598
rect 463546 710042 463782 710278
rect 463866 710042 464102 710278
rect 458426 680378 458662 680614
rect 458746 680378 458982 680614
rect 458426 680058 458662 680294
rect 458746 680058 458982 680294
rect 459826 708442 460062 708678
rect 460146 708442 460382 708678
rect 459826 708122 460062 708358
rect 460146 708122 460382 708358
rect 459826 694658 460062 694894
rect 460146 694658 460382 694894
rect 459826 694338 460062 694574
rect 460146 694338 460382 694574
rect 459826 658658 460062 658894
rect 460146 658658 460382 658894
rect 459826 658338 460062 658574
rect 460146 658338 460382 658574
rect 461226 707482 461462 707718
rect 461546 707482 461782 707718
rect 461226 707162 461462 707398
rect 461546 707162 461782 707398
rect 461226 672938 461462 673174
rect 461546 672938 461782 673174
rect 461226 672618 461462 672854
rect 461546 672618 461782 672854
rect 462626 704602 462862 704838
rect 462946 704602 463182 704838
rect 462626 704282 462862 704518
rect 462946 704282 463182 704518
rect 462626 687218 462862 687454
rect 462946 687218 463182 687454
rect 462626 686898 462862 687134
rect 462946 686898 463182 687134
rect 468666 711322 468902 711558
rect 468986 711322 469222 711558
rect 468666 711002 468902 711238
rect 468986 711002 469222 711238
rect 463546 698378 463782 698614
rect 463866 698378 464102 698614
rect 463546 698058 463782 698294
rect 463866 698058 464102 698294
rect 463546 662378 463782 662614
rect 463866 662378 464102 662614
rect 463546 662058 463782 662294
rect 463866 662058 464102 662294
rect 464946 709402 465182 709638
rect 465266 709402 465502 709638
rect 464946 709082 465182 709318
rect 465266 709082 465502 709318
rect 464946 676658 465182 676894
rect 465266 676658 465502 676894
rect 464946 676338 465182 676574
rect 465266 676338 465502 676574
rect 466346 706522 466582 706758
rect 466666 706522 466902 706758
rect 466346 706202 466582 706438
rect 466666 706202 466902 706438
rect 466346 690938 466582 691174
rect 466666 690938 466902 691174
rect 466346 690618 466582 690854
rect 466666 690618 466902 690854
rect 467746 705562 467982 705798
rect 468066 705562 468302 705798
rect 467746 705242 467982 705478
rect 468066 705242 468302 705478
rect 467746 669218 467982 669454
rect 468066 669218 468302 669454
rect 467746 668898 467982 669134
rect 468066 668898 468302 669134
rect 473786 710362 474022 710598
rect 474106 710362 474342 710598
rect 473786 710042 474022 710278
rect 474106 710042 474342 710278
rect 468666 680378 468902 680614
rect 468986 680378 469222 680614
rect 468666 680058 468902 680294
rect 468986 680058 469222 680294
rect 470066 708442 470302 708678
rect 470386 708442 470622 708678
rect 470066 708122 470302 708358
rect 470386 708122 470622 708358
rect 470066 694658 470302 694894
rect 470386 694658 470622 694894
rect 470066 694338 470302 694574
rect 470386 694338 470622 694574
rect 470066 658658 470302 658894
rect 470386 658658 470622 658894
rect 470066 658338 470302 658574
rect 470386 658338 470622 658574
rect 471466 707482 471702 707718
rect 471786 707482 472022 707718
rect 471466 707162 471702 707398
rect 471786 707162 472022 707398
rect 471466 672938 471702 673174
rect 471786 672938 472022 673174
rect 471466 672618 471702 672854
rect 471786 672618 472022 672854
rect 472866 704602 473102 704838
rect 473186 704602 473422 704838
rect 472866 704282 473102 704518
rect 473186 704282 473422 704518
rect 472866 687218 473102 687454
rect 473186 687218 473422 687454
rect 472866 686898 473102 687134
rect 473186 686898 473422 687134
rect 478906 711322 479142 711558
rect 479226 711322 479462 711558
rect 478906 711002 479142 711238
rect 479226 711002 479462 711238
rect 473786 698378 474022 698614
rect 474106 698378 474342 698614
rect 473786 698058 474022 698294
rect 474106 698058 474342 698294
rect 473786 662378 474022 662614
rect 474106 662378 474342 662614
rect 473786 662058 474022 662294
rect 474106 662058 474342 662294
rect 475186 709402 475422 709638
rect 475506 709402 475742 709638
rect 475186 709082 475422 709318
rect 475506 709082 475742 709318
rect 475186 676658 475422 676894
rect 475506 676658 475742 676894
rect 475186 676338 475422 676574
rect 475506 676338 475742 676574
rect 476586 706522 476822 706758
rect 476906 706522 477142 706758
rect 476586 706202 476822 706438
rect 476906 706202 477142 706438
rect 476586 690938 476822 691174
rect 476906 690938 477142 691174
rect 476586 690618 476822 690854
rect 476906 690618 477142 690854
rect 477986 705562 478222 705798
rect 478306 705562 478542 705798
rect 477986 705242 478222 705478
rect 478306 705242 478542 705478
rect 477986 669218 478222 669454
rect 478306 669218 478542 669454
rect 477986 668898 478222 669134
rect 478306 668898 478542 669134
rect 484026 710362 484262 710598
rect 484346 710362 484582 710598
rect 484026 710042 484262 710278
rect 484346 710042 484582 710278
rect 478906 680378 479142 680614
rect 479226 680378 479462 680614
rect 478906 680058 479142 680294
rect 479226 680058 479462 680294
rect 480306 708442 480542 708678
rect 480626 708442 480862 708678
rect 480306 708122 480542 708358
rect 480626 708122 480862 708358
rect 480306 694658 480542 694894
rect 480626 694658 480862 694894
rect 480306 694338 480542 694574
rect 480626 694338 480862 694574
rect 480306 658658 480542 658894
rect 480626 658658 480862 658894
rect 480306 658338 480542 658574
rect 480626 658338 480862 658574
rect 481706 707482 481942 707718
rect 482026 707482 482262 707718
rect 481706 707162 481942 707398
rect 482026 707162 482262 707398
rect 481706 672938 481942 673174
rect 482026 672938 482262 673174
rect 481706 672618 481942 672854
rect 482026 672618 482262 672854
rect 483106 704602 483342 704838
rect 483426 704602 483662 704838
rect 483106 704282 483342 704518
rect 483426 704282 483662 704518
rect 483106 687218 483342 687454
rect 483426 687218 483662 687454
rect 483106 686898 483342 687134
rect 483426 686898 483662 687134
rect 489146 711322 489382 711558
rect 489466 711322 489702 711558
rect 489146 711002 489382 711238
rect 489466 711002 489702 711238
rect 484026 698378 484262 698614
rect 484346 698378 484582 698614
rect 484026 698058 484262 698294
rect 484346 698058 484582 698294
rect 484026 662378 484262 662614
rect 484346 662378 484582 662614
rect 484026 662058 484262 662294
rect 484346 662058 484582 662294
rect 485426 709402 485662 709638
rect 485746 709402 485982 709638
rect 485426 709082 485662 709318
rect 485746 709082 485982 709318
rect 485426 676658 485662 676894
rect 485746 676658 485982 676894
rect 485426 676338 485662 676574
rect 485746 676338 485982 676574
rect 486826 706522 487062 706758
rect 487146 706522 487382 706758
rect 486826 706202 487062 706438
rect 487146 706202 487382 706438
rect 486826 690938 487062 691174
rect 487146 690938 487382 691174
rect 486826 690618 487062 690854
rect 487146 690618 487382 690854
rect 488226 705562 488462 705798
rect 488546 705562 488782 705798
rect 488226 705242 488462 705478
rect 488546 705242 488782 705478
rect 488226 669218 488462 669454
rect 488546 669218 488782 669454
rect 488226 668898 488462 669134
rect 488546 668898 488782 669134
rect 494266 710362 494502 710598
rect 494586 710362 494822 710598
rect 494266 710042 494502 710278
rect 494586 710042 494822 710278
rect 489146 680378 489382 680614
rect 489466 680378 489702 680614
rect 489146 680058 489382 680294
rect 489466 680058 489702 680294
rect 490546 708442 490782 708678
rect 490866 708442 491102 708678
rect 490546 708122 490782 708358
rect 490866 708122 491102 708358
rect 490546 694658 490782 694894
rect 490866 694658 491102 694894
rect 490546 694338 490782 694574
rect 490866 694338 491102 694574
rect 490546 658658 490782 658894
rect 490866 658658 491102 658894
rect 490546 658338 490782 658574
rect 490866 658338 491102 658574
rect 491946 707482 492182 707718
rect 492266 707482 492502 707718
rect 491946 707162 492182 707398
rect 492266 707162 492502 707398
rect 491946 672938 492182 673174
rect 492266 672938 492502 673174
rect 491946 672618 492182 672854
rect 492266 672618 492502 672854
rect 493346 704602 493582 704838
rect 493666 704602 493902 704838
rect 493346 704282 493582 704518
rect 493666 704282 493902 704518
rect 493346 687218 493582 687454
rect 493666 687218 493902 687454
rect 493346 686898 493582 687134
rect 493666 686898 493902 687134
rect 499386 711322 499622 711558
rect 499706 711322 499942 711558
rect 499386 711002 499622 711238
rect 499706 711002 499942 711238
rect 494266 698378 494502 698614
rect 494586 698378 494822 698614
rect 494266 698058 494502 698294
rect 494586 698058 494822 698294
rect 494266 662378 494502 662614
rect 494586 662378 494822 662614
rect 494266 662058 494502 662294
rect 494586 662058 494822 662294
rect 495666 709402 495902 709638
rect 495986 709402 496222 709638
rect 495666 709082 495902 709318
rect 495986 709082 496222 709318
rect 495666 676658 495902 676894
rect 495986 676658 496222 676894
rect 495666 676338 495902 676574
rect 495986 676338 496222 676574
rect 497066 706522 497302 706758
rect 497386 706522 497622 706758
rect 497066 706202 497302 706438
rect 497386 706202 497622 706438
rect 497066 690938 497302 691174
rect 497386 690938 497622 691174
rect 497066 690618 497302 690854
rect 497386 690618 497622 690854
rect 498466 705562 498702 705798
rect 498786 705562 499022 705798
rect 498466 705242 498702 705478
rect 498786 705242 499022 705478
rect 498466 669218 498702 669454
rect 498786 669218 499022 669454
rect 498466 668898 498702 669134
rect 498786 668898 499022 669134
rect 504506 710362 504742 710598
rect 504826 710362 505062 710598
rect 504506 710042 504742 710278
rect 504826 710042 505062 710278
rect 499386 680378 499622 680614
rect 499706 680378 499942 680614
rect 499386 680058 499622 680294
rect 499706 680058 499942 680294
rect 500786 708442 501022 708678
rect 501106 708442 501342 708678
rect 500786 708122 501022 708358
rect 501106 708122 501342 708358
rect 500786 694658 501022 694894
rect 501106 694658 501342 694894
rect 500786 694338 501022 694574
rect 501106 694338 501342 694574
rect 500786 658658 501022 658894
rect 501106 658658 501342 658894
rect 500786 658338 501022 658574
rect 501106 658338 501342 658574
rect 502186 707482 502422 707718
rect 502506 707482 502742 707718
rect 502186 707162 502422 707398
rect 502506 707162 502742 707398
rect 502186 672938 502422 673174
rect 502506 672938 502742 673174
rect 502186 672618 502422 672854
rect 502506 672618 502742 672854
rect 503586 704602 503822 704838
rect 503906 704602 504142 704838
rect 503586 704282 503822 704518
rect 503906 704282 504142 704518
rect 503586 687218 503822 687454
rect 503906 687218 504142 687454
rect 503586 686898 503822 687134
rect 503906 686898 504142 687134
rect 509626 711322 509862 711558
rect 509946 711322 510182 711558
rect 509626 711002 509862 711238
rect 509946 711002 510182 711238
rect 504506 698378 504742 698614
rect 504826 698378 505062 698614
rect 504506 698058 504742 698294
rect 504826 698058 505062 698294
rect 504506 662378 504742 662614
rect 504826 662378 505062 662614
rect 504506 662058 504742 662294
rect 504826 662058 505062 662294
rect 505906 709402 506142 709638
rect 506226 709402 506462 709638
rect 505906 709082 506142 709318
rect 506226 709082 506462 709318
rect 505906 676658 506142 676894
rect 506226 676658 506462 676894
rect 505906 676338 506142 676574
rect 506226 676338 506462 676574
rect 507306 706522 507542 706758
rect 507626 706522 507862 706758
rect 507306 706202 507542 706438
rect 507626 706202 507862 706438
rect 507306 690938 507542 691174
rect 507626 690938 507862 691174
rect 507306 690618 507542 690854
rect 507626 690618 507862 690854
rect 508706 705562 508942 705798
rect 509026 705562 509262 705798
rect 508706 705242 508942 705478
rect 509026 705242 509262 705478
rect 508706 669218 508942 669454
rect 509026 669218 509262 669454
rect 508706 668898 508942 669134
rect 509026 668898 509262 669134
rect 514746 710362 514982 710598
rect 515066 710362 515302 710598
rect 514746 710042 514982 710278
rect 515066 710042 515302 710278
rect 509626 680378 509862 680614
rect 509946 680378 510182 680614
rect 509626 680058 509862 680294
rect 509946 680058 510182 680294
rect 511026 708442 511262 708678
rect 511346 708442 511582 708678
rect 511026 708122 511262 708358
rect 511346 708122 511582 708358
rect 511026 694658 511262 694894
rect 511346 694658 511582 694894
rect 511026 694338 511262 694574
rect 511346 694338 511582 694574
rect 511026 658658 511262 658894
rect 511346 658658 511582 658894
rect 511026 658338 511262 658574
rect 511346 658338 511582 658574
rect 512426 707482 512662 707718
rect 512746 707482 512982 707718
rect 512426 707162 512662 707398
rect 512746 707162 512982 707398
rect 512426 672938 512662 673174
rect 512746 672938 512982 673174
rect 512426 672618 512662 672854
rect 512746 672618 512982 672854
rect 513826 704602 514062 704838
rect 514146 704602 514382 704838
rect 513826 704282 514062 704518
rect 514146 704282 514382 704518
rect 513826 687218 514062 687454
rect 514146 687218 514382 687454
rect 513826 686898 514062 687134
rect 514146 686898 514382 687134
rect 519866 711322 520102 711558
rect 520186 711322 520422 711558
rect 519866 711002 520102 711238
rect 520186 711002 520422 711238
rect 514746 698378 514982 698614
rect 515066 698378 515302 698614
rect 514746 698058 514982 698294
rect 515066 698058 515302 698294
rect 514746 662378 514982 662614
rect 515066 662378 515302 662614
rect 514746 662058 514982 662294
rect 515066 662058 515302 662294
rect 516146 709402 516382 709638
rect 516466 709402 516702 709638
rect 516146 709082 516382 709318
rect 516466 709082 516702 709318
rect 516146 676658 516382 676894
rect 516466 676658 516702 676894
rect 516146 676338 516382 676574
rect 516466 676338 516702 676574
rect 517546 706522 517782 706758
rect 517866 706522 518102 706758
rect 517546 706202 517782 706438
rect 517866 706202 518102 706438
rect 517546 690938 517782 691174
rect 517866 690938 518102 691174
rect 517546 690618 517782 690854
rect 517866 690618 518102 690854
rect 518946 705562 519182 705798
rect 519266 705562 519502 705798
rect 518946 705242 519182 705478
rect 519266 705242 519502 705478
rect 518946 669218 519182 669454
rect 519266 669218 519502 669454
rect 518946 668898 519182 669134
rect 519266 668898 519502 669134
rect 524986 710362 525222 710598
rect 525306 710362 525542 710598
rect 524986 710042 525222 710278
rect 525306 710042 525542 710278
rect 519866 680378 520102 680614
rect 520186 680378 520422 680614
rect 519866 680058 520102 680294
rect 520186 680058 520422 680294
rect 521266 708442 521502 708678
rect 521586 708442 521822 708678
rect 521266 708122 521502 708358
rect 521586 708122 521822 708358
rect 521266 694658 521502 694894
rect 521586 694658 521822 694894
rect 521266 694338 521502 694574
rect 521586 694338 521822 694574
rect 521266 658658 521502 658894
rect 521586 658658 521822 658894
rect 521266 658338 521502 658574
rect 521586 658338 521822 658574
rect 522666 707482 522902 707718
rect 522986 707482 523222 707718
rect 522666 707162 522902 707398
rect 522986 707162 523222 707398
rect 522666 672938 522902 673174
rect 522986 672938 523222 673174
rect 522666 672618 522902 672854
rect 522986 672618 523222 672854
rect 524066 704602 524302 704838
rect 524386 704602 524622 704838
rect 524066 704282 524302 704518
rect 524386 704282 524622 704518
rect 524066 687218 524302 687454
rect 524386 687218 524622 687454
rect 524066 686898 524302 687134
rect 524386 686898 524622 687134
rect 530106 711322 530342 711558
rect 530426 711322 530662 711558
rect 530106 711002 530342 711238
rect 530426 711002 530662 711238
rect 524986 698378 525222 698614
rect 525306 698378 525542 698614
rect 524986 698058 525222 698294
rect 525306 698058 525542 698294
rect 524986 662378 525222 662614
rect 525306 662378 525542 662614
rect 524986 662058 525222 662294
rect 525306 662058 525542 662294
rect 526386 709402 526622 709638
rect 526706 709402 526942 709638
rect 526386 709082 526622 709318
rect 526706 709082 526942 709318
rect 526386 676658 526622 676894
rect 526706 676658 526942 676894
rect 526386 676338 526622 676574
rect 526706 676338 526942 676574
rect 527786 706522 528022 706758
rect 528106 706522 528342 706758
rect 527786 706202 528022 706438
rect 528106 706202 528342 706438
rect 527786 690938 528022 691174
rect 528106 690938 528342 691174
rect 527786 690618 528022 690854
rect 528106 690618 528342 690854
rect 529186 705562 529422 705798
rect 529506 705562 529742 705798
rect 529186 705242 529422 705478
rect 529506 705242 529742 705478
rect 529186 669218 529422 669454
rect 529506 669218 529742 669454
rect 529186 668898 529422 669134
rect 529506 668898 529742 669134
rect 535226 710362 535462 710598
rect 535546 710362 535782 710598
rect 535226 710042 535462 710278
rect 535546 710042 535782 710278
rect 530106 680378 530342 680614
rect 530426 680378 530662 680614
rect 530106 680058 530342 680294
rect 530426 680058 530662 680294
rect 531506 708442 531742 708678
rect 531826 708442 532062 708678
rect 531506 708122 531742 708358
rect 531826 708122 532062 708358
rect 531506 694658 531742 694894
rect 531826 694658 532062 694894
rect 531506 694338 531742 694574
rect 531826 694338 532062 694574
rect 531506 658658 531742 658894
rect 531826 658658 532062 658894
rect 531506 658338 531742 658574
rect 531826 658338 532062 658574
rect 532906 707482 533142 707718
rect 533226 707482 533462 707718
rect 532906 707162 533142 707398
rect 533226 707162 533462 707398
rect 532906 672938 533142 673174
rect 533226 672938 533462 673174
rect 532906 672618 533142 672854
rect 533226 672618 533462 672854
rect 534306 704602 534542 704838
rect 534626 704602 534862 704838
rect 534306 704282 534542 704518
rect 534626 704282 534862 704518
rect 534306 687218 534542 687454
rect 534626 687218 534862 687454
rect 534306 686898 534542 687134
rect 534626 686898 534862 687134
rect 540346 711322 540582 711558
rect 540666 711322 540902 711558
rect 540346 711002 540582 711238
rect 540666 711002 540902 711238
rect 535226 698378 535462 698614
rect 535546 698378 535782 698614
rect 535226 698058 535462 698294
rect 535546 698058 535782 698294
rect 535226 662378 535462 662614
rect 535546 662378 535782 662614
rect 535226 662058 535462 662294
rect 535546 662058 535782 662294
rect 536626 709402 536862 709638
rect 536946 709402 537182 709638
rect 536626 709082 536862 709318
rect 536946 709082 537182 709318
rect 536626 676658 536862 676894
rect 536946 676658 537182 676894
rect 536626 676338 536862 676574
rect 536946 676338 537182 676574
rect 538026 706522 538262 706758
rect 538346 706522 538582 706758
rect 538026 706202 538262 706438
rect 538346 706202 538582 706438
rect 538026 690938 538262 691174
rect 538346 690938 538582 691174
rect 538026 690618 538262 690854
rect 538346 690618 538582 690854
rect 539426 705562 539662 705798
rect 539746 705562 539982 705798
rect 539426 705242 539662 705478
rect 539746 705242 539982 705478
rect 539426 669218 539662 669454
rect 539746 669218 539982 669454
rect 539426 668898 539662 669134
rect 539746 668898 539982 669134
rect 545466 710362 545702 710598
rect 545786 710362 546022 710598
rect 545466 710042 545702 710278
rect 545786 710042 546022 710278
rect 540346 680378 540582 680614
rect 540666 680378 540902 680614
rect 540346 680058 540582 680294
rect 540666 680058 540902 680294
rect 541746 708442 541982 708678
rect 542066 708442 542302 708678
rect 541746 708122 541982 708358
rect 542066 708122 542302 708358
rect 541746 694658 541982 694894
rect 542066 694658 542302 694894
rect 541746 694338 541982 694574
rect 542066 694338 542302 694574
rect 541746 658658 541982 658894
rect 542066 658658 542302 658894
rect 541746 658338 541982 658574
rect 542066 658338 542302 658574
rect 15786 654938 16022 655174
rect 16106 654938 16342 655174
rect 15786 654618 16022 654854
rect 16106 654618 16342 654854
rect 23330 651218 23566 651454
rect 23330 650898 23566 651134
rect 33570 651218 33806 651454
rect 33570 650898 33806 651134
rect 43810 651218 44046 651454
rect 43810 650898 44046 651134
rect 54050 651218 54286 651454
rect 54050 650898 54286 651134
rect 64290 651218 64526 651454
rect 64290 650898 64526 651134
rect 74530 651218 74766 651454
rect 74530 650898 74766 651134
rect 84770 651218 85006 651454
rect 84770 650898 85006 651134
rect 95010 651218 95246 651454
rect 95010 650898 95246 651134
rect 105250 651218 105486 651454
rect 105250 650898 105486 651134
rect 115490 651218 115726 651454
rect 115490 650898 115726 651134
rect 125730 651218 125966 651454
rect 125730 650898 125966 651134
rect 135970 651218 136206 651454
rect 135970 650898 136206 651134
rect 146210 651218 146446 651454
rect 146210 650898 146446 651134
rect 156450 651218 156686 651454
rect 156450 650898 156686 651134
rect 166690 651218 166926 651454
rect 166690 650898 166926 651134
rect 176930 651218 177166 651454
rect 176930 650898 177166 651134
rect 187170 651218 187406 651454
rect 187170 650898 187406 651134
rect 197410 651218 197646 651454
rect 197410 650898 197646 651134
rect 207650 651218 207886 651454
rect 207650 650898 207886 651134
rect 217890 651218 218126 651454
rect 217890 650898 218126 651134
rect 228130 651218 228366 651454
rect 228130 650898 228366 651134
rect 238370 651218 238606 651454
rect 238370 650898 238606 651134
rect 248610 651218 248846 651454
rect 248610 650898 248846 651134
rect 258850 651218 259086 651454
rect 258850 650898 259086 651134
rect 269090 651218 269326 651454
rect 269090 650898 269326 651134
rect 279330 651218 279566 651454
rect 279330 650898 279566 651134
rect 289570 651218 289806 651454
rect 289570 650898 289806 651134
rect 299810 651218 300046 651454
rect 299810 650898 300046 651134
rect 310050 651218 310286 651454
rect 310050 650898 310286 651134
rect 320290 651218 320526 651454
rect 320290 650898 320526 651134
rect 330530 651218 330766 651454
rect 330530 650898 330766 651134
rect 340770 651218 341006 651454
rect 340770 650898 341006 651134
rect 351010 651218 351246 651454
rect 351010 650898 351246 651134
rect 361250 651218 361486 651454
rect 361250 650898 361486 651134
rect 371490 651218 371726 651454
rect 371490 650898 371726 651134
rect 381730 651218 381966 651454
rect 381730 650898 381966 651134
rect 391970 651218 392206 651454
rect 391970 650898 392206 651134
rect 402210 651218 402446 651454
rect 402210 650898 402446 651134
rect 412450 651218 412686 651454
rect 412450 650898 412686 651134
rect 422690 651218 422926 651454
rect 422690 650898 422926 651134
rect 432930 651218 433166 651454
rect 432930 650898 433166 651134
rect 443170 651218 443406 651454
rect 443170 650898 443406 651134
rect 453410 651218 453646 651454
rect 453410 650898 453646 651134
rect 463650 651218 463886 651454
rect 463650 650898 463886 651134
rect 473890 651218 474126 651454
rect 473890 650898 474126 651134
rect 484130 651218 484366 651454
rect 484130 650898 484366 651134
rect 494370 651218 494606 651454
rect 494370 650898 494606 651134
rect 504610 651218 504846 651454
rect 504610 650898 504846 651134
rect 514850 651218 515086 651454
rect 514850 650898 515086 651134
rect 525090 651218 525326 651454
rect 525090 650898 525326 651134
rect 535330 651218 535566 651454
rect 535330 650898 535566 651134
rect 28450 633218 28686 633454
rect 28450 632898 28686 633134
rect 38690 633218 38926 633454
rect 38690 632898 38926 633134
rect 48930 633218 49166 633454
rect 48930 632898 49166 633134
rect 59170 633218 59406 633454
rect 59170 632898 59406 633134
rect 69410 633218 69646 633454
rect 69410 632898 69646 633134
rect 79650 633218 79886 633454
rect 79650 632898 79886 633134
rect 89890 633218 90126 633454
rect 89890 632898 90126 633134
rect 100130 633218 100366 633454
rect 100130 632898 100366 633134
rect 110370 633218 110606 633454
rect 110370 632898 110606 633134
rect 120610 633218 120846 633454
rect 120610 632898 120846 633134
rect 130850 633218 131086 633454
rect 130850 632898 131086 633134
rect 141090 633218 141326 633454
rect 141090 632898 141326 633134
rect 151330 633218 151566 633454
rect 151330 632898 151566 633134
rect 161570 633218 161806 633454
rect 161570 632898 161806 633134
rect 171810 633218 172046 633454
rect 171810 632898 172046 633134
rect 182050 633218 182286 633454
rect 182050 632898 182286 633134
rect 192290 633218 192526 633454
rect 192290 632898 192526 633134
rect 202530 633218 202766 633454
rect 202530 632898 202766 633134
rect 212770 633218 213006 633454
rect 212770 632898 213006 633134
rect 223010 633218 223246 633454
rect 223010 632898 223246 633134
rect 233250 633218 233486 633454
rect 233250 632898 233486 633134
rect 243490 633218 243726 633454
rect 243490 632898 243726 633134
rect 253730 633218 253966 633454
rect 253730 632898 253966 633134
rect 263970 633218 264206 633454
rect 263970 632898 264206 633134
rect 274210 633218 274446 633454
rect 274210 632898 274446 633134
rect 284450 633218 284686 633454
rect 284450 632898 284686 633134
rect 294690 633218 294926 633454
rect 294690 632898 294926 633134
rect 304930 633218 305166 633454
rect 304930 632898 305166 633134
rect 315170 633218 315406 633454
rect 315170 632898 315406 633134
rect 325410 633218 325646 633454
rect 325410 632898 325646 633134
rect 335650 633218 335886 633454
rect 335650 632898 335886 633134
rect 345890 633218 346126 633454
rect 345890 632898 346126 633134
rect 356130 633218 356366 633454
rect 356130 632898 356366 633134
rect 366370 633218 366606 633454
rect 366370 632898 366606 633134
rect 376610 633218 376846 633454
rect 376610 632898 376846 633134
rect 386850 633218 387086 633454
rect 386850 632898 387086 633134
rect 397090 633218 397326 633454
rect 397090 632898 397326 633134
rect 407330 633218 407566 633454
rect 407330 632898 407566 633134
rect 417570 633218 417806 633454
rect 417570 632898 417806 633134
rect 427810 633218 428046 633454
rect 427810 632898 428046 633134
rect 438050 633218 438286 633454
rect 438050 632898 438286 633134
rect 448290 633218 448526 633454
rect 448290 632898 448526 633134
rect 458530 633218 458766 633454
rect 458530 632898 458766 633134
rect 468770 633218 469006 633454
rect 468770 632898 469006 633134
rect 479010 633218 479246 633454
rect 479010 632898 479246 633134
rect 489250 633218 489486 633454
rect 489250 632898 489486 633134
rect 499490 633218 499726 633454
rect 499490 632898 499726 633134
rect 509730 633218 509966 633454
rect 509730 632898 509966 633134
rect 519970 633218 520206 633454
rect 519970 632898 520206 633134
rect 530210 633218 530446 633454
rect 530210 632898 530446 633134
rect 15786 618938 16022 619174
rect 16106 618938 16342 619174
rect 15786 618618 16022 618854
rect 16106 618618 16342 618854
rect 541746 622658 541982 622894
rect 542066 622658 542302 622894
rect 541746 622338 541982 622574
rect 542066 622338 542302 622574
rect 23330 615218 23566 615454
rect 23330 614898 23566 615134
rect 33570 615218 33806 615454
rect 33570 614898 33806 615134
rect 43810 615218 44046 615454
rect 43810 614898 44046 615134
rect 54050 615218 54286 615454
rect 54050 614898 54286 615134
rect 64290 615218 64526 615454
rect 64290 614898 64526 615134
rect 74530 615218 74766 615454
rect 74530 614898 74766 615134
rect 84770 615218 85006 615454
rect 84770 614898 85006 615134
rect 95010 615218 95246 615454
rect 95010 614898 95246 615134
rect 105250 615218 105486 615454
rect 105250 614898 105486 615134
rect 115490 615218 115726 615454
rect 115490 614898 115726 615134
rect 125730 615218 125966 615454
rect 125730 614898 125966 615134
rect 135970 615218 136206 615454
rect 135970 614898 136206 615134
rect 146210 615218 146446 615454
rect 146210 614898 146446 615134
rect 156450 615218 156686 615454
rect 156450 614898 156686 615134
rect 166690 615218 166926 615454
rect 166690 614898 166926 615134
rect 176930 615218 177166 615454
rect 176930 614898 177166 615134
rect 187170 615218 187406 615454
rect 187170 614898 187406 615134
rect 197410 615218 197646 615454
rect 197410 614898 197646 615134
rect 207650 615218 207886 615454
rect 207650 614898 207886 615134
rect 217890 615218 218126 615454
rect 217890 614898 218126 615134
rect 228130 615218 228366 615454
rect 228130 614898 228366 615134
rect 238370 615218 238606 615454
rect 238370 614898 238606 615134
rect 248610 615218 248846 615454
rect 248610 614898 248846 615134
rect 258850 615218 259086 615454
rect 258850 614898 259086 615134
rect 269090 615218 269326 615454
rect 269090 614898 269326 615134
rect 279330 615218 279566 615454
rect 279330 614898 279566 615134
rect 289570 615218 289806 615454
rect 289570 614898 289806 615134
rect 299810 615218 300046 615454
rect 299810 614898 300046 615134
rect 310050 615218 310286 615454
rect 310050 614898 310286 615134
rect 320290 615218 320526 615454
rect 320290 614898 320526 615134
rect 330530 615218 330766 615454
rect 330530 614898 330766 615134
rect 340770 615218 341006 615454
rect 340770 614898 341006 615134
rect 351010 615218 351246 615454
rect 351010 614898 351246 615134
rect 361250 615218 361486 615454
rect 361250 614898 361486 615134
rect 371490 615218 371726 615454
rect 371490 614898 371726 615134
rect 381730 615218 381966 615454
rect 381730 614898 381966 615134
rect 391970 615218 392206 615454
rect 391970 614898 392206 615134
rect 402210 615218 402446 615454
rect 402210 614898 402446 615134
rect 412450 615218 412686 615454
rect 412450 614898 412686 615134
rect 422690 615218 422926 615454
rect 422690 614898 422926 615134
rect 432930 615218 433166 615454
rect 432930 614898 433166 615134
rect 443170 615218 443406 615454
rect 443170 614898 443406 615134
rect 453410 615218 453646 615454
rect 453410 614898 453646 615134
rect 463650 615218 463886 615454
rect 463650 614898 463886 615134
rect 473890 615218 474126 615454
rect 473890 614898 474126 615134
rect 484130 615218 484366 615454
rect 484130 614898 484366 615134
rect 494370 615218 494606 615454
rect 494370 614898 494606 615134
rect 504610 615218 504846 615454
rect 504610 614898 504846 615134
rect 514850 615218 515086 615454
rect 514850 614898 515086 615134
rect 525090 615218 525326 615454
rect 525090 614898 525326 615134
rect 535330 615218 535566 615454
rect 535330 614898 535566 615134
rect 28450 597218 28686 597454
rect 28450 596898 28686 597134
rect 38690 597218 38926 597454
rect 38690 596898 38926 597134
rect 48930 597218 49166 597454
rect 48930 596898 49166 597134
rect 59170 597218 59406 597454
rect 59170 596898 59406 597134
rect 69410 597218 69646 597454
rect 69410 596898 69646 597134
rect 79650 597218 79886 597454
rect 79650 596898 79886 597134
rect 89890 597218 90126 597454
rect 89890 596898 90126 597134
rect 100130 597218 100366 597454
rect 100130 596898 100366 597134
rect 110370 597218 110606 597454
rect 110370 596898 110606 597134
rect 120610 597218 120846 597454
rect 120610 596898 120846 597134
rect 130850 597218 131086 597454
rect 130850 596898 131086 597134
rect 141090 597218 141326 597454
rect 141090 596898 141326 597134
rect 151330 597218 151566 597454
rect 151330 596898 151566 597134
rect 161570 597218 161806 597454
rect 161570 596898 161806 597134
rect 171810 597218 172046 597454
rect 171810 596898 172046 597134
rect 182050 597218 182286 597454
rect 182050 596898 182286 597134
rect 192290 597218 192526 597454
rect 192290 596898 192526 597134
rect 202530 597218 202766 597454
rect 202530 596898 202766 597134
rect 212770 597218 213006 597454
rect 212770 596898 213006 597134
rect 223010 597218 223246 597454
rect 223010 596898 223246 597134
rect 233250 597218 233486 597454
rect 233250 596898 233486 597134
rect 243490 597218 243726 597454
rect 243490 596898 243726 597134
rect 253730 597218 253966 597454
rect 253730 596898 253966 597134
rect 263970 597218 264206 597454
rect 263970 596898 264206 597134
rect 274210 597218 274446 597454
rect 274210 596898 274446 597134
rect 284450 597218 284686 597454
rect 284450 596898 284686 597134
rect 294690 597218 294926 597454
rect 294690 596898 294926 597134
rect 304930 597218 305166 597454
rect 304930 596898 305166 597134
rect 315170 597218 315406 597454
rect 315170 596898 315406 597134
rect 325410 597218 325646 597454
rect 325410 596898 325646 597134
rect 335650 597218 335886 597454
rect 335650 596898 335886 597134
rect 345890 597218 346126 597454
rect 345890 596898 346126 597134
rect 356130 597218 356366 597454
rect 356130 596898 356366 597134
rect 366370 597218 366606 597454
rect 366370 596898 366606 597134
rect 376610 597218 376846 597454
rect 376610 596898 376846 597134
rect 386850 597218 387086 597454
rect 386850 596898 387086 597134
rect 397090 597218 397326 597454
rect 397090 596898 397326 597134
rect 407330 597218 407566 597454
rect 407330 596898 407566 597134
rect 417570 597218 417806 597454
rect 417570 596898 417806 597134
rect 427810 597218 428046 597454
rect 427810 596898 428046 597134
rect 438050 597218 438286 597454
rect 438050 596898 438286 597134
rect 448290 597218 448526 597454
rect 448290 596898 448526 597134
rect 458530 597218 458766 597454
rect 458530 596898 458766 597134
rect 468770 597218 469006 597454
rect 468770 596898 469006 597134
rect 479010 597218 479246 597454
rect 479010 596898 479246 597134
rect 489250 597218 489486 597454
rect 489250 596898 489486 597134
rect 499490 597218 499726 597454
rect 499490 596898 499726 597134
rect 509730 597218 509966 597454
rect 509730 596898 509966 597134
rect 519970 597218 520206 597454
rect 519970 596898 520206 597134
rect 530210 597218 530446 597454
rect 530210 596898 530446 597134
rect 15786 582938 16022 583174
rect 16106 582938 16342 583174
rect 15786 582618 16022 582854
rect 16106 582618 16342 582854
rect 541746 586658 541982 586894
rect 542066 586658 542302 586894
rect 541746 586338 541982 586574
rect 542066 586338 542302 586574
rect 23330 579218 23566 579454
rect 23330 578898 23566 579134
rect 33570 579218 33806 579454
rect 33570 578898 33806 579134
rect 43810 579218 44046 579454
rect 43810 578898 44046 579134
rect 54050 579218 54286 579454
rect 54050 578898 54286 579134
rect 64290 579218 64526 579454
rect 64290 578898 64526 579134
rect 74530 579218 74766 579454
rect 74530 578898 74766 579134
rect 84770 579218 85006 579454
rect 84770 578898 85006 579134
rect 95010 579218 95246 579454
rect 95010 578898 95246 579134
rect 105250 579218 105486 579454
rect 105250 578898 105486 579134
rect 115490 579218 115726 579454
rect 115490 578898 115726 579134
rect 125730 579218 125966 579454
rect 125730 578898 125966 579134
rect 135970 579218 136206 579454
rect 135970 578898 136206 579134
rect 146210 579218 146446 579454
rect 146210 578898 146446 579134
rect 156450 579218 156686 579454
rect 156450 578898 156686 579134
rect 166690 579218 166926 579454
rect 166690 578898 166926 579134
rect 176930 579218 177166 579454
rect 176930 578898 177166 579134
rect 187170 579218 187406 579454
rect 187170 578898 187406 579134
rect 197410 579218 197646 579454
rect 197410 578898 197646 579134
rect 207650 579218 207886 579454
rect 207650 578898 207886 579134
rect 217890 579218 218126 579454
rect 217890 578898 218126 579134
rect 228130 579218 228366 579454
rect 228130 578898 228366 579134
rect 238370 579218 238606 579454
rect 238370 578898 238606 579134
rect 248610 579218 248846 579454
rect 248610 578898 248846 579134
rect 258850 579218 259086 579454
rect 258850 578898 259086 579134
rect 269090 579218 269326 579454
rect 269090 578898 269326 579134
rect 279330 579218 279566 579454
rect 279330 578898 279566 579134
rect 289570 579218 289806 579454
rect 289570 578898 289806 579134
rect 299810 579218 300046 579454
rect 299810 578898 300046 579134
rect 310050 579218 310286 579454
rect 310050 578898 310286 579134
rect 320290 579218 320526 579454
rect 320290 578898 320526 579134
rect 330530 579218 330766 579454
rect 330530 578898 330766 579134
rect 340770 579218 341006 579454
rect 340770 578898 341006 579134
rect 351010 579218 351246 579454
rect 351010 578898 351246 579134
rect 361250 579218 361486 579454
rect 361250 578898 361486 579134
rect 371490 579218 371726 579454
rect 371490 578898 371726 579134
rect 381730 579218 381966 579454
rect 381730 578898 381966 579134
rect 391970 579218 392206 579454
rect 391970 578898 392206 579134
rect 402210 579218 402446 579454
rect 402210 578898 402446 579134
rect 412450 579218 412686 579454
rect 412450 578898 412686 579134
rect 422690 579218 422926 579454
rect 422690 578898 422926 579134
rect 432930 579218 433166 579454
rect 432930 578898 433166 579134
rect 443170 579218 443406 579454
rect 443170 578898 443406 579134
rect 453410 579218 453646 579454
rect 453410 578898 453646 579134
rect 463650 579218 463886 579454
rect 463650 578898 463886 579134
rect 473890 579218 474126 579454
rect 473890 578898 474126 579134
rect 484130 579218 484366 579454
rect 484130 578898 484366 579134
rect 494370 579218 494606 579454
rect 494370 578898 494606 579134
rect 504610 579218 504846 579454
rect 504610 578898 504846 579134
rect 514850 579218 515086 579454
rect 514850 578898 515086 579134
rect 525090 579218 525326 579454
rect 525090 578898 525326 579134
rect 535330 579218 535566 579454
rect 535330 578898 535566 579134
rect 28450 561218 28686 561454
rect 28450 560898 28686 561134
rect 38690 561218 38926 561454
rect 38690 560898 38926 561134
rect 48930 561218 49166 561454
rect 48930 560898 49166 561134
rect 59170 561218 59406 561454
rect 59170 560898 59406 561134
rect 69410 561218 69646 561454
rect 69410 560898 69646 561134
rect 79650 561218 79886 561454
rect 79650 560898 79886 561134
rect 89890 561218 90126 561454
rect 89890 560898 90126 561134
rect 100130 561218 100366 561454
rect 100130 560898 100366 561134
rect 110370 561218 110606 561454
rect 110370 560898 110606 561134
rect 120610 561218 120846 561454
rect 120610 560898 120846 561134
rect 130850 561218 131086 561454
rect 130850 560898 131086 561134
rect 141090 561218 141326 561454
rect 141090 560898 141326 561134
rect 151330 561218 151566 561454
rect 151330 560898 151566 561134
rect 161570 561218 161806 561454
rect 161570 560898 161806 561134
rect 171810 561218 172046 561454
rect 171810 560898 172046 561134
rect 182050 561218 182286 561454
rect 182050 560898 182286 561134
rect 192290 561218 192526 561454
rect 192290 560898 192526 561134
rect 202530 561218 202766 561454
rect 202530 560898 202766 561134
rect 212770 561218 213006 561454
rect 212770 560898 213006 561134
rect 223010 561218 223246 561454
rect 223010 560898 223246 561134
rect 233250 561218 233486 561454
rect 233250 560898 233486 561134
rect 243490 561218 243726 561454
rect 243490 560898 243726 561134
rect 253730 561218 253966 561454
rect 253730 560898 253966 561134
rect 263970 561218 264206 561454
rect 263970 560898 264206 561134
rect 274210 561218 274446 561454
rect 274210 560898 274446 561134
rect 284450 561218 284686 561454
rect 284450 560898 284686 561134
rect 294690 561218 294926 561454
rect 294690 560898 294926 561134
rect 304930 561218 305166 561454
rect 304930 560898 305166 561134
rect 315170 561218 315406 561454
rect 315170 560898 315406 561134
rect 325410 561218 325646 561454
rect 325410 560898 325646 561134
rect 335650 561218 335886 561454
rect 335650 560898 335886 561134
rect 345890 561218 346126 561454
rect 345890 560898 346126 561134
rect 356130 561218 356366 561454
rect 356130 560898 356366 561134
rect 366370 561218 366606 561454
rect 366370 560898 366606 561134
rect 376610 561218 376846 561454
rect 376610 560898 376846 561134
rect 386850 561218 387086 561454
rect 386850 560898 387086 561134
rect 397090 561218 397326 561454
rect 397090 560898 397326 561134
rect 407330 561218 407566 561454
rect 407330 560898 407566 561134
rect 417570 561218 417806 561454
rect 417570 560898 417806 561134
rect 427810 561218 428046 561454
rect 427810 560898 428046 561134
rect 438050 561218 438286 561454
rect 438050 560898 438286 561134
rect 448290 561218 448526 561454
rect 448290 560898 448526 561134
rect 458530 561218 458766 561454
rect 458530 560898 458766 561134
rect 468770 561218 469006 561454
rect 468770 560898 469006 561134
rect 479010 561218 479246 561454
rect 479010 560898 479246 561134
rect 489250 561218 489486 561454
rect 489250 560898 489486 561134
rect 499490 561218 499726 561454
rect 499490 560898 499726 561134
rect 509730 561218 509966 561454
rect 509730 560898 509966 561134
rect 519970 561218 520206 561454
rect 519970 560898 520206 561134
rect 530210 561218 530446 561454
rect 530210 560898 530446 561134
rect 15786 546938 16022 547174
rect 16106 546938 16342 547174
rect 15786 546618 16022 546854
rect 16106 546618 16342 546854
rect 541746 550658 541982 550894
rect 542066 550658 542302 550894
rect 541746 550338 541982 550574
rect 542066 550338 542302 550574
rect 23330 543218 23566 543454
rect 23330 542898 23566 543134
rect 33570 543218 33806 543454
rect 33570 542898 33806 543134
rect 43810 543218 44046 543454
rect 43810 542898 44046 543134
rect 54050 543218 54286 543454
rect 54050 542898 54286 543134
rect 64290 543218 64526 543454
rect 64290 542898 64526 543134
rect 74530 543218 74766 543454
rect 74530 542898 74766 543134
rect 84770 543218 85006 543454
rect 84770 542898 85006 543134
rect 95010 543218 95246 543454
rect 95010 542898 95246 543134
rect 105250 543218 105486 543454
rect 105250 542898 105486 543134
rect 115490 543218 115726 543454
rect 115490 542898 115726 543134
rect 125730 543218 125966 543454
rect 125730 542898 125966 543134
rect 135970 543218 136206 543454
rect 135970 542898 136206 543134
rect 146210 543218 146446 543454
rect 146210 542898 146446 543134
rect 156450 543218 156686 543454
rect 156450 542898 156686 543134
rect 166690 543218 166926 543454
rect 166690 542898 166926 543134
rect 176930 543218 177166 543454
rect 176930 542898 177166 543134
rect 187170 543218 187406 543454
rect 187170 542898 187406 543134
rect 197410 543218 197646 543454
rect 197410 542898 197646 543134
rect 207650 543218 207886 543454
rect 207650 542898 207886 543134
rect 217890 543218 218126 543454
rect 217890 542898 218126 543134
rect 228130 543218 228366 543454
rect 228130 542898 228366 543134
rect 238370 543218 238606 543454
rect 238370 542898 238606 543134
rect 248610 543218 248846 543454
rect 248610 542898 248846 543134
rect 258850 543218 259086 543454
rect 258850 542898 259086 543134
rect 269090 543218 269326 543454
rect 269090 542898 269326 543134
rect 279330 543218 279566 543454
rect 279330 542898 279566 543134
rect 289570 543218 289806 543454
rect 289570 542898 289806 543134
rect 299810 543218 300046 543454
rect 299810 542898 300046 543134
rect 310050 543218 310286 543454
rect 310050 542898 310286 543134
rect 320290 543218 320526 543454
rect 320290 542898 320526 543134
rect 330530 543218 330766 543454
rect 330530 542898 330766 543134
rect 340770 543218 341006 543454
rect 340770 542898 341006 543134
rect 351010 543218 351246 543454
rect 351010 542898 351246 543134
rect 361250 543218 361486 543454
rect 361250 542898 361486 543134
rect 371490 543218 371726 543454
rect 371490 542898 371726 543134
rect 381730 543218 381966 543454
rect 381730 542898 381966 543134
rect 391970 543218 392206 543454
rect 391970 542898 392206 543134
rect 402210 543218 402446 543454
rect 402210 542898 402446 543134
rect 412450 543218 412686 543454
rect 412450 542898 412686 543134
rect 422690 543218 422926 543454
rect 422690 542898 422926 543134
rect 432930 543218 433166 543454
rect 432930 542898 433166 543134
rect 443170 543218 443406 543454
rect 443170 542898 443406 543134
rect 453410 543218 453646 543454
rect 453410 542898 453646 543134
rect 463650 543218 463886 543454
rect 463650 542898 463886 543134
rect 473890 543218 474126 543454
rect 473890 542898 474126 543134
rect 484130 543218 484366 543454
rect 484130 542898 484366 543134
rect 494370 543218 494606 543454
rect 494370 542898 494606 543134
rect 504610 543218 504846 543454
rect 504610 542898 504846 543134
rect 514850 543218 515086 543454
rect 514850 542898 515086 543134
rect 525090 543218 525326 543454
rect 525090 542898 525326 543134
rect 535330 543218 535566 543454
rect 535330 542898 535566 543134
rect 28450 525218 28686 525454
rect 28450 524898 28686 525134
rect 38690 525218 38926 525454
rect 38690 524898 38926 525134
rect 48930 525218 49166 525454
rect 48930 524898 49166 525134
rect 59170 525218 59406 525454
rect 59170 524898 59406 525134
rect 69410 525218 69646 525454
rect 69410 524898 69646 525134
rect 79650 525218 79886 525454
rect 79650 524898 79886 525134
rect 89890 525218 90126 525454
rect 89890 524898 90126 525134
rect 100130 525218 100366 525454
rect 100130 524898 100366 525134
rect 110370 525218 110606 525454
rect 110370 524898 110606 525134
rect 120610 525218 120846 525454
rect 120610 524898 120846 525134
rect 130850 525218 131086 525454
rect 130850 524898 131086 525134
rect 141090 525218 141326 525454
rect 141090 524898 141326 525134
rect 151330 525218 151566 525454
rect 151330 524898 151566 525134
rect 161570 525218 161806 525454
rect 161570 524898 161806 525134
rect 171810 525218 172046 525454
rect 171810 524898 172046 525134
rect 182050 525218 182286 525454
rect 182050 524898 182286 525134
rect 192290 525218 192526 525454
rect 192290 524898 192526 525134
rect 202530 525218 202766 525454
rect 202530 524898 202766 525134
rect 212770 525218 213006 525454
rect 212770 524898 213006 525134
rect 223010 525218 223246 525454
rect 223010 524898 223246 525134
rect 233250 525218 233486 525454
rect 233250 524898 233486 525134
rect 243490 525218 243726 525454
rect 243490 524898 243726 525134
rect 253730 525218 253966 525454
rect 253730 524898 253966 525134
rect 263970 525218 264206 525454
rect 263970 524898 264206 525134
rect 274210 525218 274446 525454
rect 274210 524898 274446 525134
rect 284450 525218 284686 525454
rect 284450 524898 284686 525134
rect 294690 525218 294926 525454
rect 294690 524898 294926 525134
rect 304930 525218 305166 525454
rect 304930 524898 305166 525134
rect 315170 525218 315406 525454
rect 315170 524898 315406 525134
rect 325410 525218 325646 525454
rect 325410 524898 325646 525134
rect 335650 525218 335886 525454
rect 335650 524898 335886 525134
rect 345890 525218 346126 525454
rect 345890 524898 346126 525134
rect 356130 525218 356366 525454
rect 356130 524898 356366 525134
rect 366370 525218 366606 525454
rect 366370 524898 366606 525134
rect 376610 525218 376846 525454
rect 376610 524898 376846 525134
rect 386850 525218 387086 525454
rect 386850 524898 387086 525134
rect 397090 525218 397326 525454
rect 397090 524898 397326 525134
rect 407330 525218 407566 525454
rect 407330 524898 407566 525134
rect 417570 525218 417806 525454
rect 417570 524898 417806 525134
rect 427810 525218 428046 525454
rect 427810 524898 428046 525134
rect 438050 525218 438286 525454
rect 438050 524898 438286 525134
rect 448290 525218 448526 525454
rect 448290 524898 448526 525134
rect 458530 525218 458766 525454
rect 458530 524898 458766 525134
rect 468770 525218 469006 525454
rect 468770 524898 469006 525134
rect 479010 525218 479246 525454
rect 479010 524898 479246 525134
rect 489250 525218 489486 525454
rect 489250 524898 489486 525134
rect 499490 525218 499726 525454
rect 499490 524898 499726 525134
rect 509730 525218 509966 525454
rect 509730 524898 509966 525134
rect 519970 525218 520206 525454
rect 519970 524898 520206 525134
rect 530210 525218 530446 525454
rect 530210 524898 530446 525134
rect 15786 510938 16022 511174
rect 16106 510938 16342 511174
rect 15786 510618 16022 510854
rect 16106 510618 16342 510854
rect 541746 514658 541982 514894
rect 542066 514658 542302 514894
rect 541746 514338 541982 514574
rect 542066 514338 542302 514574
rect 23330 507218 23566 507454
rect 23330 506898 23566 507134
rect 33570 507218 33806 507454
rect 33570 506898 33806 507134
rect 43810 507218 44046 507454
rect 43810 506898 44046 507134
rect 54050 507218 54286 507454
rect 54050 506898 54286 507134
rect 64290 507218 64526 507454
rect 64290 506898 64526 507134
rect 74530 507218 74766 507454
rect 74530 506898 74766 507134
rect 84770 507218 85006 507454
rect 84770 506898 85006 507134
rect 95010 507218 95246 507454
rect 95010 506898 95246 507134
rect 105250 507218 105486 507454
rect 105250 506898 105486 507134
rect 115490 507218 115726 507454
rect 115490 506898 115726 507134
rect 125730 507218 125966 507454
rect 125730 506898 125966 507134
rect 135970 507218 136206 507454
rect 135970 506898 136206 507134
rect 146210 507218 146446 507454
rect 146210 506898 146446 507134
rect 156450 507218 156686 507454
rect 156450 506898 156686 507134
rect 166690 507218 166926 507454
rect 166690 506898 166926 507134
rect 176930 507218 177166 507454
rect 176930 506898 177166 507134
rect 187170 507218 187406 507454
rect 187170 506898 187406 507134
rect 197410 507218 197646 507454
rect 197410 506898 197646 507134
rect 207650 507218 207886 507454
rect 207650 506898 207886 507134
rect 217890 507218 218126 507454
rect 217890 506898 218126 507134
rect 228130 507218 228366 507454
rect 228130 506898 228366 507134
rect 238370 507218 238606 507454
rect 238370 506898 238606 507134
rect 248610 507218 248846 507454
rect 248610 506898 248846 507134
rect 258850 507218 259086 507454
rect 258850 506898 259086 507134
rect 269090 507218 269326 507454
rect 269090 506898 269326 507134
rect 279330 507218 279566 507454
rect 279330 506898 279566 507134
rect 289570 507218 289806 507454
rect 289570 506898 289806 507134
rect 299810 507218 300046 507454
rect 299810 506898 300046 507134
rect 310050 507218 310286 507454
rect 310050 506898 310286 507134
rect 320290 507218 320526 507454
rect 320290 506898 320526 507134
rect 330530 507218 330766 507454
rect 330530 506898 330766 507134
rect 340770 507218 341006 507454
rect 340770 506898 341006 507134
rect 351010 507218 351246 507454
rect 351010 506898 351246 507134
rect 361250 507218 361486 507454
rect 361250 506898 361486 507134
rect 371490 507218 371726 507454
rect 371490 506898 371726 507134
rect 381730 507218 381966 507454
rect 381730 506898 381966 507134
rect 391970 507218 392206 507454
rect 391970 506898 392206 507134
rect 402210 507218 402446 507454
rect 402210 506898 402446 507134
rect 412450 507218 412686 507454
rect 412450 506898 412686 507134
rect 422690 507218 422926 507454
rect 422690 506898 422926 507134
rect 432930 507218 433166 507454
rect 432930 506898 433166 507134
rect 443170 507218 443406 507454
rect 443170 506898 443406 507134
rect 453410 507218 453646 507454
rect 453410 506898 453646 507134
rect 463650 507218 463886 507454
rect 463650 506898 463886 507134
rect 473890 507218 474126 507454
rect 473890 506898 474126 507134
rect 484130 507218 484366 507454
rect 484130 506898 484366 507134
rect 494370 507218 494606 507454
rect 494370 506898 494606 507134
rect 504610 507218 504846 507454
rect 504610 506898 504846 507134
rect 514850 507218 515086 507454
rect 514850 506898 515086 507134
rect 525090 507218 525326 507454
rect 525090 506898 525326 507134
rect 535330 507218 535566 507454
rect 535330 506898 535566 507134
rect 28450 489218 28686 489454
rect 28450 488898 28686 489134
rect 38690 489218 38926 489454
rect 38690 488898 38926 489134
rect 48930 489218 49166 489454
rect 48930 488898 49166 489134
rect 59170 489218 59406 489454
rect 59170 488898 59406 489134
rect 69410 489218 69646 489454
rect 69410 488898 69646 489134
rect 79650 489218 79886 489454
rect 79650 488898 79886 489134
rect 89890 489218 90126 489454
rect 89890 488898 90126 489134
rect 100130 489218 100366 489454
rect 100130 488898 100366 489134
rect 110370 489218 110606 489454
rect 110370 488898 110606 489134
rect 120610 489218 120846 489454
rect 120610 488898 120846 489134
rect 130850 489218 131086 489454
rect 130850 488898 131086 489134
rect 141090 489218 141326 489454
rect 141090 488898 141326 489134
rect 151330 489218 151566 489454
rect 151330 488898 151566 489134
rect 161570 489218 161806 489454
rect 161570 488898 161806 489134
rect 171810 489218 172046 489454
rect 171810 488898 172046 489134
rect 182050 489218 182286 489454
rect 182050 488898 182286 489134
rect 192290 489218 192526 489454
rect 192290 488898 192526 489134
rect 202530 489218 202766 489454
rect 202530 488898 202766 489134
rect 212770 489218 213006 489454
rect 212770 488898 213006 489134
rect 223010 489218 223246 489454
rect 223010 488898 223246 489134
rect 233250 489218 233486 489454
rect 233250 488898 233486 489134
rect 243490 489218 243726 489454
rect 243490 488898 243726 489134
rect 253730 489218 253966 489454
rect 253730 488898 253966 489134
rect 263970 489218 264206 489454
rect 263970 488898 264206 489134
rect 274210 489218 274446 489454
rect 274210 488898 274446 489134
rect 284450 489218 284686 489454
rect 284450 488898 284686 489134
rect 294690 489218 294926 489454
rect 294690 488898 294926 489134
rect 304930 489218 305166 489454
rect 304930 488898 305166 489134
rect 315170 489218 315406 489454
rect 315170 488898 315406 489134
rect 325410 489218 325646 489454
rect 325410 488898 325646 489134
rect 335650 489218 335886 489454
rect 335650 488898 335886 489134
rect 345890 489218 346126 489454
rect 345890 488898 346126 489134
rect 356130 489218 356366 489454
rect 356130 488898 356366 489134
rect 366370 489218 366606 489454
rect 366370 488898 366606 489134
rect 376610 489218 376846 489454
rect 376610 488898 376846 489134
rect 386850 489218 387086 489454
rect 386850 488898 387086 489134
rect 397090 489218 397326 489454
rect 397090 488898 397326 489134
rect 407330 489218 407566 489454
rect 407330 488898 407566 489134
rect 417570 489218 417806 489454
rect 417570 488898 417806 489134
rect 427810 489218 428046 489454
rect 427810 488898 428046 489134
rect 438050 489218 438286 489454
rect 438050 488898 438286 489134
rect 448290 489218 448526 489454
rect 448290 488898 448526 489134
rect 458530 489218 458766 489454
rect 458530 488898 458766 489134
rect 468770 489218 469006 489454
rect 468770 488898 469006 489134
rect 479010 489218 479246 489454
rect 479010 488898 479246 489134
rect 489250 489218 489486 489454
rect 489250 488898 489486 489134
rect 499490 489218 499726 489454
rect 499490 488898 499726 489134
rect 509730 489218 509966 489454
rect 509730 488898 509966 489134
rect 519970 489218 520206 489454
rect 519970 488898 520206 489134
rect 530210 489218 530446 489454
rect 530210 488898 530446 489134
rect 15786 474938 16022 475174
rect 16106 474938 16342 475174
rect 15786 474618 16022 474854
rect 16106 474618 16342 474854
rect 541746 478658 541982 478894
rect 542066 478658 542302 478894
rect 541746 478338 541982 478574
rect 542066 478338 542302 478574
rect 23330 471218 23566 471454
rect 23330 470898 23566 471134
rect 33570 471218 33806 471454
rect 33570 470898 33806 471134
rect 43810 471218 44046 471454
rect 43810 470898 44046 471134
rect 54050 471218 54286 471454
rect 54050 470898 54286 471134
rect 64290 471218 64526 471454
rect 64290 470898 64526 471134
rect 74530 471218 74766 471454
rect 74530 470898 74766 471134
rect 84770 471218 85006 471454
rect 84770 470898 85006 471134
rect 95010 471218 95246 471454
rect 95010 470898 95246 471134
rect 105250 471218 105486 471454
rect 105250 470898 105486 471134
rect 115490 471218 115726 471454
rect 115490 470898 115726 471134
rect 125730 471218 125966 471454
rect 125730 470898 125966 471134
rect 135970 471218 136206 471454
rect 135970 470898 136206 471134
rect 146210 471218 146446 471454
rect 146210 470898 146446 471134
rect 156450 471218 156686 471454
rect 156450 470898 156686 471134
rect 166690 471218 166926 471454
rect 166690 470898 166926 471134
rect 176930 471218 177166 471454
rect 176930 470898 177166 471134
rect 187170 471218 187406 471454
rect 187170 470898 187406 471134
rect 197410 471218 197646 471454
rect 197410 470898 197646 471134
rect 207650 471218 207886 471454
rect 207650 470898 207886 471134
rect 217890 471218 218126 471454
rect 217890 470898 218126 471134
rect 228130 471218 228366 471454
rect 228130 470898 228366 471134
rect 238370 471218 238606 471454
rect 238370 470898 238606 471134
rect 248610 471218 248846 471454
rect 248610 470898 248846 471134
rect 258850 471218 259086 471454
rect 258850 470898 259086 471134
rect 269090 471218 269326 471454
rect 269090 470898 269326 471134
rect 279330 471218 279566 471454
rect 279330 470898 279566 471134
rect 289570 471218 289806 471454
rect 289570 470898 289806 471134
rect 299810 471218 300046 471454
rect 299810 470898 300046 471134
rect 310050 471218 310286 471454
rect 310050 470898 310286 471134
rect 320290 471218 320526 471454
rect 320290 470898 320526 471134
rect 330530 471218 330766 471454
rect 330530 470898 330766 471134
rect 340770 471218 341006 471454
rect 340770 470898 341006 471134
rect 351010 471218 351246 471454
rect 351010 470898 351246 471134
rect 361250 471218 361486 471454
rect 361250 470898 361486 471134
rect 371490 471218 371726 471454
rect 371490 470898 371726 471134
rect 381730 471218 381966 471454
rect 381730 470898 381966 471134
rect 391970 471218 392206 471454
rect 391970 470898 392206 471134
rect 402210 471218 402446 471454
rect 402210 470898 402446 471134
rect 412450 471218 412686 471454
rect 412450 470898 412686 471134
rect 422690 471218 422926 471454
rect 422690 470898 422926 471134
rect 432930 471218 433166 471454
rect 432930 470898 433166 471134
rect 443170 471218 443406 471454
rect 443170 470898 443406 471134
rect 453410 471218 453646 471454
rect 453410 470898 453646 471134
rect 463650 471218 463886 471454
rect 463650 470898 463886 471134
rect 473890 471218 474126 471454
rect 473890 470898 474126 471134
rect 484130 471218 484366 471454
rect 484130 470898 484366 471134
rect 494370 471218 494606 471454
rect 494370 470898 494606 471134
rect 504610 471218 504846 471454
rect 504610 470898 504846 471134
rect 514850 471218 515086 471454
rect 514850 470898 515086 471134
rect 525090 471218 525326 471454
rect 525090 470898 525326 471134
rect 535330 471218 535566 471454
rect 535330 470898 535566 471134
rect 28450 453218 28686 453454
rect 28450 452898 28686 453134
rect 38690 453218 38926 453454
rect 38690 452898 38926 453134
rect 48930 453218 49166 453454
rect 48930 452898 49166 453134
rect 59170 453218 59406 453454
rect 59170 452898 59406 453134
rect 69410 453218 69646 453454
rect 69410 452898 69646 453134
rect 79650 453218 79886 453454
rect 79650 452898 79886 453134
rect 89890 453218 90126 453454
rect 89890 452898 90126 453134
rect 100130 453218 100366 453454
rect 100130 452898 100366 453134
rect 110370 453218 110606 453454
rect 110370 452898 110606 453134
rect 120610 453218 120846 453454
rect 120610 452898 120846 453134
rect 130850 453218 131086 453454
rect 130850 452898 131086 453134
rect 141090 453218 141326 453454
rect 141090 452898 141326 453134
rect 151330 453218 151566 453454
rect 151330 452898 151566 453134
rect 161570 453218 161806 453454
rect 161570 452898 161806 453134
rect 171810 453218 172046 453454
rect 171810 452898 172046 453134
rect 182050 453218 182286 453454
rect 182050 452898 182286 453134
rect 192290 453218 192526 453454
rect 192290 452898 192526 453134
rect 202530 453218 202766 453454
rect 202530 452898 202766 453134
rect 212770 453218 213006 453454
rect 212770 452898 213006 453134
rect 223010 453218 223246 453454
rect 223010 452898 223246 453134
rect 233250 453218 233486 453454
rect 233250 452898 233486 453134
rect 243490 453218 243726 453454
rect 243490 452898 243726 453134
rect 253730 453218 253966 453454
rect 253730 452898 253966 453134
rect 263970 453218 264206 453454
rect 263970 452898 264206 453134
rect 274210 453218 274446 453454
rect 274210 452898 274446 453134
rect 284450 453218 284686 453454
rect 284450 452898 284686 453134
rect 294690 453218 294926 453454
rect 294690 452898 294926 453134
rect 304930 453218 305166 453454
rect 304930 452898 305166 453134
rect 315170 453218 315406 453454
rect 315170 452898 315406 453134
rect 325410 453218 325646 453454
rect 325410 452898 325646 453134
rect 335650 453218 335886 453454
rect 335650 452898 335886 453134
rect 345890 453218 346126 453454
rect 345890 452898 346126 453134
rect 356130 453218 356366 453454
rect 356130 452898 356366 453134
rect 366370 453218 366606 453454
rect 366370 452898 366606 453134
rect 376610 453218 376846 453454
rect 376610 452898 376846 453134
rect 386850 453218 387086 453454
rect 386850 452898 387086 453134
rect 397090 453218 397326 453454
rect 397090 452898 397326 453134
rect 407330 453218 407566 453454
rect 407330 452898 407566 453134
rect 417570 453218 417806 453454
rect 417570 452898 417806 453134
rect 427810 453218 428046 453454
rect 427810 452898 428046 453134
rect 438050 453218 438286 453454
rect 438050 452898 438286 453134
rect 448290 453218 448526 453454
rect 448290 452898 448526 453134
rect 458530 453218 458766 453454
rect 458530 452898 458766 453134
rect 468770 453218 469006 453454
rect 468770 452898 469006 453134
rect 479010 453218 479246 453454
rect 479010 452898 479246 453134
rect 489250 453218 489486 453454
rect 489250 452898 489486 453134
rect 499490 453218 499726 453454
rect 499490 452898 499726 453134
rect 509730 453218 509966 453454
rect 509730 452898 509966 453134
rect 519970 453218 520206 453454
rect 519970 452898 520206 453134
rect 530210 453218 530446 453454
rect 530210 452898 530446 453134
rect 15786 438938 16022 439174
rect 16106 438938 16342 439174
rect 15786 438618 16022 438854
rect 16106 438618 16342 438854
rect 541746 442658 541982 442894
rect 542066 442658 542302 442894
rect 541746 442338 541982 442574
rect 542066 442338 542302 442574
rect 23330 435218 23566 435454
rect 23330 434898 23566 435134
rect 33570 435218 33806 435454
rect 33570 434898 33806 435134
rect 43810 435218 44046 435454
rect 43810 434898 44046 435134
rect 54050 435218 54286 435454
rect 54050 434898 54286 435134
rect 64290 435218 64526 435454
rect 64290 434898 64526 435134
rect 74530 435218 74766 435454
rect 74530 434898 74766 435134
rect 84770 435218 85006 435454
rect 84770 434898 85006 435134
rect 95010 435218 95246 435454
rect 95010 434898 95246 435134
rect 105250 435218 105486 435454
rect 105250 434898 105486 435134
rect 115490 435218 115726 435454
rect 115490 434898 115726 435134
rect 125730 435218 125966 435454
rect 125730 434898 125966 435134
rect 135970 435218 136206 435454
rect 135970 434898 136206 435134
rect 146210 435218 146446 435454
rect 146210 434898 146446 435134
rect 156450 435218 156686 435454
rect 156450 434898 156686 435134
rect 166690 435218 166926 435454
rect 166690 434898 166926 435134
rect 176930 435218 177166 435454
rect 176930 434898 177166 435134
rect 187170 435218 187406 435454
rect 187170 434898 187406 435134
rect 197410 435218 197646 435454
rect 197410 434898 197646 435134
rect 207650 435218 207886 435454
rect 207650 434898 207886 435134
rect 217890 435218 218126 435454
rect 217890 434898 218126 435134
rect 228130 435218 228366 435454
rect 228130 434898 228366 435134
rect 238370 435218 238606 435454
rect 238370 434898 238606 435134
rect 248610 435218 248846 435454
rect 248610 434898 248846 435134
rect 258850 435218 259086 435454
rect 258850 434898 259086 435134
rect 269090 435218 269326 435454
rect 269090 434898 269326 435134
rect 279330 435218 279566 435454
rect 279330 434898 279566 435134
rect 289570 435218 289806 435454
rect 289570 434898 289806 435134
rect 299810 435218 300046 435454
rect 299810 434898 300046 435134
rect 310050 435218 310286 435454
rect 310050 434898 310286 435134
rect 320290 435218 320526 435454
rect 320290 434898 320526 435134
rect 330530 435218 330766 435454
rect 330530 434898 330766 435134
rect 340770 435218 341006 435454
rect 340770 434898 341006 435134
rect 351010 435218 351246 435454
rect 351010 434898 351246 435134
rect 361250 435218 361486 435454
rect 361250 434898 361486 435134
rect 371490 435218 371726 435454
rect 371490 434898 371726 435134
rect 381730 435218 381966 435454
rect 381730 434898 381966 435134
rect 391970 435218 392206 435454
rect 391970 434898 392206 435134
rect 402210 435218 402446 435454
rect 402210 434898 402446 435134
rect 412450 435218 412686 435454
rect 412450 434898 412686 435134
rect 422690 435218 422926 435454
rect 422690 434898 422926 435134
rect 432930 435218 433166 435454
rect 432930 434898 433166 435134
rect 443170 435218 443406 435454
rect 443170 434898 443406 435134
rect 453410 435218 453646 435454
rect 453410 434898 453646 435134
rect 463650 435218 463886 435454
rect 463650 434898 463886 435134
rect 473890 435218 474126 435454
rect 473890 434898 474126 435134
rect 484130 435218 484366 435454
rect 484130 434898 484366 435134
rect 494370 435218 494606 435454
rect 494370 434898 494606 435134
rect 504610 435218 504846 435454
rect 504610 434898 504846 435134
rect 514850 435218 515086 435454
rect 514850 434898 515086 435134
rect 525090 435218 525326 435454
rect 525090 434898 525326 435134
rect 535330 435218 535566 435454
rect 535330 434898 535566 435134
rect 28450 417218 28686 417454
rect 28450 416898 28686 417134
rect 38690 417218 38926 417454
rect 38690 416898 38926 417134
rect 48930 417218 49166 417454
rect 48930 416898 49166 417134
rect 59170 417218 59406 417454
rect 59170 416898 59406 417134
rect 69410 417218 69646 417454
rect 69410 416898 69646 417134
rect 79650 417218 79886 417454
rect 79650 416898 79886 417134
rect 89890 417218 90126 417454
rect 89890 416898 90126 417134
rect 100130 417218 100366 417454
rect 100130 416898 100366 417134
rect 110370 417218 110606 417454
rect 110370 416898 110606 417134
rect 120610 417218 120846 417454
rect 120610 416898 120846 417134
rect 130850 417218 131086 417454
rect 130850 416898 131086 417134
rect 141090 417218 141326 417454
rect 141090 416898 141326 417134
rect 151330 417218 151566 417454
rect 151330 416898 151566 417134
rect 161570 417218 161806 417454
rect 161570 416898 161806 417134
rect 171810 417218 172046 417454
rect 171810 416898 172046 417134
rect 182050 417218 182286 417454
rect 182050 416898 182286 417134
rect 192290 417218 192526 417454
rect 192290 416898 192526 417134
rect 202530 417218 202766 417454
rect 202530 416898 202766 417134
rect 212770 417218 213006 417454
rect 212770 416898 213006 417134
rect 223010 417218 223246 417454
rect 223010 416898 223246 417134
rect 233250 417218 233486 417454
rect 233250 416898 233486 417134
rect 243490 417218 243726 417454
rect 243490 416898 243726 417134
rect 253730 417218 253966 417454
rect 253730 416898 253966 417134
rect 263970 417218 264206 417454
rect 263970 416898 264206 417134
rect 274210 417218 274446 417454
rect 274210 416898 274446 417134
rect 284450 417218 284686 417454
rect 284450 416898 284686 417134
rect 294690 417218 294926 417454
rect 294690 416898 294926 417134
rect 304930 417218 305166 417454
rect 304930 416898 305166 417134
rect 315170 417218 315406 417454
rect 315170 416898 315406 417134
rect 325410 417218 325646 417454
rect 325410 416898 325646 417134
rect 335650 417218 335886 417454
rect 335650 416898 335886 417134
rect 345890 417218 346126 417454
rect 345890 416898 346126 417134
rect 356130 417218 356366 417454
rect 356130 416898 356366 417134
rect 366370 417218 366606 417454
rect 366370 416898 366606 417134
rect 376610 417218 376846 417454
rect 376610 416898 376846 417134
rect 386850 417218 387086 417454
rect 386850 416898 387086 417134
rect 397090 417218 397326 417454
rect 397090 416898 397326 417134
rect 407330 417218 407566 417454
rect 407330 416898 407566 417134
rect 417570 417218 417806 417454
rect 417570 416898 417806 417134
rect 427810 417218 428046 417454
rect 427810 416898 428046 417134
rect 438050 417218 438286 417454
rect 438050 416898 438286 417134
rect 448290 417218 448526 417454
rect 448290 416898 448526 417134
rect 458530 417218 458766 417454
rect 458530 416898 458766 417134
rect 468770 417218 469006 417454
rect 468770 416898 469006 417134
rect 479010 417218 479246 417454
rect 479010 416898 479246 417134
rect 489250 417218 489486 417454
rect 489250 416898 489486 417134
rect 499490 417218 499726 417454
rect 499490 416898 499726 417134
rect 509730 417218 509966 417454
rect 509730 416898 509966 417134
rect 519970 417218 520206 417454
rect 519970 416898 520206 417134
rect 530210 417218 530446 417454
rect 530210 416898 530446 417134
rect 15786 402938 16022 403174
rect 16106 402938 16342 403174
rect 15786 402618 16022 402854
rect 16106 402618 16342 402854
rect 541746 406658 541982 406894
rect 542066 406658 542302 406894
rect 541746 406338 541982 406574
rect 542066 406338 542302 406574
rect 23330 399218 23566 399454
rect 23330 398898 23566 399134
rect 33570 399218 33806 399454
rect 33570 398898 33806 399134
rect 43810 399218 44046 399454
rect 43810 398898 44046 399134
rect 54050 399218 54286 399454
rect 54050 398898 54286 399134
rect 64290 399218 64526 399454
rect 64290 398898 64526 399134
rect 74530 399218 74766 399454
rect 74530 398898 74766 399134
rect 84770 399218 85006 399454
rect 84770 398898 85006 399134
rect 95010 399218 95246 399454
rect 95010 398898 95246 399134
rect 105250 399218 105486 399454
rect 105250 398898 105486 399134
rect 115490 399218 115726 399454
rect 115490 398898 115726 399134
rect 125730 399218 125966 399454
rect 125730 398898 125966 399134
rect 135970 399218 136206 399454
rect 135970 398898 136206 399134
rect 146210 399218 146446 399454
rect 146210 398898 146446 399134
rect 156450 399218 156686 399454
rect 156450 398898 156686 399134
rect 166690 399218 166926 399454
rect 166690 398898 166926 399134
rect 176930 399218 177166 399454
rect 176930 398898 177166 399134
rect 187170 399218 187406 399454
rect 187170 398898 187406 399134
rect 197410 399218 197646 399454
rect 197410 398898 197646 399134
rect 207650 399218 207886 399454
rect 207650 398898 207886 399134
rect 217890 399218 218126 399454
rect 217890 398898 218126 399134
rect 228130 399218 228366 399454
rect 228130 398898 228366 399134
rect 238370 399218 238606 399454
rect 238370 398898 238606 399134
rect 248610 399218 248846 399454
rect 248610 398898 248846 399134
rect 258850 399218 259086 399454
rect 258850 398898 259086 399134
rect 269090 399218 269326 399454
rect 269090 398898 269326 399134
rect 279330 399218 279566 399454
rect 279330 398898 279566 399134
rect 289570 399218 289806 399454
rect 289570 398898 289806 399134
rect 299810 399218 300046 399454
rect 299810 398898 300046 399134
rect 310050 399218 310286 399454
rect 310050 398898 310286 399134
rect 320290 399218 320526 399454
rect 320290 398898 320526 399134
rect 330530 399218 330766 399454
rect 330530 398898 330766 399134
rect 340770 399218 341006 399454
rect 340770 398898 341006 399134
rect 351010 399218 351246 399454
rect 351010 398898 351246 399134
rect 361250 399218 361486 399454
rect 361250 398898 361486 399134
rect 371490 399218 371726 399454
rect 371490 398898 371726 399134
rect 381730 399218 381966 399454
rect 381730 398898 381966 399134
rect 391970 399218 392206 399454
rect 391970 398898 392206 399134
rect 402210 399218 402446 399454
rect 402210 398898 402446 399134
rect 412450 399218 412686 399454
rect 412450 398898 412686 399134
rect 422690 399218 422926 399454
rect 422690 398898 422926 399134
rect 432930 399218 433166 399454
rect 432930 398898 433166 399134
rect 443170 399218 443406 399454
rect 443170 398898 443406 399134
rect 453410 399218 453646 399454
rect 453410 398898 453646 399134
rect 463650 399218 463886 399454
rect 463650 398898 463886 399134
rect 473890 399218 474126 399454
rect 473890 398898 474126 399134
rect 484130 399218 484366 399454
rect 484130 398898 484366 399134
rect 494370 399218 494606 399454
rect 494370 398898 494606 399134
rect 504610 399218 504846 399454
rect 504610 398898 504846 399134
rect 514850 399218 515086 399454
rect 514850 398898 515086 399134
rect 525090 399218 525326 399454
rect 525090 398898 525326 399134
rect 535330 399218 535566 399454
rect 535330 398898 535566 399134
rect 28450 381218 28686 381454
rect 28450 380898 28686 381134
rect 38690 381218 38926 381454
rect 38690 380898 38926 381134
rect 48930 381218 49166 381454
rect 48930 380898 49166 381134
rect 59170 381218 59406 381454
rect 59170 380898 59406 381134
rect 69410 381218 69646 381454
rect 69410 380898 69646 381134
rect 79650 381218 79886 381454
rect 79650 380898 79886 381134
rect 89890 381218 90126 381454
rect 89890 380898 90126 381134
rect 100130 381218 100366 381454
rect 100130 380898 100366 381134
rect 110370 381218 110606 381454
rect 110370 380898 110606 381134
rect 120610 381218 120846 381454
rect 120610 380898 120846 381134
rect 130850 381218 131086 381454
rect 130850 380898 131086 381134
rect 141090 381218 141326 381454
rect 141090 380898 141326 381134
rect 151330 381218 151566 381454
rect 151330 380898 151566 381134
rect 161570 381218 161806 381454
rect 161570 380898 161806 381134
rect 171810 381218 172046 381454
rect 171810 380898 172046 381134
rect 182050 381218 182286 381454
rect 182050 380898 182286 381134
rect 192290 381218 192526 381454
rect 192290 380898 192526 381134
rect 202530 381218 202766 381454
rect 202530 380898 202766 381134
rect 212770 381218 213006 381454
rect 212770 380898 213006 381134
rect 223010 381218 223246 381454
rect 223010 380898 223246 381134
rect 233250 381218 233486 381454
rect 233250 380898 233486 381134
rect 243490 381218 243726 381454
rect 243490 380898 243726 381134
rect 253730 381218 253966 381454
rect 253730 380898 253966 381134
rect 263970 381218 264206 381454
rect 263970 380898 264206 381134
rect 274210 381218 274446 381454
rect 274210 380898 274446 381134
rect 284450 381218 284686 381454
rect 284450 380898 284686 381134
rect 294690 381218 294926 381454
rect 294690 380898 294926 381134
rect 304930 381218 305166 381454
rect 304930 380898 305166 381134
rect 315170 381218 315406 381454
rect 315170 380898 315406 381134
rect 325410 381218 325646 381454
rect 325410 380898 325646 381134
rect 335650 381218 335886 381454
rect 335650 380898 335886 381134
rect 345890 381218 346126 381454
rect 345890 380898 346126 381134
rect 356130 381218 356366 381454
rect 356130 380898 356366 381134
rect 366370 381218 366606 381454
rect 366370 380898 366606 381134
rect 376610 381218 376846 381454
rect 376610 380898 376846 381134
rect 386850 381218 387086 381454
rect 386850 380898 387086 381134
rect 397090 381218 397326 381454
rect 397090 380898 397326 381134
rect 407330 381218 407566 381454
rect 407330 380898 407566 381134
rect 417570 381218 417806 381454
rect 417570 380898 417806 381134
rect 427810 381218 428046 381454
rect 427810 380898 428046 381134
rect 438050 381218 438286 381454
rect 438050 380898 438286 381134
rect 448290 381218 448526 381454
rect 448290 380898 448526 381134
rect 458530 381218 458766 381454
rect 458530 380898 458766 381134
rect 468770 381218 469006 381454
rect 468770 380898 469006 381134
rect 479010 381218 479246 381454
rect 479010 380898 479246 381134
rect 489250 381218 489486 381454
rect 489250 380898 489486 381134
rect 499490 381218 499726 381454
rect 499490 380898 499726 381134
rect 509730 381218 509966 381454
rect 509730 380898 509966 381134
rect 519970 381218 520206 381454
rect 519970 380898 520206 381134
rect 530210 381218 530446 381454
rect 530210 380898 530446 381134
rect 15786 366938 16022 367174
rect 16106 366938 16342 367174
rect 15786 366618 16022 366854
rect 16106 366618 16342 366854
rect 541746 370658 541982 370894
rect 542066 370658 542302 370894
rect 541746 370338 541982 370574
rect 542066 370338 542302 370574
rect 23330 363218 23566 363454
rect 23330 362898 23566 363134
rect 33570 363218 33806 363454
rect 33570 362898 33806 363134
rect 43810 363218 44046 363454
rect 43810 362898 44046 363134
rect 54050 363218 54286 363454
rect 54050 362898 54286 363134
rect 64290 363218 64526 363454
rect 64290 362898 64526 363134
rect 74530 363218 74766 363454
rect 74530 362898 74766 363134
rect 84770 363218 85006 363454
rect 84770 362898 85006 363134
rect 95010 363218 95246 363454
rect 95010 362898 95246 363134
rect 105250 363218 105486 363454
rect 105250 362898 105486 363134
rect 115490 363218 115726 363454
rect 115490 362898 115726 363134
rect 125730 363218 125966 363454
rect 125730 362898 125966 363134
rect 135970 363218 136206 363454
rect 135970 362898 136206 363134
rect 146210 363218 146446 363454
rect 146210 362898 146446 363134
rect 156450 363218 156686 363454
rect 156450 362898 156686 363134
rect 166690 363218 166926 363454
rect 166690 362898 166926 363134
rect 176930 363218 177166 363454
rect 176930 362898 177166 363134
rect 187170 363218 187406 363454
rect 187170 362898 187406 363134
rect 197410 363218 197646 363454
rect 197410 362898 197646 363134
rect 207650 363218 207886 363454
rect 207650 362898 207886 363134
rect 217890 363218 218126 363454
rect 217890 362898 218126 363134
rect 228130 363218 228366 363454
rect 228130 362898 228366 363134
rect 238370 363218 238606 363454
rect 238370 362898 238606 363134
rect 248610 363218 248846 363454
rect 248610 362898 248846 363134
rect 258850 363218 259086 363454
rect 258850 362898 259086 363134
rect 269090 363218 269326 363454
rect 269090 362898 269326 363134
rect 279330 363218 279566 363454
rect 279330 362898 279566 363134
rect 289570 363218 289806 363454
rect 289570 362898 289806 363134
rect 299810 363218 300046 363454
rect 299810 362898 300046 363134
rect 310050 363218 310286 363454
rect 310050 362898 310286 363134
rect 320290 363218 320526 363454
rect 320290 362898 320526 363134
rect 330530 363218 330766 363454
rect 330530 362898 330766 363134
rect 340770 363218 341006 363454
rect 340770 362898 341006 363134
rect 351010 363218 351246 363454
rect 351010 362898 351246 363134
rect 361250 363218 361486 363454
rect 361250 362898 361486 363134
rect 371490 363218 371726 363454
rect 371490 362898 371726 363134
rect 381730 363218 381966 363454
rect 381730 362898 381966 363134
rect 391970 363218 392206 363454
rect 391970 362898 392206 363134
rect 402210 363218 402446 363454
rect 402210 362898 402446 363134
rect 412450 363218 412686 363454
rect 412450 362898 412686 363134
rect 422690 363218 422926 363454
rect 422690 362898 422926 363134
rect 432930 363218 433166 363454
rect 432930 362898 433166 363134
rect 443170 363218 443406 363454
rect 443170 362898 443406 363134
rect 453410 363218 453646 363454
rect 453410 362898 453646 363134
rect 463650 363218 463886 363454
rect 463650 362898 463886 363134
rect 473890 363218 474126 363454
rect 473890 362898 474126 363134
rect 484130 363218 484366 363454
rect 484130 362898 484366 363134
rect 494370 363218 494606 363454
rect 494370 362898 494606 363134
rect 504610 363218 504846 363454
rect 504610 362898 504846 363134
rect 514850 363218 515086 363454
rect 514850 362898 515086 363134
rect 525090 363218 525326 363454
rect 525090 362898 525326 363134
rect 535330 363218 535566 363454
rect 535330 362898 535566 363134
rect 28450 345218 28686 345454
rect 28450 344898 28686 345134
rect 38690 345218 38926 345454
rect 38690 344898 38926 345134
rect 48930 345218 49166 345454
rect 48930 344898 49166 345134
rect 59170 345218 59406 345454
rect 59170 344898 59406 345134
rect 69410 345218 69646 345454
rect 69410 344898 69646 345134
rect 79650 345218 79886 345454
rect 79650 344898 79886 345134
rect 89890 345218 90126 345454
rect 89890 344898 90126 345134
rect 100130 345218 100366 345454
rect 100130 344898 100366 345134
rect 110370 345218 110606 345454
rect 110370 344898 110606 345134
rect 120610 345218 120846 345454
rect 120610 344898 120846 345134
rect 130850 345218 131086 345454
rect 130850 344898 131086 345134
rect 141090 345218 141326 345454
rect 141090 344898 141326 345134
rect 151330 345218 151566 345454
rect 151330 344898 151566 345134
rect 161570 345218 161806 345454
rect 161570 344898 161806 345134
rect 171810 345218 172046 345454
rect 171810 344898 172046 345134
rect 182050 345218 182286 345454
rect 182050 344898 182286 345134
rect 192290 345218 192526 345454
rect 192290 344898 192526 345134
rect 202530 345218 202766 345454
rect 202530 344898 202766 345134
rect 212770 345218 213006 345454
rect 212770 344898 213006 345134
rect 223010 345218 223246 345454
rect 223010 344898 223246 345134
rect 233250 345218 233486 345454
rect 233250 344898 233486 345134
rect 243490 345218 243726 345454
rect 243490 344898 243726 345134
rect 253730 345218 253966 345454
rect 253730 344898 253966 345134
rect 263970 345218 264206 345454
rect 263970 344898 264206 345134
rect 274210 345218 274446 345454
rect 274210 344898 274446 345134
rect 284450 345218 284686 345454
rect 284450 344898 284686 345134
rect 294690 345218 294926 345454
rect 294690 344898 294926 345134
rect 304930 345218 305166 345454
rect 304930 344898 305166 345134
rect 315170 345218 315406 345454
rect 315170 344898 315406 345134
rect 325410 345218 325646 345454
rect 325410 344898 325646 345134
rect 335650 345218 335886 345454
rect 335650 344898 335886 345134
rect 345890 345218 346126 345454
rect 345890 344898 346126 345134
rect 356130 345218 356366 345454
rect 356130 344898 356366 345134
rect 366370 345218 366606 345454
rect 366370 344898 366606 345134
rect 376610 345218 376846 345454
rect 376610 344898 376846 345134
rect 386850 345218 387086 345454
rect 386850 344898 387086 345134
rect 397090 345218 397326 345454
rect 397090 344898 397326 345134
rect 407330 345218 407566 345454
rect 407330 344898 407566 345134
rect 417570 345218 417806 345454
rect 417570 344898 417806 345134
rect 427810 345218 428046 345454
rect 427810 344898 428046 345134
rect 438050 345218 438286 345454
rect 438050 344898 438286 345134
rect 448290 345218 448526 345454
rect 448290 344898 448526 345134
rect 458530 345218 458766 345454
rect 458530 344898 458766 345134
rect 468770 345218 469006 345454
rect 468770 344898 469006 345134
rect 479010 345218 479246 345454
rect 479010 344898 479246 345134
rect 489250 345218 489486 345454
rect 489250 344898 489486 345134
rect 499490 345218 499726 345454
rect 499490 344898 499726 345134
rect 509730 345218 509966 345454
rect 509730 344898 509966 345134
rect 519970 345218 520206 345454
rect 519970 344898 520206 345134
rect 530210 345218 530446 345454
rect 530210 344898 530446 345134
rect 15786 330938 16022 331174
rect 16106 330938 16342 331174
rect 15786 330618 16022 330854
rect 16106 330618 16342 330854
rect 541746 334658 541982 334894
rect 542066 334658 542302 334894
rect 541746 334338 541982 334574
rect 542066 334338 542302 334574
rect 23330 327218 23566 327454
rect 23330 326898 23566 327134
rect 33570 327218 33806 327454
rect 33570 326898 33806 327134
rect 43810 327218 44046 327454
rect 43810 326898 44046 327134
rect 54050 327218 54286 327454
rect 54050 326898 54286 327134
rect 64290 327218 64526 327454
rect 64290 326898 64526 327134
rect 74530 327218 74766 327454
rect 74530 326898 74766 327134
rect 84770 327218 85006 327454
rect 84770 326898 85006 327134
rect 95010 327218 95246 327454
rect 95010 326898 95246 327134
rect 105250 327218 105486 327454
rect 105250 326898 105486 327134
rect 115490 327218 115726 327454
rect 115490 326898 115726 327134
rect 125730 327218 125966 327454
rect 125730 326898 125966 327134
rect 135970 327218 136206 327454
rect 135970 326898 136206 327134
rect 146210 327218 146446 327454
rect 146210 326898 146446 327134
rect 156450 327218 156686 327454
rect 156450 326898 156686 327134
rect 166690 327218 166926 327454
rect 166690 326898 166926 327134
rect 176930 327218 177166 327454
rect 176930 326898 177166 327134
rect 187170 327218 187406 327454
rect 187170 326898 187406 327134
rect 197410 327218 197646 327454
rect 197410 326898 197646 327134
rect 207650 327218 207886 327454
rect 207650 326898 207886 327134
rect 217890 327218 218126 327454
rect 217890 326898 218126 327134
rect 228130 327218 228366 327454
rect 228130 326898 228366 327134
rect 238370 327218 238606 327454
rect 238370 326898 238606 327134
rect 248610 327218 248846 327454
rect 248610 326898 248846 327134
rect 258850 327218 259086 327454
rect 258850 326898 259086 327134
rect 269090 327218 269326 327454
rect 269090 326898 269326 327134
rect 279330 327218 279566 327454
rect 279330 326898 279566 327134
rect 289570 327218 289806 327454
rect 289570 326898 289806 327134
rect 299810 327218 300046 327454
rect 299810 326898 300046 327134
rect 310050 327218 310286 327454
rect 310050 326898 310286 327134
rect 320290 327218 320526 327454
rect 320290 326898 320526 327134
rect 330530 327218 330766 327454
rect 330530 326898 330766 327134
rect 340770 327218 341006 327454
rect 340770 326898 341006 327134
rect 351010 327218 351246 327454
rect 351010 326898 351246 327134
rect 361250 327218 361486 327454
rect 361250 326898 361486 327134
rect 371490 327218 371726 327454
rect 371490 326898 371726 327134
rect 381730 327218 381966 327454
rect 381730 326898 381966 327134
rect 391970 327218 392206 327454
rect 391970 326898 392206 327134
rect 402210 327218 402446 327454
rect 402210 326898 402446 327134
rect 412450 327218 412686 327454
rect 412450 326898 412686 327134
rect 422690 327218 422926 327454
rect 422690 326898 422926 327134
rect 432930 327218 433166 327454
rect 432930 326898 433166 327134
rect 443170 327218 443406 327454
rect 443170 326898 443406 327134
rect 453410 327218 453646 327454
rect 453410 326898 453646 327134
rect 463650 327218 463886 327454
rect 463650 326898 463886 327134
rect 473890 327218 474126 327454
rect 473890 326898 474126 327134
rect 484130 327218 484366 327454
rect 484130 326898 484366 327134
rect 494370 327218 494606 327454
rect 494370 326898 494606 327134
rect 504610 327218 504846 327454
rect 504610 326898 504846 327134
rect 514850 327218 515086 327454
rect 514850 326898 515086 327134
rect 525090 327218 525326 327454
rect 525090 326898 525326 327134
rect 535330 327218 535566 327454
rect 535330 326898 535566 327134
rect 28450 309218 28686 309454
rect 28450 308898 28686 309134
rect 38690 309218 38926 309454
rect 38690 308898 38926 309134
rect 48930 309218 49166 309454
rect 48930 308898 49166 309134
rect 59170 309218 59406 309454
rect 59170 308898 59406 309134
rect 69410 309218 69646 309454
rect 69410 308898 69646 309134
rect 79650 309218 79886 309454
rect 79650 308898 79886 309134
rect 89890 309218 90126 309454
rect 89890 308898 90126 309134
rect 100130 309218 100366 309454
rect 100130 308898 100366 309134
rect 110370 309218 110606 309454
rect 110370 308898 110606 309134
rect 120610 309218 120846 309454
rect 120610 308898 120846 309134
rect 130850 309218 131086 309454
rect 130850 308898 131086 309134
rect 141090 309218 141326 309454
rect 141090 308898 141326 309134
rect 151330 309218 151566 309454
rect 151330 308898 151566 309134
rect 161570 309218 161806 309454
rect 161570 308898 161806 309134
rect 171810 309218 172046 309454
rect 171810 308898 172046 309134
rect 182050 309218 182286 309454
rect 182050 308898 182286 309134
rect 192290 309218 192526 309454
rect 192290 308898 192526 309134
rect 202530 309218 202766 309454
rect 202530 308898 202766 309134
rect 212770 309218 213006 309454
rect 212770 308898 213006 309134
rect 223010 309218 223246 309454
rect 223010 308898 223246 309134
rect 233250 309218 233486 309454
rect 233250 308898 233486 309134
rect 243490 309218 243726 309454
rect 243490 308898 243726 309134
rect 253730 309218 253966 309454
rect 253730 308898 253966 309134
rect 263970 309218 264206 309454
rect 263970 308898 264206 309134
rect 274210 309218 274446 309454
rect 274210 308898 274446 309134
rect 284450 309218 284686 309454
rect 284450 308898 284686 309134
rect 294690 309218 294926 309454
rect 294690 308898 294926 309134
rect 304930 309218 305166 309454
rect 304930 308898 305166 309134
rect 315170 309218 315406 309454
rect 315170 308898 315406 309134
rect 325410 309218 325646 309454
rect 325410 308898 325646 309134
rect 335650 309218 335886 309454
rect 335650 308898 335886 309134
rect 345890 309218 346126 309454
rect 345890 308898 346126 309134
rect 356130 309218 356366 309454
rect 356130 308898 356366 309134
rect 366370 309218 366606 309454
rect 366370 308898 366606 309134
rect 376610 309218 376846 309454
rect 376610 308898 376846 309134
rect 386850 309218 387086 309454
rect 386850 308898 387086 309134
rect 397090 309218 397326 309454
rect 397090 308898 397326 309134
rect 407330 309218 407566 309454
rect 407330 308898 407566 309134
rect 417570 309218 417806 309454
rect 417570 308898 417806 309134
rect 427810 309218 428046 309454
rect 427810 308898 428046 309134
rect 438050 309218 438286 309454
rect 438050 308898 438286 309134
rect 448290 309218 448526 309454
rect 448290 308898 448526 309134
rect 458530 309218 458766 309454
rect 458530 308898 458766 309134
rect 468770 309218 469006 309454
rect 468770 308898 469006 309134
rect 479010 309218 479246 309454
rect 479010 308898 479246 309134
rect 489250 309218 489486 309454
rect 489250 308898 489486 309134
rect 499490 309218 499726 309454
rect 499490 308898 499726 309134
rect 509730 309218 509966 309454
rect 509730 308898 509966 309134
rect 519970 309218 520206 309454
rect 519970 308898 520206 309134
rect 530210 309218 530446 309454
rect 530210 308898 530446 309134
rect 15786 294938 16022 295174
rect 16106 294938 16342 295174
rect 15786 294618 16022 294854
rect 16106 294618 16342 294854
rect 541746 298658 541982 298894
rect 542066 298658 542302 298894
rect 541746 298338 541982 298574
rect 542066 298338 542302 298574
rect 23330 291218 23566 291454
rect 23330 290898 23566 291134
rect 33570 291218 33806 291454
rect 33570 290898 33806 291134
rect 43810 291218 44046 291454
rect 43810 290898 44046 291134
rect 54050 291218 54286 291454
rect 54050 290898 54286 291134
rect 64290 291218 64526 291454
rect 64290 290898 64526 291134
rect 74530 291218 74766 291454
rect 74530 290898 74766 291134
rect 84770 291218 85006 291454
rect 84770 290898 85006 291134
rect 95010 291218 95246 291454
rect 95010 290898 95246 291134
rect 105250 291218 105486 291454
rect 105250 290898 105486 291134
rect 115490 291218 115726 291454
rect 115490 290898 115726 291134
rect 125730 291218 125966 291454
rect 125730 290898 125966 291134
rect 135970 291218 136206 291454
rect 135970 290898 136206 291134
rect 146210 291218 146446 291454
rect 146210 290898 146446 291134
rect 156450 291218 156686 291454
rect 156450 290898 156686 291134
rect 166690 291218 166926 291454
rect 166690 290898 166926 291134
rect 176930 291218 177166 291454
rect 176930 290898 177166 291134
rect 187170 291218 187406 291454
rect 187170 290898 187406 291134
rect 197410 291218 197646 291454
rect 197410 290898 197646 291134
rect 207650 291218 207886 291454
rect 207650 290898 207886 291134
rect 217890 291218 218126 291454
rect 217890 290898 218126 291134
rect 228130 291218 228366 291454
rect 228130 290898 228366 291134
rect 238370 291218 238606 291454
rect 238370 290898 238606 291134
rect 248610 291218 248846 291454
rect 248610 290898 248846 291134
rect 258850 291218 259086 291454
rect 258850 290898 259086 291134
rect 269090 291218 269326 291454
rect 269090 290898 269326 291134
rect 279330 291218 279566 291454
rect 279330 290898 279566 291134
rect 289570 291218 289806 291454
rect 289570 290898 289806 291134
rect 299810 291218 300046 291454
rect 299810 290898 300046 291134
rect 310050 291218 310286 291454
rect 310050 290898 310286 291134
rect 320290 291218 320526 291454
rect 320290 290898 320526 291134
rect 330530 291218 330766 291454
rect 330530 290898 330766 291134
rect 340770 291218 341006 291454
rect 340770 290898 341006 291134
rect 351010 291218 351246 291454
rect 351010 290898 351246 291134
rect 361250 291218 361486 291454
rect 361250 290898 361486 291134
rect 371490 291218 371726 291454
rect 371490 290898 371726 291134
rect 381730 291218 381966 291454
rect 381730 290898 381966 291134
rect 391970 291218 392206 291454
rect 391970 290898 392206 291134
rect 402210 291218 402446 291454
rect 402210 290898 402446 291134
rect 412450 291218 412686 291454
rect 412450 290898 412686 291134
rect 422690 291218 422926 291454
rect 422690 290898 422926 291134
rect 432930 291218 433166 291454
rect 432930 290898 433166 291134
rect 443170 291218 443406 291454
rect 443170 290898 443406 291134
rect 453410 291218 453646 291454
rect 453410 290898 453646 291134
rect 463650 291218 463886 291454
rect 463650 290898 463886 291134
rect 473890 291218 474126 291454
rect 473890 290898 474126 291134
rect 484130 291218 484366 291454
rect 484130 290898 484366 291134
rect 494370 291218 494606 291454
rect 494370 290898 494606 291134
rect 504610 291218 504846 291454
rect 504610 290898 504846 291134
rect 514850 291218 515086 291454
rect 514850 290898 515086 291134
rect 525090 291218 525326 291454
rect 525090 290898 525326 291134
rect 535330 291218 535566 291454
rect 535330 290898 535566 291134
rect 28450 273218 28686 273454
rect 28450 272898 28686 273134
rect 38690 273218 38926 273454
rect 38690 272898 38926 273134
rect 48930 273218 49166 273454
rect 48930 272898 49166 273134
rect 59170 273218 59406 273454
rect 59170 272898 59406 273134
rect 69410 273218 69646 273454
rect 69410 272898 69646 273134
rect 79650 273218 79886 273454
rect 79650 272898 79886 273134
rect 89890 273218 90126 273454
rect 89890 272898 90126 273134
rect 100130 273218 100366 273454
rect 100130 272898 100366 273134
rect 110370 273218 110606 273454
rect 110370 272898 110606 273134
rect 120610 273218 120846 273454
rect 120610 272898 120846 273134
rect 130850 273218 131086 273454
rect 130850 272898 131086 273134
rect 141090 273218 141326 273454
rect 141090 272898 141326 273134
rect 151330 273218 151566 273454
rect 151330 272898 151566 273134
rect 161570 273218 161806 273454
rect 161570 272898 161806 273134
rect 171810 273218 172046 273454
rect 171810 272898 172046 273134
rect 182050 273218 182286 273454
rect 182050 272898 182286 273134
rect 192290 273218 192526 273454
rect 192290 272898 192526 273134
rect 202530 273218 202766 273454
rect 202530 272898 202766 273134
rect 212770 273218 213006 273454
rect 212770 272898 213006 273134
rect 223010 273218 223246 273454
rect 223010 272898 223246 273134
rect 233250 273218 233486 273454
rect 233250 272898 233486 273134
rect 243490 273218 243726 273454
rect 243490 272898 243726 273134
rect 253730 273218 253966 273454
rect 253730 272898 253966 273134
rect 263970 273218 264206 273454
rect 263970 272898 264206 273134
rect 274210 273218 274446 273454
rect 274210 272898 274446 273134
rect 284450 273218 284686 273454
rect 284450 272898 284686 273134
rect 294690 273218 294926 273454
rect 294690 272898 294926 273134
rect 304930 273218 305166 273454
rect 304930 272898 305166 273134
rect 315170 273218 315406 273454
rect 315170 272898 315406 273134
rect 325410 273218 325646 273454
rect 325410 272898 325646 273134
rect 335650 273218 335886 273454
rect 335650 272898 335886 273134
rect 345890 273218 346126 273454
rect 345890 272898 346126 273134
rect 356130 273218 356366 273454
rect 356130 272898 356366 273134
rect 366370 273218 366606 273454
rect 366370 272898 366606 273134
rect 376610 273218 376846 273454
rect 376610 272898 376846 273134
rect 386850 273218 387086 273454
rect 386850 272898 387086 273134
rect 397090 273218 397326 273454
rect 397090 272898 397326 273134
rect 407330 273218 407566 273454
rect 407330 272898 407566 273134
rect 417570 273218 417806 273454
rect 417570 272898 417806 273134
rect 427810 273218 428046 273454
rect 427810 272898 428046 273134
rect 438050 273218 438286 273454
rect 438050 272898 438286 273134
rect 448290 273218 448526 273454
rect 448290 272898 448526 273134
rect 458530 273218 458766 273454
rect 458530 272898 458766 273134
rect 468770 273218 469006 273454
rect 468770 272898 469006 273134
rect 479010 273218 479246 273454
rect 479010 272898 479246 273134
rect 489250 273218 489486 273454
rect 489250 272898 489486 273134
rect 499490 273218 499726 273454
rect 499490 272898 499726 273134
rect 509730 273218 509966 273454
rect 509730 272898 509966 273134
rect 519970 273218 520206 273454
rect 519970 272898 520206 273134
rect 530210 273218 530446 273454
rect 530210 272898 530446 273134
rect 15786 258938 16022 259174
rect 16106 258938 16342 259174
rect 15786 258618 16022 258854
rect 16106 258618 16342 258854
rect 541746 262658 541982 262894
rect 542066 262658 542302 262894
rect 541746 262338 541982 262574
rect 542066 262338 542302 262574
rect 23330 255218 23566 255454
rect 23330 254898 23566 255134
rect 33570 255218 33806 255454
rect 33570 254898 33806 255134
rect 43810 255218 44046 255454
rect 43810 254898 44046 255134
rect 54050 255218 54286 255454
rect 54050 254898 54286 255134
rect 64290 255218 64526 255454
rect 64290 254898 64526 255134
rect 74530 255218 74766 255454
rect 74530 254898 74766 255134
rect 84770 255218 85006 255454
rect 84770 254898 85006 255134
rect 95010 255218 95246 255454
rect 95010 254898 95246 255134
rect 105250 255218 105486 255454
rect 105250 254898 105486 255134
rect 115490 255218 115726 255454
rect 115490 254898 115726 255134
rect 125730 255218 125966 255454
rect 125730 254898 125966 255134
rect 135970 255218 136206 255454
rect 135970 254898 136206 255134
rect 146210 255218 146446 255454
rect 146210 254898 146446 255134
rect 156450 255218 156686 255454
rect 156450 254898 156686 255134
rect 166690 255218 166926 255454
rect 166690 254898 166926 255134
rect 176930 255218 177166 255454
rect 176930 254898 177166 255134
rect 187170 255218 187406 255454
rect 187170 254898 187406 255134
rect 197410 255218 197646 255454
rect 197410 254898 197646 255134
rect 207650 255218 207886 255454
rect 207650 254898 207886 255134
rect 217890 255218 218126 255454
rect 217890 254898 218126 255134
rect 228130 255218 228366 255454
rect 228130 254898 228366 255134
rect 238370 255218 238606 255454
rect 238370 254898 238606 255134
rect 248610 255218 248846 255454
rect 248610 254898 248846 255134
rect 258850 255218 259086 255454
rect 258850 254898 259086 255134
rect 269090 255218 269326 255454
rect 269090 254898 269326 255134
rect 279330 255218 279566 255454
rect 279330 254898 279566 255134
rect 289570 255218 289806 255454
rect 289570 254898 289806 255134
rect 299810 255218 300046 255454
rect 299810 254898 300046 255134
rect 310050 255218 310286 255454
rect 310050 254898 310286 255134
rect 320290 255218 320526 255454
rect 320290 254898 320526 255134
rect 330530 255218 330766 255454
rect 330530 254898 330766 255134
rect 340770 255218 341006 255454
rect 340770 254898 341006 255134
rect 351010 255218 351246 255454
rect 351010 254898 351246 255134
rect 361250 255218 361486 255454
rect 361250 254898 361486 255134
rect 371490 255218 371726 255454
rect 371490 254898 371726 255134
rect 381730 255218 381966 255454
rect 381730 254898 381966 255134
rect 391970 255218 392206 255454
rect 391970 254898 392206 255134
rect 402210 255218 402446 255454
rect 402210 254898 402446 255134
rect 412450 255218 412686 255454
rect 412450 254898 412686 255134
rect 422690 255218 422926 255454
rect 422690 254898 422926 255134
rect 432930 255218 433166 255454
rect 432930 254898 433166 255134
rect 443170 255218 443406 255454
rect 443170 254898 443406 255134
rect 453410 255218 453646 255454
rect 453410 254898 453646 255134
rect 463650 255218 463886 255454
rect 463650 254898 463886 255134
rect 473890 255218 474126 255454
rect 473890 254898 474126 255134
rect 484130 255218 484366 255454
rect 484130 254898 484366 255134
rect 494370 255218 494606 255454
rect 494370 254898 494606 255134
rect 504610 255218 504846 255454
rect 504610 254898 504846 255134
rect 514850 255218 515086 255454
rect 514850 254898 515086 255134
rect 525090 255218 525326 255454
rect 525090 254898 525326 255134
rect 535330 255218 535566 255454
rect 535330 254898 535566 255134
rect 28450 237218 28686 237454
rect 28450 236898 28686 237134
rect 38690 237218 38926 237454
rect 38690 236898 38926 237134
rect 48930 237218 49166 237454
rect 48930 236898 49166 237134
rect 59170 237218 59406 237454
rect 59170 236898 59406 237134
rect 69410 237218 69646 237454
rect 69410 236898 69646 237134
rect 79650 237218 79886 237454
rect 79650 236898 79886 237134
rect 89890 237218 90126 237454
rect 89890 236898 90126 237134
rect 100130 237218 100366 237454
rect 100130 236898 100366 237134
rect 110370 237218 110606 237454
rect 110370 236898 110606 237134
rect 120610 237218 120846 237454
rect 120610 236898 120846 237134
rect 130850 237218 131086 237454
rect 130850 236898 131086 237134
rect 141090 237218 141326 237454
rect 141090 236898 141326 237134
rect 151330 237218 151566 237454
rect 151330 236898 151566 237134
rect 161570 237218 161806 237454
rect 161570 236898 161806 237134
rect 171810 237218 172046 237454
rect 171810 236898 172046 237134
rect 182050 237218 182286 237454
rect 182050 236898 182286 237134
rect 192290 237218 192526 237454
rect 192290 236898 192526 237134
rect 202530 237218 202766 237454
rect 202530 236898 202766 237134
rect 212770 237218 213006 237454
rect 212770 236898 213006 237134
rect 223010 237218 223246 237454
rect 223010 236898 223246 237134
rect 233250 237218 233486 237454
rect 233250 236898 233486 237134
rect 243490 237218 243726 237454
rect 243490 236898 243726 237134
rect 253730 237218 253966 237454
rect 253730 236898 253966 237134
rect 263970 237218 264206 237454
rect 263970 236898 264206 237134
rect 274210 237218 274446 237454
rect 274210 236898 274446 237134
rect 284450 237218 284686 237454
rect 284450 236898 284686 237134
rect 294690 237218 294926 237454
rect 294690 236898 294926 237134
rect 304930 237218 305166 237454
rect 304930 236898 305166 237134
rect 315170 237218 315406 237454
rect 315170 236898 315406 237134
rect 325410 237218 325646 237454
rect 325410 236898 325646 237134
rect 335650 237218 335886 237454
rect 335650 236898 335886 237134
rect 345890 237218 346126 237454
rect 345890 236898 346126 237134
rect 356130 237218 356366 237454
rect 356130 236898 356366 237134
rect 366370 237218 366606 237454
rect 366370 236898 366606 237134
rect 376610 237218 376846 237454
rect 376610 236898 376846 237134
rect 386850 237218 387086 237454
rect 386850 236898 387086 237134
rect 397090 237218 397326 237454
rect 397090 236898 397326 237134
rect 407330 237218 407566 237454
rect 407330 236898 407566 237134
rect 417570 237218 417806 237454
rect 417570 236898 417806 237134
rect 427810 237218 428046 237454
rect 427810 236898 428046 237134
rect 438050 237218 438286 237454
rect 438050 236898 438286 237134
rect 448290 237218 448526 237454
rect 448290 236898 448526 237134
rect 458530 237218 458766 237454
rect 458530 236898 458766 237134
rect 468770 237218 469006 237454
rect 468770 236898 469006 237134
rect 479010 237218 479246 237454
rect 479010 236898 479246 237134
rect 489250 237218 489486 237454
rect 489250 236898 489486 237134
rect 499490 237218 499726 237454
rect 499490 236898 499726 237134
rect 509730 237218 509966 237454
rect 509730 236898 509966 237134
rect 519970 237218 520206 237454
rect 519970 236898 520206 237134
rect 530210 237218 530446 237454
rect 530210 236898 530446 237134
rect 15786 222938 16022 223174
rect 16106 222938 16342 223174
rect 15786 222618 16022 222854
rect 16106 222618 16342 222854
rect 541746 226658 541982 226894
rect 542066 226658 542302 226894
rect 541746 226338 541982 226574
rect 542066 226338 542302 226574
rect 23330 219218 23566 219454
rect 23330 218898 23566 219134
rect 33570 219218 33806 219454
rect 33570 218898 33806 219134
rect 43810 219218 44046 219454
rect 43810 218898 44046 219134
rect 54050 219218 54286 219454
rect 54050 218898 54286 219134
rect 64290 219218 64526 219454
rect 64290 218898 64526 219134
rect 74530 219218 74766 219454
rect 74530 218898 74766 219134
rect 84770 219218 85006 219454
rect 84770 218898 85006 219134
rect 95010 219218 95246 219454
rect 95010 218898 95246 219134
rect 105250 219218 105486 219454
rect 105250 218898 105486 219134
rect 115490 219218 115726 219454
rect 115490 218898 115726 219134
rect 125730 219218 125966 219454
rect 125730 218898 125966 219134
rect 135970 219218 136206 219454
rect 135970 218898 136206 219134
rect 146210 219218 146446 219454
rect 146210 218898 146446 219134
rect 156450 219218 156686 219454
rect 156450 218898 156686 219134
rect 166690 219218 166926 219454
rect 166690 218898 166926 219134
rect 176930 219218 177166 219454
rect 176930 218898 177166 219134
rect 187170 219218 187406 219454
rect 187170 218898 187406 219134
rect 197410 219218 197646 219454
rect 197410 218898 197646 219134
rect 207650 219218 207886 219454
rect 207650 218898 207886 219134
rect 217890 219218 218126 219454
rect 217890 218898 218126 219134
rect 228130 219218 228366 219454
rect 228130 218898 228366 219134
rect 238370 219218 238606 219454
rect 238370 218898 238606 219134
rect 248610 219218 248846 219454
rect 248610 218898 248846 219134
rect 258850 219218 259086 219454
rect 258850 218898 259086 219134
rect 269090 219218 269326 219454
rect 269090 218898 269326 219134
rect 279330 219218 279566 219454
rect 279330 218898 279566 219134
rect 289570 219218 289806 219454
rect 289570 218898 289806 219134
rect 299810 219218 300046 219454
rect 299810 218898 300046 219134
rect 310050 219218 310286 219454
rect 310050 218898 310286 219134
rect 320290 219218 320526 219454
rect 320290 218898 320526 219134
rect 330530 219218 330766 219454
rect 330530 218898 330766 219134
rect 340770 219218 341006 219454
rect 340770 218898 341006 219134
rect 351010 219218 351246 219454
rect 351010 218898 351246 219134
rect 361250 219218 361486 219454
rect 361250 218898 361486 219134
rect 371490 219218 371726 219454
rect 371490 218898 371726 219134
rect 381730 219218 381966 219454
rect 381730 218898 381966 219134
rect 391970 219218 392206 219454
rect 391970 218898 392206 219134
rect 402210 219218 402446 219454
rect 402210 218898 402446 219134
rect 412450 219218 412686 219454
rect 412450 218898 412686 219134
rect 422690 219218 422926 219454
rect 422690 218898 422926 219134
rect 432930 219218 433166 219454
rect 432930 218898 433166 219134
rect 443170 219218 443406 219454
rect 443170 218898 443406 219134
rect 453410 219218 453646 219454
rect 453410 218898 453646 219134
rect 463650 219218 463886 219454
rect 463650 218898 463886 219134
rect 473890 219218 474126 219454
rect 473890 218898 474126 219134
rect 484130 219218 484366 219454
rect 484130 218898 484366 219134
rect 494370 219218 494606 219454
rect 494370 218898 494606 219134
rect 504610 219218 504846 219454
rect 504610 218898 504846 219134
rect 514850 219218 515086 219454
rect 514850 218898 515086 219134
rect 525090 219218 525326 219454
rect 525090 218898 525326 219134
rect 535330 219218 535566 219454
rect 535330 218898 535566 219134
rect 28450 201218 28686 201454
rect 28450 200898 28686 201134
rect 38690 201218 38926 201454
rect 38690 200898 38926 201134
rect 48930 201218 49166 201454
rect 48930 200898 49166 201134
rect 59170 201218 59406 201454
rect 59170 200898 59406 201134
rect 69410 201218 69646 201454
rect 69410 200898 69646 201134
rect 79650 201218 79886 201454
rect 79650 200898 79886 201134
rect 89890 201218 90126 201454
rect 89890 200898 90126 201134
rect 100130 201218 100366 201454
rect 100130 200898 100366 201134
rect 110370 201218 110606 201454
rect 110370 200898 110606 201134
rect 120610 201218 120846 201454
rect 120610 200898 120846 201134
rect 130850 201218 131086 201454
rect 130850 200898 131086 201134
rect 141090 201218 141326 201454
rect 141090 200898 141326 201134
rect 151330 201218 151566 201454
rect 151330 200898 151566 201134
rect 161570 201218 161806 201454
rect 161570 200898 161806 201134
rect 171810 201218 172046 201454
rect 171810 200898 172046 201134
rect 182050 201218 182286 201454
rect 182050 200898 182286 201134
rect 192290 201218 192526 201454
rect 192290 200898 192526 201134
rect 202530 201218 202766 201454
rect 202530 200898 202766 201134
rect 212770 201218 213006 201454
rect 212770 200898 213006 201134
rect 223010 201218 223246 201454
rect 223010 200898 223246 201134
rect 233250 201218 233486 201454
rect 233250 200898 233486 201134
rect 243490 201218 243726 201454
rect 243490 200898 243726 201134
rect 253730 201218 253966 201454
rect 253730 200898 253966 201134
rect 263970 201218 264206 201454
rect 263970 200898 264206 201134
rect 274210 201218 274446 201454
rect 274210 200898 274446 201134
rect 284450 201218 284686 201454
rect 284450 200898 284686 201134
rect 294690 201218 294926 201454
rect 294690 200898 294926 201134
rect 304930 201218 305166 201454
rect 304930 200898 305166 201134
rect 315170 201218 315406 201454
rect 315170 200898 315406 201134
rect 325410 201218 325646 201454
rect 325410 200898 325646 201134
rect 335650 201218 335886 201454
rect 335650 200898 335886 201134
rect 345890 201218 346126 201454
rect 345890 200898 346126 201134
rect 356130 201218 356366 201454
rect 356130 200898 356366 201134
rect 366370 201218 366606 201454
rect 366370 200898 366606 201134
rect 376610 201218 376846 201454
rect 376610 200898 376846 201134
rect 386850 201218 387086 201454
rect 386850 200898 387086 201134
rect 397090 201218 397326 201454
rect 397090 200898 397326 201134
rect 407330 201218 407566 201454
rect 407330 200898 407566 201134
rect 417570 201218 417806 201454
rect 417570 200898 417806 201134
rect 427810 201218 428046 201454
rect 427810 200898 428046 201134
rect 438050 201218 438286 201454
rect 438050 200898 438286 201134
rect 448290 201218 448526 201454
rect 448290 200898 448526 201134
rect 458530 201218 458766 201454
rect 458530 200898 458766 201134
rect 468770 201218 469006 201454
rect 468770 200898 469006 201134
rect 479010 201218 479246 201454
rect 479010 200898 479246 201134
rect 489250 201218 489486 201454
rect 489250 200898 489486 201134
rect 499490 201218 499726 201454
rect 499490 200898 499726 201134
rect 509730 201218 509966 201454
rect 509730 200898 509966 201134
rect 519970 201218 520206 201454
rect 519970 200898 520206 201134
rect 530210 201218 530446 201454
rect 530210 200898 530446 201134
rect 15786 186938 16022 187174
rect 16106 186938 16342 187174
rect 15786 186618 16022 186854
rect 16106 186618 16342 186854
rect 541746 190658 541982 190894
rect 542066 190658 542302 190894
rect 541746 190338 541982 190574
rect 542066 190338 542302 190574
rect 23330 183218 23566 183454
rect 23330 182898 23566 183134
rect 33570 183218 33806 183454
rect 33570 182898 33806 183134
rect 43810 183218 44046 183454
rect 43810 182898 44046 183134
rect 54050 183218 54286 183454
rect 54050 182898 54286 183134
rect 64290 183218 64526 183454
rect 64290 182898 64526 183134
rect 74530 183218 74766 183454
rect 74530 182898 74766 183134
rect 84770 183218 85006 183454
rect 84770 182898 85006 183134
rect 95010 183218 95246 183454
rect 95010 182898 95246 183134
rect 105250 183218 105486 183454
rect 105250 182898 105486 183134
rect 115490 183218 115726 183454
rect 115490 182898 115726 183134
rect 125730 183218 125966 183454
rect 125730 182898 125966 183134
rect 135970 183218 136206 183454
rect 135970 182898 136206 183134
rect 146210 183218 146446 183454
rect 146210 182898 146446 183134
rect 156450 183218 156686 183454
rect 156450 182898 156686 183134
rect 166690 183218 166926 183454
rect 166690 182898 166926 183134
rect 176930 183218 177166 183454
rect 176930 182898 177166 183134
rect 187170 183218 187406 183454
rect 187170 182898 187406 183134
rect 197410 183218 197646 183454
rect 197410 182898 197646 183134
rect 207650 183218 207886 183454
rect 207650 182898 207886 183134
rect 217890 183218 218126 183454
rect 217890 182898 218126 183134
rect 228130 183218 228366 183454
rect 228130 182898 228366 183134
rect 238370 183218 238606 183454
rect 238370 182898 238606 183134
rect 248610 183218 248846 183454
rect 248610 182898 248846 183134
rect 258850 183218 259086 183454
rect 258850 182898 259086 183134
rect 269090 183218 269326 183454
rect 269090 182898 269326 183134
rect 279330 183218 279566 183454
rect 279330 182898 279566 183134
rect 289570 183218 289806 183454
rect 289570 182898 289806 183134
rect 299810 183218 300046 183454
rect 299810 182898 300046 183134
rect 310050 183218 310286 183454
rect 310050 182898 310286 183134
rect 320290 183218 320526 183454
rect 320290 182898 320526 183134
rect 330530 183218 330766 183454
rect 330530 182898 330766 183134
rect 340770 183218 341006 183454
rect 340770 182898 341006 183134
rect 351010 183218 351246 183454
rect 351010 182898 351246 183134
rect 361250 183218 361486 183454
rect 361250 182898 361486 183134
rect 371490 183218 371726 183454
rect 371490 182898 371726 183134
rect 381730 183218 381966 183454
rect 381730 182898 381966 183134
rect 391970 183218 392206 183454
rect 391970 182898 392206 183134
rect 402210 183218 402446 183454
rect 402210 182898 402446 183134
rect 412450 183218 412686 183454
rect 412450 182898 412686 183134
rect 422690 183218 422926 183454
rect 422690 182898 422926 183134
rect 432930 183218 433166 183454
rect 432930 182898 433166 183134
rect 443170 183218 443406 183454
rect 443170 182898 443406 183134
rect 453410 183218 453646 183454
rect 453410 182898 453646 183134
rect 463650 183218 463886 183454
rect 463650 182898 463886 183134
rect 473890 183218 474126 183454
rect 473890 182898 474126 183134
rect 484130 183218 484366 183454
rect 484130 182898 484366 183134
rect 494370 183218 494606 183454
rect 494370 182898 494606 183134
rect 504610 183218 504846 183454
rect 504610 182898 504846 183134
rect 514850 183218 515086 183454
rect 514850 182898 515086 183134
rect 525090 183218 525326 183454
rect 525090 182898 525326 183134
rect 535330 183218 535566 183454
rect 535330 182898 535566 183134
rect 28450 165218 28686 165454
rect 28450 164898 28686 165134
rect 38690 165218 38926 165454
rect 38690 164898 38926 165134
rect 48930 165218 49166 165454
rect 48930 164898 49166 165134
rect 59170 165218 59406 165454
rect 59170 164898 59406 165134
rect 69410 165218 69646 165454
rect 69410 164898 69646 165134
rect 79650 165218 79886 165454
rect 79650 164898 79886 165134
rect 89890 165218 90126 165454
rect 89890 164898 90126 165134
rect 100130 165218 100366 165454
rect 100130 164898 100366 165134
rect 110370 165218 110606 165454
rect 110370 164898 110606 165134
rect 120610 165218 120846 165454
rect 120610 164898 120846 165134
rect 130850 165218 131086 165454
rect 130850 164898 131086 165134
rect 141090 165218 141326 165454
rect 141090 164898 141326 165134
rect 151330 165218 151566 165454
rect 151330 164898 151566 165134
rect 161570 165218 161806 165454
rect 161570 164898 161806 165134
rect 171810 165218 172046 165454
rect 171810 164898 172046 165134
rect 182050 165218 182286 165454
rect 182050 164898 182286 165134
rect 192290 165218 192526 165454
rect 192290 164898 192526 165134
rect 202530 165218 202766 165454
rect 202530 164898 202766 165134
rect 212770 165218 213006 165454
rect 212770 164898 213006 165134
rect 223010 165218 223246 165454
rect 223010 164898 223246 165134
rect 233250 165218 233486 165454
rect 233250 164898 233486 165134
rect 243490 165218 243726 165454
rect 243490 164898 243726 165134
rect 253730 165218 253966 165454
rect 253730 164898 253966 165134
rect 263970 165218 264206 165454
rect 263970 164898 264206 165134
rect 274210 165218 274446 165454
rect 274210 164898 274446 165134
rect 284450 165218 284686 165454
rect 284450 164898 284686 165134
rect 294690 165218 294926 165454
rect 294690 164898 294926 165134
rect 304930 165218 305166 165454
rect 304930 164898 305166 165134
rect 315170 165218 315406 165454
rect 315170 164898 315406 165134
rect 325410 165218 325646 165454
rect 325410 164898 325646 165134
rect 335650 165218 335886 165454
rect 335650 164898 335886 165134
rect 345890 165218 346126 165454
rect 345890 164898 346126 165134
rect 356130 165218 356366 165454
rect 356130 164898 356366 165134
rect 366370 165218 366606 165454
rect 366370 164898 366606 165134
rect 376610 165218 376846 165454
rect 376610 164898 376846 165134
rect 386850 165218 387086 165454
rect 386850 164898 387086 165134
rect 397090 165218 397326 165454
rect 397090 164898 397326 165134
rect 407330 165218 407566 165454
rect 407330 164898 407566 165134
rect 417570 165218 417806 165454
rect 417570 164898 417806 165134
rect 427810 165218 428046 165454
rect 427810 164898 428046 165134
rect 438050 165218 438286 165454
rect 438050 164898 438286 165134
rect 448290 165218 448526 165454
rect 448290 164898 448526 165134
rect 458530 165218 458766 165454
rect 458530 164898 458766 165134
rect 468770 165218 469006 165454
rect 468770 164898 469006 165134
rect 479010 165218 479246 165454
rect 479010 164898 479246 165134
rect 489250 165218 489486 165454
rect 489250 164898 489486 165134
rect 499490 165218 499726 165454
rect 499490 164898 499726 165134
rect 509730 165218 509966 165454
rect 509730 164898 509966 165134
rect 519970 165218 520206 165454
rect 519970 164898 520206 165134
rect 530210 165218 530446 165454
rect 530210 164898 530446 165134
rect 15786 150938 16022 151174
rect 16106 150938 16342 151174
rect 15786 150618 16022 150854
rect 16106 150618 16342 150854
rect 541746 154658 541982 154894
rect 542066 154658 542302 154894
rect 541746 154338 541982 154574
rect 542066 154338 542302 154574
rect 23330 147218 23566 147454
rect 23330 146898 23566 147134
rect 33570 147218 33806 147454
rect 33570 146898 33806 147134
rect 43810 147218 44046 147454
rect 43810 146898 44046 147134
rect 54050 147218 54286 147454
rect 54050 146898 54286 147134
rect 64290 147218 64526 147454
rect 64290 146898 64526 147134
rect 74530 147218 74766 147454
rect 74530 146898 74766 147134
rect 84770 147218 85006 147454
rect 84770 146898 85006 147134
rect 95010 147218 95246 147454
rect 95010 146898 95246 147134
rect 105250 147218 105486 147454
rect 105250 146898 105486 147134
rect 115490 147218 115726 147454
rect 115490 146898 115726 147134
rect 125730 147218 125966 147454
rect 125730 146898 125966 147134
rect 135970 147218 136206 147454
rect 135970 146898 136206 147134
rect 146210 147218 146446 147454
rect 146210 146898 146446 147134
rect 156450 147218 156686 147454
rect 156450 146898 156686 147134
rect 166690 147218 166926 147454
rect 166690 146898 166926 147134
rect 176930 147218 177166 147454
rect 176930 146898 177166 147134
rect 187170 147218 187406 147454
rect 187170 146898 187406 147134
rect 197410 147218 197646 147454
rect 197410 146898 197646 147134
rect 207650 147218 207886 147454
rect 207650 146898 207886 147134
rect 217890 147218 218126 147454
rect 217890 146898 218126 147134
rect 228130 147218 228366 147454
rect 228130 146898 228366 147134
rect 238370 147218 238606 147454
rect 238370 146898 238606 147134
rect 248610 147218 248846 147454
rect 248610 146898 248846 147134
rect 258850 147218 259086 147454
rect 258850 146898 259086 147134
rect 269090 147218 269326 147454
rect 269090 146898 269326 147134
rect 279330 147218 279566 147454
rect 279330 146898 279566 147134
rect 289570 147218 289806 147454
rect 289570 146898 289806 147134
rect 299810 147218 300046 147454
rect 299810 146898 300046 147134
rect 310050 147218 310286 147454
rect 310050 146898 310286 147134
rect 320290 147218 320526 147454
rect 320290 146898 320526 147134
rect 330530 147218 330766 147454
rect 330530 146898 330766 147134
rect 340770 147218 341006 147454
rect 340770 146898 341006 147134
rect 351010 147218 351246 147454
rect 351010 146898 351246 147134
rect 361250 147218 361486 147454
rect 361250 146898 361486 147134
rect 371490 147218 371726 147454
rect 371490 146898 371726 147134
rect 381730 147218 381966 147454
rect 381730 146898 381966 147134
rect 391970 147218 392206 147454
rect 391970 146898 392206 147134
rect 402210 147218 402446 147454
rect 402210 146898 402446 147134
rect 412450 147218 412686 147454
rect 412450 146898 412686 147134
rect 422690 147218 422926 147454
rect 422690 146898 422926 147134
rect 432930 147218 433166 147454
rect 432930 146898 433166 147134
rect 443170 147218 443406 147454
rect 443170 146898 443406 147134
rect 453410 147218 453646 147454
rect 453410 146898 453646 147134
rect 463650 147218 463886 147454
rect 463650 146898 463886 147134
rect 473890 147218 474126 147454
rect 473890 146898 474126 147134
rect 484130 147218 484366 147454
rect 484130 146898 484366 147134
rect 494370 147218 494606 147454
rect 494370 146898 494606 147134
rect 504610 147218 504846 147454
rect 504610 146898 504846 147134
rect 514850 147218 515086 147454
rect 514850 146898 515086 147134
rect 525090 147218 525326 147454
rect 525090 146898 525326 147134
rect 535330 147218 535566 147454
rect 535330 146898 535566 147134
rect 28450 129218 28686 129454
rect 28450 128898 28686 129134
rect 38690 129218 38926 129454
rect 38690 128898 38926 129134
rect 48930 129218 49166 129454
rect 48930 128898 49166 129134
rect 59170 129218 59406 129454
rect 59170 128898 59406 129134
rect 69410 129218 69646 129454
rect 69410 128898 69646 129134
rect 79650 129218 79886 129454
rect 79650 128898 79886 129134
rect 89890 129218 90126 129454
rect 89890 128898 90126 129134
rect 100130 129218 100366 129454
rect 100130 128898 100366 129134
rect 110370 129218 110606 129454
rect 110370 128898 110606 129134
rect 120610 129218 120846 129454
rect 120610 128898 120846 129134
rect 130850 129218 131086 129454
rect 130850 128898 131086 129134
rect 141090 129218 141326 129454
rect 141090 128898 141326 129134
rect 151330 129218 151566 129454
rect 151330 128898 151566 129134
rect 161570 129218 161806 129454
rect 161570 128898 161806 129134
rect 171810 129218 172046 129454
rect 171810 128898 172046 129134
rect 182050 129218 182286 129454
rect 182050 128898 182286 129134
rect 192290 129218 192526 129454
rect 192290 128898 192526 129134
rect 202530 129218 202766 129454
rect 202530 128898 202766 129134
rect 212770 129218 213006 129454
rect 212770 128898 213006 129134
rect 223010 129218 223246 129454
rect 223010 128898 223246 129134
rect 233250 129218 233486 129454
rect 233250 128898 233486 129134
rect 243490 129218 243726 129454
rect 243490 128898 243726 129134
rect 253730 129218 253966 129454
rect 253730 128898 253966 129134
rect 263970 129218 264206 129454
rect 263970 128898 264206 129134
rect 274210 129218 274446 129454
rect 274210 128898 274446 129134
rect 284450 129218 284686 129454
rect 284450 128898 284686 129134
rect 294690 129218 294926 129454
rect 294690 128898 294926 129134
rect 304930 129218 305166 129454
rect 304930 128898 305166 129134
rect 315170 129218 315406 129454
rect 315170 128898 315406 129134
rect 325410 129218 325646 129454
rect 325410 128898 325646 129134
rect 335650 129218 335886 129454
rect 335650 128898 335886 129134
rect 345890 129218 346126 129454
rect 345890 128898 346126 129134
rect 356130 129218 356366 129454
rect 356130 128898 356366 129134
rect 366370 129218 366606 129454
rect 366370 128898 366606 129134
rect 376610 129218 376846 129454
rect 376610 128898 376846 129134
rect 386850 129218 387086 129454
rect 386850 128898 387086 129134
rect 397090 129218 397326 129454
rect 397090 128898 397326 129134
rect 407330 129218 407566 129454
rect 407330 128898 407566 129134
rect 417570 129218 417806 129454
rect 417570 128898 417806 129134
rect 427810 129218 428046 129454
rect 427810 128898 428046 129134
rect 438050 129218 438286 129454
rect 438050 128898 438286 129134
rect 448290 129218 448526 129454
rect 448290 128898 448526 129134
rect 458530 129218 458766 129454
rect 458530 128898 458766 129134
rect 468770 129218 469006 129454
rect 468770 128898 469006 129134
rect 479010 129218 479246 129454
rect 479010 128898 479246 129134
rect 489250 129218 489486 129454
rect 489250 128898 489486 129134
rect 499490 129218 499726 129454
rect 499490 128898 499726 129134
rect 509730 129218 509966 129454
rect 509730 128898 509966 129134
rect 519970 129218 520206 129454
rect 519970 128898 520206 129134
rect 530210 129218 530446 129454
rect 530210 128898 530446 129134
rect 15786 114938 16022 115174
rect 16106 114938 16342 115174
rect 15786 114618 16022 114854
rect 16106 114618 16342 114854
rect 541746 118658 541982 118894
rect 542066 118658 542302 118894
rect 541746 118338 541982 118574
rect 542066 118338 542302 118574
rect 23330 111218 23566 111454
rect 23330 110898 23566 111134
rect 33570 111218 33806 111454
rect 33570 110898 33806 111134
rect 43810 111218 44046 111454
rect 43810 110898 44046 111134
rect 54050 111218 54286 111454
rect 54050 110898 54286 111134
rect 64290 111218 64526 111454
rect 64290 110898 64526 111134
rect 74530 111218 74766 111454
rect 74530 110898 74766 111134
rect 84770 111218 85006 111454
rect 84770 110898 85006 111134
rect 95010 111218 95246 111454
rect 95010 110898 95246 111134
rect 105250 111218 105486 111454
rect 105250 110898 105486 111134
rect 115490 111218 115726 111454
rect 115490 110898 115726 111134
rect 125730 111218 125966 111454
rect 125730 110898 125966 111134
rect 135970 111218 136206 111454
rect 135970 110898 136206 111134
rect 146210 111218 146446 111454
rect 146210 110898 146446 111134
rect 156450 111218 156686 111454
rect 156450 110898 156686 111134
rect 166690 111218 166926 111454
rect 166690 110898 166926 111134
rect 176930 111218 177166 111454
rect 176930 110898 177166 111134
rect 187170 111218 187406 111454
rect 187170 110898 187406 111134
rect 197410 111218 197646 111454
rect 197410 110898 197646 111134
rect 207650 111218 207886 111454
rect 207650 110898 207886 111134
rect 217890 111218 218126 111454
rect 217890 110898 218126 111134
rect 228130 111218 228366 111454
rect 228130 110898 228366 111134
rect 238370 111218 238606 111454
rect 238370 110898 238606 111134
rect 248610 111218 248846 111454
rect 248610 110898 248846 111134
rect 258850 111218 259086 111454
rect 258850 110898 259086 111134
rect 269090 111218 269326 111454
rect 269090 110898 269326 111134
rect 279330 111218 279566 111454
rect 279330 110898 279566 111134
rect 289570 111218 289806 111454
rect 289570 110898 289806 111134
rect 299810 111218 300046 111454
rect 299810 110898 300046 111134
rect 310050 111218 310286 111454
rect 310050 110898 310286 111134
rect 320290 111218 320526 111454
rect 320290 110898 320526 111134
rect 330530 111218 330766 111454
rect 330530 110898 330766 111134
rect 340770 111218 341006 111454
rect 340770 110898 341006 111134
rect 351010 111218 351246 111454
rect 351010 110898 351246 111134
rect 361250 111218 361486 111454
rect 361250 110898 361486 111134
rect 371490 111218 371726 111454
rect 371490 110898 371726 111134
rect 381730 111218 381966 111454
rect 381730 110898 381966 111134
rect 391970 111218 392206 111454
rect 391970 110898 392206 111134
rect 402210 111218 402446 111454
rect 402210 110898 402446 111134
rect 412450 111218 412686 111454
rect 412450 110898 412686 111134
rect 422690 111218 422926 111454
rect 422690 110898 422926 111134
rect 432930 111218 433166 111454
rect 432930 110898 433166 111134
rect 443170 111218 443406 111454
rect 443170 110898 443406 111134
rect 453410 111218 453646 111454
rect 453410 110898 453646 111134
rect 463650 111218 463886 111454
rect 463650 110898 463886 111134
rect 473890 111218 474126 111454
rect 473890 110898 474126 111134
rect 484130 111218 484366 111454
rect 484130 110898 484366 111134
rect 494370 111218 494606 111454
rect 494370 110898 494606 111134
rect 504610 111218 504846 111454
rect 504610 110898 504846 111134
rect 514850 111218 515086 111454
rect 514850 110898 515086 111134
rect 525090 111218 525326 111454
rect 525090 110898 525326 111134
rect 535330 111218 535566 111454
rect 535330 110898 535566 111134
rect 28450 93218 28686 93454
rect 28450 92898 28686 93134
rect 38690 93218 38926 93454
rect 38690 92898 38926 93134
rect 48930 93218 49166 93454
rect 48930 92898 49166 93134
rect 59170 93218 59406 93454
rect 59170 92898 59406 93134
rect 69410 93218 69646 93454
rect 69410 92898 69646 93134
rect 79650 93218 79886 93454
rect 79650 92898 79886 93134
rect 89890 93218 90126 93454
rect 89890 92898 90126 93134
rect 100130 93218 100366 93454
rect 100130 92898 100366 93134
rect 110370 93218 110606 93454
rect 110370 92898 110606 93134
rect 120610 93218 120846 93454
rect 120610 92898 120846 93134
rect 130850 93218 131086 93454
rect 130850 92898 131086 93134
rect 141090 93218 141326 93454
rect 141090 92898 141326 93134
rect 151330 93218 151566 93454
rect 151330 92898 151566 93134
rect 161570 93218 161806 93454
rect 161570 92898 161806 93134
rect 171810 93218 172046 93454
rect 171810 92898 172046 93134
rect 182050 93218 182286 93454
rect 182050 92898 182286 93134
rect 192290 93218 192526 93454
rect 192290 92898 192526 93134
rect 202530 93218 202766 93454
rect 202530 92898 202766 93134
rect 212770 93218 213006 93454
rect 212770 92898 213006 93134
rect 223010 93218 223246 93454
rect 223010 92898 223246 93134
rect 233250 93218 233486 93454
rect 233250 92898 233486 93134
rect 243490 93218 243726 93454
rect 243490 92898 243726 93134
rect 253730 93218 253966 93454
rect 253730 92898 253966 93134
rect 263970 93218 264206 93454
rect 263970 92898 264206 93134
rect 274210 93218 274446 93454
rect 274210 92898 274446 93134
rect 284450 93218 284686 93454
rect 284450 92898 284686 93134
rect 294690 93218 294926 93454
rect 294690 92898 294926 93134
rect 304930 93218 305166 93454
rect 304930 92898 305166 93134
rect 315170 93218 315406 93454
rect 315170 92898 315406 93134
rect 325410 93218 325646 93454
rect 325410 92898 325646 93134
rect 335650 93218 335886 93454
rect 335650 92898 335886 93134
rect 345890 93218 346126 93454
rect 345890 92898 346126 93134
rect 356130 93218 356366 93454
rect 356130 92898 356366 93134
rect 366370 93218 366606 93454
rect 366370 92898 366606 93134
rect 376610 93218 376846 93454
rect 376610 92898 376846 93134
rect 386850 93218 387086 93454
rect 386850 92898 387086 93134
rect 397090 93218 397326 93454
rect 397090 92898 397326 93134
rect 407330 93218 407566 93454
rect 407330 92898 407566 93134
rect 417570 93218 417806 93454
rect 417570 92898 417806 93134
rect 427810 93218 428046 93454
rect 427810 92898 428046 93134
rect 438050 93218 438286 93454
rect 438050 92898 438286 93134
rect 448290 93218 448526 93454
rect 448290 92898 448526 93134
rect 458530 93218 458766 93454
rect 458530 92898 458766 93134
rect 468770 93218 469006 93454
rect 468770 92898 469006 93134
rect 479010 93218 479246 93454
rect 479010 92898 479246 93134
rect 489250 93218 489486 93454
rect 489250 92898 489486 93134
rect 499490 93218 499726 93454
rect 499490 92898 499726 93134
rect 509730 93218 509966 93454
rect 509730 92898 509966 93134
rect 519970 93218 520206 93454
rect 519970 92898 520206 93134
rect 530210 93218 530446 93454
rect 530210 92898 530446 93134
rect 15786 78938 16022 79174
rect 16106 78938 16342 79174
rect 15786 78618 16022 78854
rect 16106 78618 16342 78854
rect 541746 82658 541982 82894
rect 542066 82658 542302 82894
rect 541746 82338 541982 82574
rect 542066 82338 542302 82574
rect 23330 75218 23566 75454
rect 23330 74898 23566 75134
rect 33570 75218 33806 75454
rect 33570 74898 33806 75134
rect 43810 75218 44046 75454
rect 43810 74898 44046 75134
rect 54050 75218 54286 75454
rect 54050 74898 54286 75134
rect 64290 75218 64526 75454
rect 64290 74898 64526 75134
rect 74530 75218 74766 75454
rect 74530 74898 74766 75134
rect 84770 75218 85006 75454
rect 84770 74898 85006 75134
rect 95010 75218 95246 75454
rect 95010 74898 95246 75134
rect 105250 75218 105486 75454
rect 105250 74898 105486 75134
rect 115490 75218 115726 75454
rect 115490 74898 115726 75134
rect 125730 75218 125966 75454
rect 125730 74898 125966 75134
rect 135970 75218 136206 75454
rect 135970 74898 136206 75134
rect 146210 75218 146446 75454
rect 146210 74898 146446 75134
rect 156450 75218 156686 75454
rect 156450 74898 156686 75134
rect 166690 75218 166926 75454
rect 166690 74898 166926 75134
rect 176930 75218 177166 75454
rect 176930 74898 177166 75134
rect 187170 75218 187406 75454
rect 187170 74898 187406 75134
rect 197410 75218 197646 75454
rect 197410 74898 197646 75134
rect 207650 75218 207886 75454
rect 207650 74898 207886 75134
rect 217890 75218 218126 75454
rect 217890 74898 218126 75134
rect 228130 75218 228366 75454
rect 228130 74898 228366 75134
rect 238370 75218 238606 75454
rect 238370 74898 238606 75134
rect 248610 75218 248846 75454
rect 248610 74898 248846 75134
rect 258850 75218 259086 75454
rect 258850 74898 259086 75134
rect 269090 75218 269326 75454
rect 269090 74898 269326 75134
rect 279330 75218 279566 75454
rect 279330 74898 279566 75134
rect 289570 75218 289806 75454
rect 289570 74898 289806 75134
rect 299810 75218 300046 75454
rect 299810 74898 300046 75134
rect 310050 75218 310286 75454
rect 310050 74898 310286 75134
rect 320290 75218 320526 75454
rect 320290 74898 320526 75134
rect 330530 75218 330766 75454
rect 330530 74898 330766 75134
rect 340770 75218 341006 75454
rect 340770 74898 341006 75134
rect 351010 75218 351246 75454
rect 351010 74898 351246 75134
rect 361250 75218 361486 75454
rect 361250 74898 361486 75134
rect 371490 75218 371726 75454
rect 371490 74898 371726 75134
rect 381730 75218 381966 75454
rect 381730 74898 381966 75134
rect 391970 75218 392206 75454
rect 391970 74898 392206 75134
rect 402210 75218 402446 75454
rect 402210 74898 402446 75134
rect 412450 75218 412686 75454
rect 412450 74898 412686 75134
rect 422690 75218 422926 75454
rect 422690 74898 422926 75134
rect 432930 75218 433166 75454
rect 432930 74898 433166 75134
rect 443170 75218 443406 75454
rect 443170 74898 443406 75134
rect 453410 75218 453646 75454
rect 453410 74898 453646 75134
rect 463650 75218 463886 75454
rect 463650 74898 463886 75134
rect 473890 75218 474126 75454
rect 473890 74898 474126 75134
rect 484130 75218 484366 75454
rect 484130 74898 484366 75134
rect 494370 75218 494606 75454
rect 494370 74898 494606 75134
rect 504610 75218 504846 75454
rect 504610 74898 504846 75134
rect 514850 75218 515086 75454
rect 514850 74898 515086 75134
rect 525090 75218 525326 75454
rect 525090 74898 525326 75134
rect 535330 75218 535566 75454
rect 535330 74898 535566 75134
rect 28450 57218 28686 57454
rect 28450 56898 28686 57134
rect 38690 57218 38926 57454
rect 38690 56898 38926 57134
rect 48930 57218 49166 57454
rect 48930 56898 49166 57134
rect 59170 57218 59406 57454
rect 59170 56898 59406 57134
rect 69410 57218 69646 57454
rect 69410 56898 69646 57134
rect 79650 57218 79886 57454
rect 79650 56898 79886 57134
rect 89890 57218 90126 57454
rect 89890 56898 90126 57134
rect 100130 57218 100366 57454
rect 100130 56898 100366 57134
rect 110370 57218 110606 57454
rect 110370 56898 110606 57134
rect 120610 57218 120846 57454
rect 120610 56898 120846 57134
rect 130850 57218 131086 57454
rect 130850 56898 131086 57134
rect 141090 57218 141326 57454
rect 141090 56898 141326 57134
rect 151330 57218 151566 57454
rect 151330 56898 151566 57134
rect 161570 57218 161806 57454
rect 161570 56898 161806 57134
rect 171810 57218 172046 57454
rect 171810 56898 172046 57134
rect 182050 57218 182286 57454
rect 182050 56898 182286 57134
rect 192290 57218 192526 57454
rect 192290 56898 192526 57134
rect 202530 57218 202766 57454
rect 202530 56898 202766 57134
rect 212770 57218 213006 57454
rect 212770 56898 213006 57134
rect 223010 57218 223246 57454
rect 223010 56898 223246 57134
rect 233250 57218 233486 57454
rect 233250 56898 233486 57134
rect 243490 57218 243726 57454
rect 243490 56898 243726 57134
rect 253730 57218 253966 57454
rect 253730 56898 253966 57134
rect 263970 57218 264206 57454
rect 263970 56898 264206 57134
rect 274210 57218 274446 57454
rect 274210 56898 274446 57134
rect 284450 57218 284686 57454
rect 284450 56898 284686 57134
rect 294690 57218 294926 57454
rect 294690 56898 294926 57134
rect 304930 57218 305166 57454
rect 304930 56898 305166 57134
rect 315170 57218 315406 57454
rect 315170 56898 315406 57134
rect 325410 57218 325646 57454
rect 325410 56898 325646 57134
rect 335650 57218 335886 57454
rect 335650 56898 335886 57134
rect 345890 57218 346126 57454
rect 345890 56898 346126 57134
rect 356130 57218 356366 57454
rect 356130 56898 356366 57134
rect 366370 57218 366606 57454
rect 366370 56898 366606 57134
rect 376610 57218 376846 57454
rect 376610 56898 376846 57134
rect 386850 57218 387086 57454
rect 386850 56898 387086 57134
rect 397090 57218 397326 57454
rect 397090 56898 397326 57134
rect 407330 57218 407566 57454
rect 407330 56898 407566 57134
rect 417570 57218 417806 57454
rect 417570 56898 417806 57134
rect 427810 57218 428046 57454
rect 427810 56898 428046 57134
rect 438050 57218 438286 57454
rect 438050 56898 438286 57134
rect 448290 57218 448526 57454
rect 448290 56898 448526 57134
rect 458530 57218 458766 57454
rect 458530 56898 458766 57134
rect 468770 57218 469006 57454
rect 468770 56898 469006 57134
rect 479010 57218 479246 57454
rect 479010 56898 479246 57134
rect 489250 57218 489486 57454
rect 489250 56898 489486 57134
rect 499490 57218 499726 57454
rect 499490 56898 499726 57134
rect 509730 57218 509966 57454
rect 509730 56898 509966 57134
rect 519970 57218 520206 57454
rect 519970 56898 520206 57134
rect 530210 57218 530446 57454
rect 530210 56898 530446 57134
rect 15786 42938 16022 43174
rect 16106 42938 16342 43174
rect 15786 42618 16022 42854
rect 16106 42618 16342 42854
rect 541746 46658 541982 46894
rect 542066 46658 542302 46894
rect 541746 46338 541982 46574
rect 542066 46338 542302 46574
rect 23330 39218 23566 39454
rect 23330 38898 23566 39134
rect 33570 39218 33806 39454
rect 33570 38898 33806 39134
rect 43810 39218 44046 39454
rect 43810 38898 44046 39134
rect 54050 39218 54286 39454
rect 54050 38898 54286 39134
rect 64290 39218 64526 39454
rect 64290 38898 64526 39134
rect 74530 39218 74766 39454
rect 74530 38898 74766 39134
rect 84770 39218 85006 39454
rect 84770 38898 85006 39134
rect 95010 39218 95246 39454
rect 95010 38898 95246 39134
rect 105250 39218 105486 39454
rect 105250 38898 105486 39134
rect 115490 39218 115726 39454
rect 115490 38898 115726 39134
rect 125730 39218 125966 39454
rect 125730 38898 125966 39134
rect 135970 39218 136206 39454
rect 135970 38898 136206 39134
rect 146210 39218 146446 39454
rect 146210 38898 146446 39134
rect 156450 39218 156686 39454
rect 156450 38898 156686 39134
rect 166690 39218 166926 39454
rect 166690 38898 166926 39134
rect 176930 39218 177166 39454
rect 176930 38898 177166 39134
rect 187170 39218 187406 39454
rect 187170 38898 187406 39134
rect 197410 39218 197646 39454
rect 197410 38898 197646 39134
rect 207650 39218 207886 39454
rect 207650 38898 207886 39134
rect 217890 39218 218126 39454
rect 217890 38898 218126 39134
rect 228130 39218 228366 39454
rect 228130 38898 228366 39134
rect 238370 39218 238606 39454
rect 238370 38898 238606 39134
rect 248610 39218 248846 39454
rect 248610 38898 248846 39134
rect 258850 39218 259086 39454
rect 258850 38898 259086 39134
rect 269090 39218 269326 39454
rect 269090 38898 269326 39134
rect 279330 39218 279566 39454
rect 279330 38898 279566 39134
rect 289570 39218 289806 39454
rect 289570 38898 289806 39134
rect 299810 39218 300046 39454
rect 299810 38898 300046 39134
rect 310050 39218 310286 39454
rect 310050 38898 310286 39134
rect 320290 39218 320526 39454
rect 320290 38898 320526 39134
rect 330530 39218 330766 39454
rect 330530 38898 330766 39134
rect 340770 39218 341006 39454
rect 340770 38898 341006 39134
rect 351010 39218 351246 39454
rect 351010 38898 351246 39134
rect 361250 39218 361486 39454
rect 361250 38898 361486 39134
rect 371490 39218 371726 39454
rect 371490 38898 371726 39134
rect 381730 39218 381966 39454
rect 381730 38898 381966 39134
rect 391970 39218 392206 39454
rect 391970 38898 392206 39134
rect 402210 39218 402446 39454
rect 402210 38898 402446 39134
rect 412450 39218 412686 39454
rect 412450 38898 412686 39134
rect 422690 39218 422926 39454
rect 422690 38898 422926 39134
rect 432930 39218 433166 39454
rect 432930 38898 433166 39134
rect 443170 39218 443406 39454
rect 443170 38898 443406 39134
rect 453410 39218 453646 39454
rect 453410 38898 453646 39134
rect 463650 39218 463886 39454
rect 463650 38898 463886 39134
rect 473890 39218 474126 39454
rect 473890 38898 474126 39134
rect 484130 39218 484366 39454
rect 484130 38898 484366 39134
rect 494370 39218 494606 39454
rect 494370 38898 494606 39134
rect 504610 39218 504846 39454
rect 504610 38898 504846 39134
rect 514850 39218 515086 39454
rect 514850 38898 515086 39134
rect 525090 39218 525326 39454
rect 525090 38898 525326 39134
rect 535330 39218 535566 39454
rect 535330 38898 535566 39134
rect 28450 21218 28686 21454
rect 28450 20898 28686 21134
rect 38690 21218 38926 21454
rect 38690 20898 38926 21134
rect 48930 21218 49166 21454
rect 48930 20898 49166 21134
rect 59170 21218 59406 21454
rect 59170 20898 59406 21134
rect 69410 21218 69646 21454
rect 69410 20898 69646 21134
rect 79650 21218 79886 21454
rect 79650 20898 79886 21134
rect 89890 21218 90126 21454
rect 89890 20898 90126 21134
rect 100130 21218 100366 21454
rect 100130 20898 100366 21134
rect 110370 21218 110606 21454
rect 110370 20898 110606 21134
rect 120610 21218 120846 21454
rect 120610 20898 120846 21134
rect 130850 21218 131086 21454
rect 130850 20898 131086 21134
rect 141090 21218 141326 21454
rect 141090 20898 141326 21134
rect 151330 21218 151566 21454
rect 151330 20898 151566 21134
rect 161570 21218 161806 21454
rect 161570 20898 161806 21134
rect 171810 21218 172046 21454
rect 171810 20898 172046 21134
rect 182050 21218 182286 21454
rect 182050 20898 182286 21134
rect 192290 21218 192526 21454
rect 192290 20898 192526 21134
rect 202530 21218 202766 21454
rect 202530 20898 202766 21134
rect 212770 21218 213006 21454
rect 212770 20898 213006 21134
rect 223010 21218 223246 21454
rect 223010 20898 223246 21134
rect 233250 21218 233486 21454
rect 233250 20898 233486 21134
rect 243490 21218 243726 21454
rect 243490 20898 243726 21134
rect 253730 21218 253966 21454
rect 253730 20898 253966 21134
rect 263970 21218 264206 21454
rect 263970 20898 264206 21134
rect 274210 21218 274446 21454
rect 274210 20898 274446 21134
rect 284450 21218 284686 21454
rect 284450 20898 284686 21134
rect 294690 21218 294926 21454
rect 294690 20898 294926 21134
rect 304930 21218 305166 21454
rect 304930 20898 305166 21134
rect 315170 21218 315406 21454
rect 315170 20898 315406 21134
rect 325410 21218 325646 21454
rect 325410 20898 325646 21134
rect 335650 21218 335886 21454
rect 335650 20898 335886 21134
rect 345890 21218 346126 21454
rect 345890 20898 346126 21134
rect 356130 21218 356366 21454
rect 356130 20898 356366 21134
rect 366370 21218 366606 21454
rect 366370 20898 366606 21134
rect 376610 21218 376846 21454
rect 376610 20898 376846 21134
rect 386850 21218 387086 21454
rect 386850 20898 387086 21134
rect 397090 21218 397326 21454
rect 397090 20898 397326 21134
rect 407330 21218 407566 21454
rect 407330 20898 407566 21134
rect 417570 21218 417806 21454
rect 417570 20898 417806 21134
rect 427810 21218 428046 21454
rect 427810 20898 428046 21134
rect 438050 21218 438286 21454
rect 438050 20898 438286 21134
rect 448290 21218 448526 21454
rect 448290 20898 448526 21134
rect 458530 21218 458766 21454
rect 458530 20898 458766 21134
rect 468770 21218 469006 21454
rect 468770 20898 469006 21134
rect 479010 21218 479246 21454
rect 479010 20898 479246 21134
rect 489250 21218 489486 21454
rect 489250 20898 489486 21134
rect 499490 21218 499726 21454
rect 499490 20898 499726 21134
rect 509730 21218 509966 21454
rect 509730 20898 509966 21134
rect 519970 21218 520206 21454
rect 519970 20898 520206 21134
rect 530210 21218 530446 21454
rect 530210 20898 530446 21134
rect 15786 6938 16022 7174
rect 16106 6938 16342 7174
rect 15786 6618 16022 6854
rect 16106 6618 16342 6854
rect 17186 -1542 17422 -1306
rect 17506 -1542 17742 -1306
rect 17186 -1862 17422 -1626
rect 17506 -1862 17742 -1626
rect 15786 -2502 16022 -2266
rect 16106 -2502 16342 -2266
rect 15786 -2822 16022 -2586
rect 16106 -2822 16342 -2586
rect 14386 -5382 14622 -5146
rect 14706 -5382 14942 -5146
rect 14386 -5702 14622 -5466
rect 14706 -5702 14942 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 19506 10658 19742 10894
rect 19826 10658 20062 10894
rect 19506 10338 19742 10574
rect 19826 10338 20062 10574
rect 22306 3218 22542 3454
rect 22626 3218 22862 3454
rect 22306 2898 22542 3134
rect 22626 2898 22862 3134
rect 22306 -582 22542 -346
rect 22626 -582 22862 -346
rect 22306 -902 22542 -666
rect 22626 -902 22862 -666
rect 20906 -3462 21142 -3226
rect 21226 -3462 21462 -3226
rect 20906 -3782 21142 -3546
rect 21226 -3782 21462 -3546
rect 19506 -4422 19742 -4186
rect 19826 -4422 20062 -4186
rect 19506 -4742 19742 -4506
rect 19826 -4742 20062 -4506
rect 18106 -7302 18342 -7066
rect 18426 -7302 18662 -7066
rect 18106 -7622 18342 -7386
rect 18426 -7622 18662 -7386
rect 26026 6938 26262 7174
rect 26346 6938 26582 7174
rect 26026 6618 26262 6854
rect 26346 6618 26582 6854
rect 27426 -1542 27662 -1306
rect 27746 -1542 27982 -1306
rect 27426 -1862 27662 -1626
rect 27746 -1862 27982 -1626
rect 26026 -2502 26262 -2266
rect 26346 -2502 26582 -2266
rect 26026 -2822 26262 -2586
rect 26346 -2822 26582 -2586
rect 24626 -5382 24862 -5146
rect 24946 -5382 25182 -5146
rect 24626 -5702 24862 -5466
rect 24946 -5702 25182 -5466
rect 23226 -6342 23462 -6106
rect 23546 -6342 23782 -6106
rect 23226 -6662 23462 -6426
rect 23546 -6662 23782 -6426
rect 29746 10658 29982 10894
rect 30066 10658 30302 10894
rect 29746 10338 29982 10574
rect 30066 10338 30302 10574
rect 32546 3218 32782 3454
rect 32866 3218 33102 3454
rect 32546 2898 32782 3134
rect 32866 2898 33102 3134
rect 32546 -582 32782 -346
rect 32866 -582 33102 -346
rect 32546 -902 32782 -666
rect 32866 -902 33102 -666
rect 31146 -3462 31382 -3226
rect 31466 -3462 31702 -3226
rect 31146 -3782 31382 -3546
rect 31466 -3782 31702 -3546
rect 29746 -4422 29982 -4186
rect 30066 -4422 30302 -4186
rect 29746 -4742 29982 -4506
rect 30066 -4742 30302 -4506
rect 28346 -7302 28582 -7066
rect 28666 -7302 28902 -7066
rect 28346 -7622 28582 -7386
rect 28666 -7622 28902 -7386
rect 36266 6938 36502 7174
rect 36586 6938 36822 7174
rect 36266 6618 36502 6854
rect 36586 6618 36822 6854
rect 37666 -1542 37902 -1306
rect 37986 -1542 38222 -1306
rect 37666 -1862 37902 -1626
rect 37986 -1862 38222 -1626
rect 36266 -2502 36502 -2266
rect 36586 -2502 36822 -2266
rect 36266 -2822 36502 -2586
rect 36586 -2822 36822 -2586
rect 34866 -5382 35102 -5146
rect 35186 -5382 35422 -5146
rect 34866 -5702 35102 -5466
rect 35186 -5702 35422 -5466
rect 33466 -6342 33702 -6106
rect 33786 -6342 34022 -6106
rect 33466 -6662 33702 -6426
rect 33786 -6662 34022 -6426
rect 39986 10658 40222 10894
rect 40306 10658 40542 10894
rect 39986 10338 40222 10574
rect 40306 10338 40542 10574
rect 42786 3218 43022 3454
rect 43106 3218 43342 3454
rect 42786 2898 43022 3134
rect 43106 2898 43342 3134
rect 42786 -582 43022 -346
rect 43106 -582 43342 -346
rect 42786 -902 43022 -666
rect 43106 -902 43342 -666
rect 41386 -3462 41622 -3226
rect 41706 -3462 41942 -3226
rect 41386 -3782 41622 -3546
rect 41706 -3782 41942 -3546
rect 39986 -4422 40222 -4186
rect 40306 -4422 40542 -4186
rect 39986 -4742 40222 -4506
rect 40306 -4742 40542 -4506
rect 38586 -7302 38822 -7066
rect 38906 -7302 39142 -7066
rect 38586 -7622 38822 -7386
rect 38906 -7622 39142 -7386
rect 46506 6938 46742 7174
rect 46826 6938 47062 7174
rect 46506 6618 46742 6854
rect 46826 6618 47062 6854
rect 47906 -1542 48142 -1306
rect 48226 -1542 48462 -1306
rect 47906 -1862 48142 -1626
rect 48226 -1862 48462 -1626
rect 46506 -2502 46742 -2266
rect 46826 -2502 47062 -2266
rect 46506 -2822 46742 -2586
rect 46826 -2822 47062 -2586
rect 45106 -5382 45342 -5146
rect 45426 -5382 45662 -5146
rect 45106 -5702 45342 -5466
rect 45426 -5702 45662 -5466
rect 43706 -6342 43942 -6106
rect 44026 -6342 44262 -6106
rect 43706 -6662 43942 -6426
rect 44026 -6662 44262 -6426
rect 50226 10658 50462 10894
rect 50546 10658 50782 10894
rect 50226 10338 50462 10574
rect 50546 10338 50782 10574
rect 53026 3218 53262 3454
rect 53346 3218 53582 3454
rect 53026 2898 53262 3134
rect 53346 2898 53582 3134
rect 53026 -582 53262 -346
rect 53346 -582 53582 -346
rect 53026 -902 53262 -666
rect 53346 -902 53582 -666
rect 51626 -3462 51862 -3226
rect 51946 -3462 52182 -3226
rect 51626 -3782 51862 -3546
rect 51946 -3782 52182 -3546
rect 50226 -4422 50462 -4186
rect 50546 -4422 50782 -4186
rect 50226 -4742 50462 -4506
rect 50546 -4742 50782 -4506
rect 48826 -7302 49062 -7066
rect 49146 -7302 49382 -7066
rect 48826 -7622 49062 -7386
rect 49146 -7622 49382 -7386
rect 56746 6938 56982 7174
rect 57066 6938 57302 7174
rect 56746 6618 56982 6854
rect 57066 6618 57302 6854
rect 58146 -1542 58382 -1306
rect 58466 -1542 58702 -1306
rect 58146 -1862 58382 -1626
rect 58466 -1862 58702 -1626
rect 56746 -2502 56982 -2266
rect 57066 -2502 57302 -2266
rect 56746 -2822 56982 -2586
rect 57066 -2822 57302 -2586
rect 55346 -5382 55582 -5146
rect 55666 -5382 55902 -5146
rect 55346 -5702 55582 -5466
rect 55666 -5702 55902 -5466
rect 53946 -6342 54182 -6106
rect 54266 -6342 54502 -6106
rect 53946 -6662 54182 -6426
rect 54266 -6662 54502 -6426
rect 60466 10658 60702 10894
rect 60786 10658 61022 10894
rect 60466 10338 60702 10574
rect 60786 10338 61022 10574
rect 63266 3218 63502 3454
rect 63586 3218 63822 3454
rect 63266 2898 63502 3134
rect 63586 2898 63822 3134
rect 63266 -582 63502 -346
rect 63586 -582 63822 -346
rect 63266 -902 63502 -666
rect 63586 -902 63822 -666
rect 61866 -3462 62102 -3226
rect 62186 -3462 62422 -3226
rect 61866 -3782 62102 -3546
rect 62186 -3782 62422 -3546
rect 60466 -4422 60702 -4186
rect 60786 -4422 61022 -4186
rect 60466 -4742 60702 -4506
rect 60786 -4742 61022 -4506
rect 59066 -7302 59302 -7066
rect 59386 -7302 59622 -7066
rect 59066 -7622 59302 -7386
rect 59386 -7622 59622 -7386
rect 66986 6938 67222 7174
rect 67306 6938 67542 7174
rect 66986 6618 67222 6854
rect 67306 6618 67542 6854
rect 68386 -1542 68622 -1306
rect 68706 -1542 68942 -1306
rect 68386 -1862 68622 -1626
rect 68706 -1862 68942 -1626
rect 66986 -2502 67222 -2266
rect 67306 -2502 67542 -2266
rect 66986 -2822 67222 -2586
rect 67306 -2822 67542 -2586
rect 65586 -5382 65822 -5146
rect 65906 -5382 66142 -5146
rect 65586 -5702 65822 -5466
rect 65906 -5702 66142 -5466
rect 64186 -6342 64422 -6106
rect 64506 -6342 64742 -6106
rect 64186 -6662 64422 -6426
rect 64506 -6662 64742 -6426
rect 70706 10658 70942 10894
rect 71026 10658 71262 10894
rect 70706 10338 70942 10574
rect 71026 10338 71262 10574
rect 73506 3218 73742 3454
rect 73826 3218 74062 3454
rect 73506 2898 73742 3134
rect 73826 2898 74062 3134
rect 73506 -582 73742 -346
rect 73826 -582 74062 -346
rect 73506 -902 73742 -666
rect 73826 -902 74062 -666
rect 72106 -3462 72342 -3226
rect 72426 -3462 72662 -3226
rect 72106 -3782 72342 -3546
rect 72426 -3782 72662 -3546
rect 70706 -4422 70942 -4186
rect 71026 -4422 71262 -4186
rect 70706 -4742 70942 -4506
rect 71026 -4742 71262 -4506
rect 69306 -7302 69542 -7066
rect 69626 -7302 69862 -7066
rect 69306 -7622 69542 -7386
rect 69626 -7622 69862 -7386
rect 77226 6938 77462 7174
rect 77546 6938 77782 7174
rect 77226 6618 77462 6854
rect 77546 6618 77782 6854
rect 78626 -1542 78862 -1306
rect 78946 -1542 79182 -1306
rect 78626 -1862 78862 -1626
rect 78946 -1862 79182 -1626
rect 77226 -2502 77462 -2266
rect 77546 -2502 77782 -2266
rect 77226 -2822 77462 -2586
rect 77546 -2822 77782 -2586
rect 75826 -5382 76062 -5146
rect 76146 -5382 76382 -5146
rect 75826 -5702 76062 -5466
rect 76146 -5702 76382 -5466
rect 74426 -6342 74662 -6106
rect 74746 -6342 74982 -6106
rect 74426 -6662 74662 -6426
rect 74746 -6662 74982 -6426
rect 80946 10658 81182 10894
rect 81266 10658 81502 10894
rect 80946 10338 81182 10574
rect 81266 10338 81502 10574
rect 83746 3218 83982 3454
rect 84066 3218 84302 3454
rect 83746 2898 83982 3134
rect 84066 2898 84302 3134
rect 83746 -582 83982 -346
rect 84066 -582 84302 -346
rect 83746 -902 83982 -666
rect 84066 -902 84302 -666
rect 82346 -3462 82582 -3226
rect 82666 -3462 82902 -3226
rect 82346 -3782 82582 -3546
rect 82666 -3782 82902 -3546
rect 80946 -4422 81182 -4186
rect 81266 -4422 81502 -4186
rect 80946 -4742 81182 -4506
rect 81266 -4742 81502 -4506
rect 79546 -7302 79782 -7066
rect 79866 -7302 80102 -7066
rect 79546 -7622 79782 -7386
rect 79866 -7622 80102 -7386
rect 87466 6938 87702 7174
rect 87786 6938 88022 7174
rect 87466 6618 87702 6854
rect 87786 6618 88022 6854
rect 88866 -1542 89102 -1306
rect 89186 -1542 89422 -1306
rect 88866 -1862 89102 -1626
rect 89186 -1862 89422 -1626
rect 87466 -2502 87702 -2266
rect 87786 -2502 88022 -2266
rect 87466 -2822 87702 -2586
rect 87786 -2822 88022 -2586
rect 86066 -5382 86302 -5146
rect 86386 -5382 86622 -5146
rect 86066 -5702 86302 -5466
rect 86386 -5702 86622 -5466
rect 84666 -6342 84902 -6106
rect 84986 -6342 85222 -6106
rect 84666 -6662 84902 -6426
rect 84986 -6662 85222 -6426
rect 91186 10658 91422 10894
rect 91506 10658 91742 10894
rect 91186 10338 91422 10574
rect 91506 10338 91742 10574
rect 93986 3218 94222 3454
rect 94306 3218 94542 3454
rect 93986 2898 94222 3134
rect 94306 2898 94542 3134
rect 93986 -582 94222 -346
rect 94306 -582 94542 -346
rect 93986 -902 94222 -666
rect 94306 -902 94542 -666
rect 92586 -3462 92822 -3226
rect 92906 -3462 93142 -3226
rect 92586 -3782 92822 -3546
rect 92906 -3782 93142 -3546
rect 91186 -4422 91422 -4186
rect 91506 -4422 91742 -4186
rect 91186 -4742 91422 -4506
rect 91506 -4742 91742 -4506
rect 89786 -7302 90022 -7066
rect 90106 -7302 90342 -7066
rect 89786 -7622 90022 -7386
rect 90106 -7622 90342 -7386
rect 97706 6938 97942 7174
rect 98026 6938 98262 7174
rect 97706 6618 97942 6854
rect 98026 6618 98262 6854
rect 99106 -1542 99342 -1306
rect 99426 -1542 99662 -1306
rect 99106 -1862 99342 -1626
rect 99426 -1862 99662 -1626
rect 97706 -2502 97942 -2266
rect 98026 -2502 98262 -2266
rect 97706 -2822 97942 -2586
rect 98026 -2822 98262 -2586
rect 96306 -5382 96542 -5146
rect 96626 -5382 96862 -5146
rect 96306 -5702 96542 -5466
rect 96626 -5702 96862 -5466
rect 94906 -6342 95142 -6106
rect 95226 -6342 95462 -6106
rect 94906 -6662 95142 -6426
rect 95226 -6662 95462 -6426
rect 101426 10658 101662 10894
rect 101746 10658 101982 10894
rect 101426 10338 101662 10574
rect 101746 10338 101982 10574
rect 104226 3218 104462 3454
rect 104546 3218 104782 3454
rect 104226 2898 104462 3134
rect 104546 2898 104782 3134
rect 104226 -582 104462 -346
rect 104546 -582 104782 -346
rect 104226 -902 104462 -666
rect 104546 -902 104782 -666
rect 102826 -3462 103062 -3226
rect 103146 -3462 103382 -3226
rect 102826 -3782 103062 -3546
rect 103146 -3782 103382 -3546
rect 101426 -4422 101662 -4186
rect 101746 -4422 101982 -4186
rect 101426 -4742 101662 -4506
rect 101746 -4742 101982 -4506
rect 100026 -7302 100262 -7066
rect 100346 -7302 100582 -7066
rect 100026 -7622 100262 -7386
rect 100346 -7622 100582 -7386
rect 107946 6938 108182 7174
rect 108266 6938 108502 7174
rect 107946 6618 108182 6854
rect 108266 6618 108502 6854
rect 109346 -1542 109582 -1306
rect 109666 -1542 109902 -1306
rect 109346 -1862 109582 -1626
rect 109666 -1862 109902 -1626
rect 107946 -2502 108182 -2266
rect 108266 -2502 108502 -2266
rect 107946 -2822 108182 -2586
rect 108266 -2822 108502 -2586
rect 106546 -5382 106782 -5146
rect 106866 -5382 107102 -5146
rect 106546 -5702 106782 -5466
rect 106866 -5702 107102 -5466
rect 105146 -6342 105382 -6106
rect 105466 -6342 105702 -6106
rect 105146 -6662 105382 -6426
rect 105466 -6662 105702 -6426
rect 111666 10658 111902 10894
rect 111986 10658 112222 10894
rect 111666 10338 111902 10574
rect 111986 10338 112222 10574
rect 114466 3218 114702 3454
rect 114786 3218 115022 3454
rect 114466 2898 114702 3134
rect 114786 2898 115022 3134
rect 114466 -582 114702 -346
rect 114786 -582 115022 -346
rect 114466 -902 114702 -666
rect 114786 -902 115022 -666
rect 113066 -3462 113302 -3226
rect 113386 -3462 113622 -3226
rect 113066 -3782 113302 -3546
rect 113386 -3782 113622 -3546
rect 111666 -4422 111902 -4186
rect 111986 -4422 112222 -4186
rect 111666 -4742 111902 -4506
rect 111986 -4742 112222 -4506
rect 110266 -7302 110502 -7066
rect 110586 -7302 110822 -7066
rect 110266 -7622 110502 -7386
rect 110586 -7622 110822 -7386
rect 118186 6938 118422 7174
rect 118506 6938 118742 7174
rect 118186 6618 118422 6854
rect 118506 6618 118742 6854
rect 119586 -1542 119822 -1306
rect 119906 -1542 120142 -1306
rect 119586 -1862 119822 -1626
rect 119906 -1862 120142 -1626
rect 118186 -2502 118422 -2266
rect 118506 -2502 118742 -2266
rect 118186 -2822 118422 -2586
rect 118506 -2822 118742 -2586
rect 116786 -5382 117022 -5146
rect 117106 -5382 117342 -5146
rect 116786 -5702 117022 -5466
rect 117106 -5702 117342 -5466
rect 115386 -6342 115622 -6106
rect 115706 -6342 115942 -6106
rect 115386 -6662 115622 -6426
rect 115706 -6662 115942 -6426
rect 121906 10658 122142 10894
rect 122226 10658 122462 10894
rect 121906 10338 122142 10574
rect 122226 10338 122462 10574
rect 124706 3218 124942 3454
rect 125026 3218 125262 3454
rect 124706 2898 124942 3134
rect 125026 2898 125262 3134
rect 124706 -582 124942 -346
rect 125026 -582 125262 -346
rect 124706 -902 124942 -666
rect 125026 -902 125262 -666
rect 123306 -3462 123542 -3226
rect 123626 -3462 123862 -3226
rect 123306 -3782 123542 -3546
rect 123626 -3782 123862 -3546
rect 121906 -4422 122142 -4186
rect 122226 -4422 122462 -4186
rect 121906 -4742 122142 -4506
rect 122226 -4742 122462 -4506
rect 120506 -7302 120742 -7066
rect 120826 -7302 121062 -7066
rect 120506 -7622 120742 -7386
rect 120826 -7622 121062 -7386
rect 128426 6938 128662 7174
rect 128746 6938 128982 7174
rect 128426 6618 128662 6854
rect 128746 6618 128982 6854
rect 129826 -1542 130062 -1306
rect 130146 -1542 130382 -1306
rect 129826 -1862 130062 -1626
rect 130146 -1862 130382 -1626
rect 128426 -2502 128662 -2266
rect 128746 -2502 128982 -2266
rect 128426 -2822 128662 -2586
rect 128746 -2822 128982 -2586
rect 127026 -5382 127262 -5146
rect 127346 -5382 127582 -5146
rect 127026 -5702 127262 -5466
rect 127346 -5702 127582 -5466
rect 125626 -6342 125862 -6106
rect 125946 -6342 126182 -6106
rect 125626 -6662 125862 -6426
rect 125946 -6662 126182 -6426
rect 132146 10658 132382 10894
rect 132466 10658 132702 10894
rect 132146 10338 132382 10574
rect 132466 10338 132702 10574
rect 134946 3218 135182 3454
rect 135266 3218 135502 3454
rect 134946 2898 135182 3134
rect 135266 2898 135502 3134
rect 134946 -582 135182 -346
rect 135266 -582 135502 -346
rect 134946 -902 135182 -666
rect 135266 -902 135502 -666
rect 133546 -3462 133782 -3226
rect 133866 -3462 134102 -3226
rect 133546 -3782 133782 -3546
rect 133866 -3782 134102 -3546
rect 132146 -4422 132382 -4186
rect 132466 -4422 132702 -4186
rect 132146 -4742 132382 -4506
rect 132466 -4742 132702 -4506
rect 130746 -7302 130982 -7066
rect 131066 -7302 131302 -7066
rect 130746 -7622 130982 -7386
rect 131066 -7622 131302 -7386
rect 138666 6938 138902 7174
rect 138986 6938 139222 7174
rect 138666 6618 138902 6854
rect 138986 6618 139222 6854
rect 140066 -1542 140302 -1306
rect 140386 -1542 140622 -1306
rect 140066 -1862 140302 -1626
rect 140386 -1862 140622 -1626
rect 138666 -2502 138902 -2266
rect 138986 -2502 139222 -2266
rect 138666 -2822 138902 -2586
rect 138986 -2822 139222 -2586
rect 137266 -5382 137502 -5146
rect 137586 -5382 137822 -5146
rect 137266 -5702 137502 -5466
rect 137586 -5702 137822 -5466
rect 135866 -6342 136102 -6106
rect 136186 -6342 136422 -6106
rect 135866 -6662 136102 -6426
rect 136186 -6662 136422 -6426
rect 142386 10658 142622 10894
rect 142706 10658 142942 10894
rect 142386 10338 142622 10574
rect 142706 10338 142942 10574
rect 145186 3218 145422 3454
rect 145506 3218 145742 3454
rect 145186 2898 145422 3134
rect 145506 2898 145742 3134
rect 145186 -582 145422 -346
rect 145506 -582 145742 -346
rect 145186 -902 145422 -666
rect 145506 -902 145742 -666
rect 143786 -3462 144022 -3226
rect 144106 -3462 144342 -3226
rect 143786 -3782 144022 -3546
rect 144106 -3782 144342 -3546
rect 142386 -4422 142622 -4186
rect 142706 -4422 142942 -4186
rect 142386 -4742 142622 -4506
rect 142706 -4742 142942 -4506
rect 140986 -7302 141222 -7066
rect 141306 -7302 141542 -7066
rect 140986 -7622 141222 -7386
rect 141306 -7622 141542 -7386
rect 148906 6938 149142 7174
rect 149226 6938 149462 7174
rect 148906 6618 149142 6854
rect 149226 6618 149462 6854
rect 150306 -1542 150542 -1306
rect 150626 -1542 150862 -1306
rect 150306 -1862 150542 -1626
rect 150626 -1862 150862 -1626
rect 148906 -2502 149142 -2266
rect 149226 -2502 149462 -2266
rect 148906 -2822 149142 -2586
rect 149226 -2822 149462 -2586
rect 147506 -5382 147742 -5146
rect 147826 -5382 148062 -5146
rect 147506 -5702 147742 -5466
rect 147826 -5702 148062 -5466
rect 146106 -6342 146342 -6106
rect 146426 -6342 146662 -6106
rect 146106 -6662 146342 -6426
rect 146426 -6662 146662 -6426
rect 152626 10658 152862 10894
rect 152946 10658 153182 10894
rect 152626 10338 152862 10574
rect 152946 10338 153182 10574
rect 155426 3218 155662 3454
rect 155746 3218 155982 3454
rect 155426 2898 155662 3134
rect 155746 2898 155982 3134
rect 155426 -582 155662 -346
rect 155746 -582 155982 -346
rect 155426 -902 155662 -666
rect 155746 -902 155982 -666
rect 154026 -3462 154262 -3226
rect 154346 -3462 154582 -3226
rect 154026 -3782 154262 -3546
rect 154346 -3782 154582 -3546
rect 152626 -4422 152862 -4186
rect 152946 -4422 153182 -4186
rect 152626 -4742 152862 -4506
rect 152946 -4742 153182 -4506
rect 151226 -7302 151462 -7066
rect 151546 -7302 151782 -7066
rect 151226 -7622 151462 -7386
rect 151546 -7622 151782 -7386
rect 159146 6938 159382 7174
rect 159466 6938 159702 7174
rect 159146 6618 159382 6854
rect 159466 6618 159702 6854
rect 160546 -1542 160782 -1306
rect 160866 -1542 161102 -1306
rect 160546 -1862 160782 -1626
rect 160866 -1862 161102 -1626
rect 159146 -2502 159382 -2266
rect 159466 -2502 159702 -2266
rect 159146 -2822 159382 -2586
rect 159466 -2822 159702 -2586
rect 157746 -5382 157982 -5146
rect 158066 -5382 158302 -5146
rect 157746 -5702 157982 -5466
rect 158066 -5702 158302 -5466
rect 156346 -6342 156582 -6106
rect 156666 -6342 156902 -6106
rect 156346 -6662 156582 -6426
rect 156666 -6662 156902 -6426
rect 162866 10658 163102 10894
rect 163186 10658 163422 10894
rect 162866 10338 163102 10574
rect 163186 10338 163422 10574
rect 165666 3218 165902 3454
rect 165986 3218 166222 3454
rect 165666 2898 165902 3134
rect 165986 2898 166222 3134
rect 165666 -582 165902 -346
rect 165986 -582 166222 -346
rect 165666 -902 165902 -666
rect 165986 -902 166222 -666
rect 164266 -3462 164502 -3226
rect 164586 -3462 164822 -3226
rect 164266 -3782 164502 -3546
rect 164586 -3782 164822 -3546
rect 162866 -4422 163102 -4186
rect 163186 -4422 163422 -4186
rect 162866 -4742 163102 -4506
rect 163186 -4742 163422 -4506
rect 161466 -7302 161702 -7066
rect 161786 -7302 162022 -7066
rect 161466 -7622 161702 -7386
rect 161786 -7622 162022 -7386
rect 169386 6938 169622 7174
rect 169706 6938 169942 7174
rect 169386 6618 169622 6854
rect 169706 6618 169942 6854
rect 170786 -1542 171022 -1306
rect 171106 -1542 171342 -1306
rect 170786 -1862 171022 -1626
rect 171106 -1862 171342 -1626
rect 169386 -2502 169622 -2266
rect 169706 -2502 169942 -2266
rect 169386 -2822 169622 -2586
rect 169706 -2822 169942 -2586
rect 167986 -5382 168222 -5146
rect 168306 -5382 168542 -5146
rect 167986 -5702 168222 -5466
rect 168306 -5702 168542 -5466
rect 166586 -6342 166822 -6106
rect 166906 -6342 167142 -6106
rect 166586 -6662 166822 -6426
rect 166906 -6662 167142 -6426
rect 173106 10658 173342 10894
rect 173426 10658 173662 10894
rect 173106 10338 173342 10574
rect 173426 10338 173662 10574
rect 175906 3218 176142 3454
rect 176226 3218 176462 3454
rect 175906 2898 176142 3134
rect 176226 2898 176462 3134
rect 175906 -582 176142 -346
rect 176226 -582 176462 -346
rect 175906 -902 176142 -666
rect 176226 -902 176462 -666
rect 174506 -3462 174742 -3226
rect 174826 -3462 175062 -3226
rect 174506 -3782 174742 -3546
rect 174826 -3782 175062 -3546
rect 173106 -4422 173342 -4186
rect 173426 -4422 173662 -4186
rect 173106 -4742 173342 -4506
rect 173426 -4742 173662 -4506
rect 171706 -7302 171942 -7066
rect 172026 -7302 172262 -7066
rect 171706 -7622 171942 -7386
rect 172026 -7622 172262 -7386
rect 179626 6938 179862 7174
rect 179946 6938 180182 7174
rect 179626 6618 179862 6854
rect 179946 6618 180182 6854
rect 181026 -1542 181262 -1306
rect 181346 -1542 181582 -1306
rect 181026 -1862 181262 -1626
rect 181346 -1862 181582 -1626
rect 179626 -2502 179862 -2266
rect 179946 -2502 180182 -2266
rect 179626 -2822 179862 -2586
rect 179946 -2822 180182 -2586
rect 178226 -5382 178462 -5146
rect 178546 -5382 178782 -5146
rect 178226 -5702 178462 -5466
rect 178546 -5702 178782 -5466
rect 176826 -6342 177062 -6106
rect 177146 -6342 177382 -6106
rect 176826 -6662 177062 -6426
rect 177146 -6662 177382 -6426
rect 183346 10658 183582 10894
rect 183666 10658 183902 10894
rect 183346 10338 183582 10574
rect 183666 10338 183902 10574
rect 186146 3218 186382 3454
rect 186466 3218 186702 3454
rect 186146 2898 186382 3134
rect 186466 2898 186702 3134
rect 186146 -582 186382 -346
rect 186466 -582 186702 -346
rect 186146 -902 186382 -666
rect 186466 -902 186702 -666
rect 184746 -3462 184982 -3226
rect 185066 -3462 185302 -3226
rect 184746 -3782 184982 -3546
rect 185066 -3782 185302 -3546
rect 183346 -4422 183582 -4186
rect 183666 -4422 183902 -4186
rect 183346 -4742 183582 -4506
rect 183666 -4742 183902 -4506
rect 181946 -7302 182182 -7066
rect 182266 -7302 182502 -7066
rect 181946 -7622 182182 -7386
rect 182266 -7622 182502 -7386
rect 189866 6938 190102 7174
rect 190186 6938 190422 7174
rect 189866 6618 190102 6854
rect 190186 6618 190422 6854
rect 191266 -1542 191502 -1306
rect 191586 -1542 191822 -1306
rect 191266 -1862 191502 -1626
rect 191586 -1862 191822 -1626
rect 189866 -2502 190102 -2266
rect 190186 -2502 190422 -2266
rect 189866 -2822 190102 -2586
rect 190186 -2822 190422 -2586
rect 188466 -5382 188702 -5146
rect 188786 -5382 189022 -5146
rect 188466 -5702 188702 -5466
rect 188786 -5702 189022 -5466
rect 187066 -6342 187302 -6106
rect 187386 -6342 187622 -6106
rect 187066 -6662 187302 -6426
rect 187386 -6662 187622 -6426
rect 193586 10658 193822 10894
rect 193906 10658 194142 10894
rect 193586 10338 193822 10574
rect 193906 10338 194142 10574
rect 196386 3218 196622 3454
rect 196706 3218 196942 3454
rect 196386 2898 196622 3134
rect 196706 2898 196942 3134
rect 196386 -582 196622 -346
rect 196706 -582 196942 -346
rect 196386 -902 196622 -666
rect 196706 -902 196942 -666
rect 194986 -3462 195222 -3226
rect 195306 -3462 195542 -3226
rect 194986 -3782 195222 -3546
rect 195306 -3782 195542 -3546
rect 193586 -4422 193822 -4186
rect 193906 -4422 194142 -4186
rect 193586 -4742 193822 -4506
rect 193906 -4742 194142 -4506
rect 192186 -7302 192422 -7066
rect 192506 -7302 192742 -7066
rect 192186 -7622 192422 -7386
rect 192506 -7622 192742 -7386
rect 200106 6938 200342 7174
rect 200426 6938 200662 7174
rect 200106 6618 200342 6854
rect 200426 6618 200662 6854
rect 201506 -1542 201742 -1306
rect 201826 -1542 202062 -1306
rect 201506 -1862 201742 -1626
rect 201826 -1862 202062 -1626
rect 200106 -2502 200342 -2266
rect 200426 -2502 200662 -2266
rect 200106 -2822 200342 -2586
rect 200426 -2822 200662 -2586
rect 198706 -5382 198942 -5146
rect 199026 -5382 199262 -5146
rect 198706 -5702 198942 -5466
rect 199026 -5702 199262 -5466
rect 197306 -6342 197542 -6106
rect 197626 -6342 197862 -6106
rect 197306 -6662 197542 -6426
rect 197626 -6662 197862 -6426
rect 203826 10658 204062 10894
rect 204146 10658 204382 10894
rect 203826 10338 204062 10574
rect 204146 10338 204382 10574
rect 206626 3218 206862 3454
rect 206946 3218 207182 3454
rect 206626 2898 206862 3134
rect 206946 2898 207182 3134
rect 206626 -582 206862 -346
rect 206946 -582 207182 -346
rect 206626 -902 206862 -666
rect 206946 -902 207182 -666
rect 205226 -3462 205462 -3226
rect 205546 -3462 205782 -3226
rect 205226 -3782 205462 -3546
rect 205546 -3782 205782 -3546
rect 203826 -4422 204062 -4186
rect 204146 -4422 204382 -4186
rect 203826 -4742 204062 -4506
rect 204146 -4742 204382 -4506
rect 202426 -7302 202662 -7066
rect 202746 -7302 202982 -7066
rect 202426 -7622 202662 -7386
rect 202746 -7622 202982 -7386
rect 210346 6938 210582 7174
rect 210666 6938 210902 7174
rect 210346 6618 210582 6854
rect 210666 6618 210902 6854
rect 211746 -1542 211982 -1306
rect 212066 -1542 212302 -1306
rect 211746 -1862 211982 -1626
rect 212066 -1862 212302 -1626
rect 210346 -2502 210582 -2266
rect 210666 -2502 210902 -2266
rect 210346 -2822 210582 -2586
rect 210666 -2822 210902 -2586
rect 208946 -5382 209182 -5146
rect 209266 -5382 209502 -5146
rect 208946 -5702 209182 -5466
rect 209266 -5702 209502 -5466
rect 207546 -6342 207782 -6106
rect 207866 -6342 208102 -6106
rect 207546 -6662 207782 -6426
rect 207866 -6662 208102 -6426
rect 214066 10658 214302 10894
rect 214386 10658 214622 10894
rect 214066 10338 214302 10574
rect 214386 10338 214622 10574
rect 216866 3218 217102 3454
rect 217186 3218 217422 3454
rect 216866 2898 217102 3134
rect 217186 2898 217422 3134
rect 216866 -582 217102 -346
rect 217186 -582 217422 -346
rect 216866 -902 217102 -666
rect 217186 -902 217422 -666
rect 215466 -3462 215702 -3226
rect 215786 -3462 216022 -3226
rect 215466 -3782 215702 -3546
rect 215786 -3782 216022 -3546
rect 214066 -4422 214302 -4186
rect 214386 -4422 214622 -4186
rect 214066 -4742 214302 -4506
rect 214386 -4742 214622 -4506
rect 212666 -7302 212902 -7066
rect 212986 -7302 213222 -7066
rect 212666 -7622 212902 -7386
rect 212986 -7622 213222 -7386
rect 220586 6938 220822 7174
rect 220906 6938 221142 7174
rect 220586 6618 220822 6854
rect 220906 6618 221142 6854
rect 221986 -1542 222222 -1306
rect 222306 -1542 222542 -1306
rect 221986 -1862 222222 -1626
rect 222306 -1862 222542 -1626
rect 220586 -2502 220822 -2266
rect 220906 -2502 221142 -2266
rect 220586 -2822 220822 -2586
rect 220906 -2822 221142 -2586
rect 219186 -5382 219422 -5146
rect 219506 -5382 219742 -5146
rect 219186 -5702 219422 -5466
rect 219506 -5702 219742 -5466
rect 217786 -6342 218022 -6106
rect 218106 -6342 218342 -6106
rect 217786 -6662 218022 -6426
rect 218106 -6662 218342 -6426
rect 224306 10658 224542 10894
rect 224626 10658 224862 10894
rect 224306 10338 224542 10574
rect 224626 10338 224862 10574
rect 227106 3218 227342 3454
rect 227426 3218 227662 3454
rect 227106 2898 227342 3134
rect 227426 2898 227662 3134
rect 227106 -582 227342 -346
rect 227426 -582 227662 -346
rect 227106 -902 227342 -666
rect 227426 -902 227662 -666
rect 225706 -3462 225942 -3226
rect 226026 -3462 226262 -3226
rect 225706 -3782 225942 -3546
rect 226026 -3782 226262 -3546
rect 224306 -4422 224542 -4186
rect 224626 -4422 224862 -4186
rect 224306 -4742 224542 -4506
rect 224626 -4742 224862 -4506
rect 222906 -7302 223142 -7066
rect 223226 -7302 223462 -7066
rect 222906 -7622 223142 -7386
rect 223226 -7622 223462 -7386
rect 230826 6938 231062 7174
rect 231146 6938 231382 7174
rect 230826 6618 231062 6854
rect 231146 6618 231382 6854
rect 232226 -1542 232462 -1306
rect 232546 -1542 232782 -1306
rect 232226 -1862 232462 -1626
rect 232546 -1862 232782 -1626
rect 230826 -2502 231062 -2266
rect 231146 -2502 231382 -2266
rect 230826 -2822 231062 -2586
rect 231146 -2822 231382 -2586
rect 229426 -5382 229662 -5146
rect 229746 -5382 229982 -5146
rect 229426 -5702 229662 -5466
rect 229746 -5702 229982 -5466
rect 228026 -6342 228262 -6106
rect 228346 -6342 228582 -6106
rect 228026 -6662 228262 -6426
rect 228346 -6662 228582 -6426
rect 234546 10658 234782 10894
rect 234866 10658 235102 10894
rect 234546 10338 234782 10574
rect 234866 10338 235102 10574
rect 237346 3218 237582 3454
rect 237666 3218 237902 3454
rect 237346 2898 237582 3134
rect 237666 2898 237902 3134
rect 237346 -582 237582 -346
rect 237666 -582 237902 -346
rect 237346 -902 237582 -666
rect 237666 -902 237902 -666
rect 235946 -3462 236182 -3226
rect 236266 -3462 236502 -3226
rect 235946 -3782 236182 -3546
rect 236266 -3782 236502 -3546
rect 234546 -4422 234782 -4186
rect 234866 -4422 235102 -4186
rect 234546 -4742 234782 -4506
rect 234866 -4742 235102 -4506
rect 233146 -7302 233382 -7066
rect 233466 -7302 233702 -7066
rect 233146 -7622 233382 -7386
rect 233466 -7622 233702 -7386
rect 241066 6938 241302 7174
rect 241386 6938 241622 7174
rect 241066 6618 241302 6854
rect 241386 6618 241622 6854
rect 242466 -1542 242702 -1306
rect 242786 -1542 243022 -1306
rect 242466 -1862 242702 -1626
rect 242786 -1862 243022 -1626
rect 241066 -2502 241302 -2266
rect 241386 -2502 241622 -2266
rect 241066 -2822 241302 -2586
rect 241386 -2822 241622 -2586
rect 239666 -5382 239902 -5146
rect 239986 -5382 240222 -5146
rect 239666 -5702 239902 -5466
rect 239986 -5702 240222 -5466
rect 238266 -6342 238502 -6106
rect 238586 -6342 238822 -6106
rect 238266 -6662 238502 -6426
rect 238586 -6662 238822 -6426
rect 244786 10658 245022 10894
rect 245106 10658 245342 10894
rect 244786 10338 245022 10574
rect 245106 10338 245342 10574
rect 247586 3218 247822 3454
rect 247906 3218 248142 3454
rect 247586 2898 247822 3134
rect 247906 2898 248142 3134
rect 247586 -582 247822 -346
rect 247906 -582 248142 -346
rect 247586 -902 247822 -666
rect 247906 -902 248142 -666
rect 246186 -3462 246422 -3226
rect 246506 -3462 246742 -3226
rect 246186 -3782 246422 -3546
rect 246506 -3782 246742 -3546
rect 244786 -4422 245022 -4186
rect 245106 -4422 245342 -4186
rect 244786 -4742 245022 -4506
rect 245106 -4742 245342 -4506
rect 243386 -7302 243622 -7066
rect 243706 -7302 243942 -7066
rect 243386 -7622 243622 -7386
rect 243706 -7622 243942 -7386
rect 251306 6938 251542 7174
rect 251626 6938 251862 7174
rect 251306 6618 251542 6854
rect 251626 6618 251862 6854
rect 252706 -1542 252942 -1306
rect 253026 -1542 253262 -1306
rect 252706 -1862 252942 -1626
rect 253026 -1862 253262 -1626
rect 251306 -2502 251542 -2266
rect 251626 -2502 251862 -2266
rect 251306 -2822 251542 -2586
rect 251626 -2822 251862 -2586
rect 249906 -5382 250142 -5146
rect 250226 -5382 250462 -5146
rect 249906 -5702 250142 -5466
rect 250226 -5702 250462 -5466
rect 248506 -6342 248742 -6106
rect 248826 -6342 249062 -6106
rect 248506 -6662 248742 -6426
rect 248826 -6662 249062 -6426
rect 255026 10658 255262 10894
rect 255346 10658 255582 10894
rect 255026 10338 255262 10574
rect 255346 10338 255582 10574
rect 257826 3218 258062 3454
rect 258146 3218 258382 3454
rect 257826 2898 258062 3134
rect 258146 2898 258382 3134
rect 257826 -582 258062 -346
rect 258146 -582 258382 -346
rect 257826 -902 258062 -666
rect 258146 -902 258382 -666
rect 256426 -3462 256662 -3226
rect 256746 -3462 256982 -3226
rect 256426 -3782 256662 -3546
rect 256746 -3782 256982 -3546
rect 255026 -4422 255262 -4186
rect 255346 -4422 255582 -4186
rect 255026 -4742 255262 -4506
rect 255346 -4742 255582 -4506
rect 253626 -7302 253862 -7066
rect 253946 -7302 254182 -7066
rect 253626 -7622 253862 -7386
rect 253946 -7622 254182 -7386
rect 261546 6938 261782 7174
rect 261866 6938 262102 7174
rect 261546 6618 261782 6854
rect 261866 6618 262102 6854
rect 262946 -1542 263182 -1306
rect 263266 -1542 263502 -1306
rect 262946 -1862 263182 -1626
rect 263266 -1862 263502 -1626
rect 261546 -2502 261782 -2266
rect 261866 -2502 262102 -2266
rect 261546 -2822 261782 -2586
rect 261866 -2822 262102 -2586
rect 260146 -5382 260382 -5146
rect 260466 -5382 260702 -5146
rect 260146 -5702 260382 -5466
rect 260466 -5702 260702 -5466
rect 258746 -6342 258982 -6106
rect 259066 -6342 259302 -6106
rect 258746 -6662 258982 -6426
rect 259066 -6662 259302 -6426
rect 265266 10658 265502 10894
rect 265586 10658 265822 10894
rect 265266 10338 265502 10574
rect 265586 10338 265822 10574
rect 268066 3218 268302 3454
rect 268386 3218 268622 3454
rect 268066 2898 268302 3134
rect 268386 2898 268622 3134
rect 268066 -582 268302 -346
rect 268386 -582 268622 -346
rect 268066 -902 268302 -666
rect 268386 -902 268622 -666
rect 266666 -3462 266902 -3226
rect 266986 -3462 267222 -3226
rect 266666 -3782 266902 -3546
rect 266986 -3782 267222 -3546
rect 265266 -4422 265502 -4186
rect 265586 -4422 265822 -4186
rect 265266 -4742 265502 -4506
rect 265586 -4742 265822 -4506
rect 263866 -7302 264102 -7066
rect 264186 -7302 264422 -7066
rect 263866 -7622 264102 -7386
rect 264186 -7622 264422 -7386
rect 271786 6938 272022 7174
rect 272106 6938 272342 7174
rect 271786 6618 272022 6854
rect 272106 6618 272342 6854
rect 273186 -1542 273422 -1306
rect 273506 -1542 273742 -1306
rect 273186 -1862 273422 -1626
rect 273506 -1862 273742 -1626
rect 271786 -2502 272022 -2266
rect 272106 -2502 272342 -2266
rect 271786 -2822 272022 -2586
rect 272106 -2822 272342 -2586
rect 270386 -5382 270622 -5146
rect 270706 -5382 270942 -5146
rect 270386 -5702 270622 -5466
rect 270706 -5702 270942 -5466
rect 268986 -6342 269222 -6106
rect 269306 -6342 269542 -6106
rect 268986 -6662 269222 -6426
rect 269306 -6662 269542 -6426
rect 275506 10658 275742 10894
rect 275826 10658 276062 10894
rect 275506 10338 275742 10574
rect 275826 10338 276062 10574
rect 278306 3218 278542 3454
rect 278626 3218 278862 3454
rect 278306 2898 278542 3134
rect 278626 2898 278862 3134
rect 278306 -582 278542 -346
rect 278626 -582 278862 -346
rect 278306 -902 278542 -666
rect 278626 -902 278862 -666
rect 276906 -3462 277142 -3226
rect 277226 -3462 277462 -3226
rect 276906 -3782 277142 -3546
rect 277226 -3782 277462 -3546
rect 275506 -4422 275742 -4186
rect 275826 -4422 276062 -4186
rect 275506 -4742 275742 -4506
rect 275826 -4742 276062 -4506
rect 274106 -7302 274342 -7066
rect 274426 -7302 274662 -7066
rect 274106 -7622 274342 -7386
rect 274426 -7622 274662 -7386
rect 282026 6938 282262 7174
rect 282346 6938 282582 7174
rect 282026 6618 282262 6854
rect 282346 6618 282582 6854
rect 283426 -1542 283662 -1306
rect 283746 -1542 283982 -1306
rect 283426 -1862 283662 -1626
rect 283746 -1862 283982 -1626
rect 282026 -2502 282262 -2266
rect 282346 -2502 282582 -2266
rect 282026 -2822 282262 -2586
rect 282346 -2822 282582 -2586
rect 280626 -5382 280862 -5146
rect 280946 -5382 281182 -5146
rect 280626 -5702 280862 -5466
rect 280946 -5702 281182 -5466
rect 279226 -6342 279462 -6106
rect 279546 -6342 279782 -6106
rect 279226 -6662 279462 -6426
rect 279546 -6662 279782 -6426
rect 285746 10658 285982 10894
rect 286066 10658 286302 10894
rect 285746 10338 285982 10574
rect 286066 10338 286302 10574
rect 288546 3218 288782 3454
rect 288866 3218 289102 3454
rect 288546 2898 288782 3134
rect 288866 2898 289102 3134
rect 288546 -582 288782 -346
rect 288866 -582 289102 -346
rect 288546 -902 288782 -666
rect 288866 -902 289102 -666
rect 287146 -3462 287382 -3226
rect 287466 -3462 287702 -3226
rect 287146 -3782 287382 -3546
rect 287466 -3782 287702 -3546
rect 285746 -4422 285982 -4186
rect 286066 -4422 286302 -4186
rect 285746 -4742 285982 -4506
rect 286066 -4742 286302 -4506
rect 284346 -7302 284582 -7066
rect 284666 -7302 284902 -7066
rect 284346 -7622 284582 -7386
rect 284666 -7622 284902 -7386
rect 292266 6938 292502 7174
rect 292586 6938 292822 7174
rect 292266 6618 292502 6854
rect 292586 6618 292822 6854
rect 293666 -1542 293902 -1306
rect 293986 -1542 294222 -1306
rect 293666 -1862 293902 -1626
rect 293986 -1862 294222 -1626
rect 292266 -2502 292502 -2266
rect 292586 -2502 292822 -2266
rect 292266 -2822 292502 -2586
rect 292586 -2822 292822 -2586
rect 290866 -5382 291102 -5146
rect 291186 -5382 291422 -5146
rect 290866 -5702 291102 -5466
rect 291186 -5702 291422 -5466
rect 289466 -6342 289702 -6106
rect 289786 -6342 290022 -6106
rect 289466 -6662 289702 -6426
rect 289786 -6662 290022 -6426
rect 295986 10658 296222 10894
rect 296306 10658 296542 10894
rect 295986 10338 296222 10574
rect 296306 10338 296542 10574
rect 298786 3218 299022 3454
rect 299106 3218 299342 3454
rect 298786 2898 299022 3134
rect 299106 2898 299342 3134
rect 298786 -582 299022 -346
rect 299106 -582 299342 -346
rect 298786 -902 299022 -666
rect 299106 -902 299342 -666
rect 297386 -3462 297622 -3226
rect 297706 -3462 297942 -3226
rect 297386 -3782 297622 -3546
rect 297706 -3782 297942 -3546
rect 295986 -4422 296222 -4186
rect 296306 -4422 296542 -4186
rect 295986 -4742 296222 -4506
rect 296306 -4742 296542 -4506
rect 294586 -7302 294822 -7066
rect 294906 -7302 295142 -7066
rect 294586 -7622 294822 -7386
rect 294906 -7622 295142 -7386
rect 302506 6938 302742 7174
rect 302826 6938 303062 7174
rect 302506 6618 302742 6854
rect 302826 6618 303062 6854
rect 303906 -1542 304142 -1306
rect 304226 -1542 304462 -1306
rect 303906 -1862 304142 -1626
rect 304226 -1862 304462 -1626
rect 302506 -2502 302742 -2266
rect 302826 -2502 303062 -2266
rect 302506 -2822 302742 -2586
rect 302826 -2822 303062 -2586
rect 301106 -5382 301342 -5146
rect 301426 -5382 301662 -5146
rect 301106 -5702 301342 -5466
rect 301426 -5702 301662 -5466
rect 299706 -6342 299942 -6106
rect 300026 -6342 300262 -6106
rect 299706 -6662 299942 -6426
rect 300026 -6662 300262 -6426
rect 306226 10658 306462 10894
rect 306546 10658 306782 10894
rect 306226 10338 306462 10574
rect 306546 10338 306782 10574
rect 309026 3218 309262 3454
rect 309346 3218 309582 3454
rect 309026 2898 309262 3134
rect 309346 2898 309582 3134
rect 309026 -582 309262 -346
rect 309346 -582 309582 -346
rect 309026 -902 309262 -666
rect 309346 -902 309582 -666
rect 307626 -3462 307862 -3226
rect 307946 -3462 308182 -3226
rect 307626 -3782 307862 -3546
rect 307946 -3782 308182 -3546
rect 306226 -4422 306462 -4186
rect 306546 -4422 306782 -4186
rect 306226 -4742 306462 -4506
rect 306546 -4742 306782 -4506
rect 304826 -7302 305062 -7066
rect 305146 -7302 305382 -7066
rect 304826 -7622 305062 -7386
rect 305146 -7622 305382 -7386
rect 312746 6938 312982 7174
rect 313066 6938 313302 7174
rect 312746 6618 312982 6854
rect 313066 6618 313302 6854
rect 314146 -1542 314382 -1306
rect 314466 -1542 314702 -1306
rect 314146 -1862 314382 -1626
rect 314466 -1862 314702 -1626
rect 312746 -2502 312982 -2266
rect 313066 -2502 313302 -2266
rect 312746 -2822 312982 -2586
rect 313066 -2822 313302 -2586
rect 311346 -5382 311582 -5146
rect 311666 -5382 311902 -5146
rect 311346 -5702 311582 -5466
rect 311666 -5702 311902 -5466
rect 309946 -6342 310182 -6106
rect 310266 -6342 310502 -6106
rect 309946 -6662 310182 -6426
rect 310266 -6662 310502 -6426
rect 316466 10658 316702 10894
rect 316786 10658 317022 10894
rect 316466 10338 316702 10574
rect 316786 10338 317022 10574
rect 319266 3218 319502 3454
rect 319586 3218 319822 3454
rect 319266 2898 319502 3134
rect 319586 2898 319822 3134
rect 319266 -582 319502 -346
rect 319586 -582 319822 -346
rect 319266 -902 319502 -666
rect 319586 -902 319822 -666
rect 317866 -3462 318102 -3226
rect 318186 -3462 318422 -3226
rect 317866 -3782 318102 -3546
rect 318186 -3782 318422 -3546
rect 316466 -4422 316702 -4186
rect 316786 -4422 317022 -4186
rect 316466 -4742 316702 -4506
rect 316786 -4742 317022 -4506
rect 315066 -7302 315302 -7066
rect 315386 -7302 315622 -7066
rect 315066 -7622 315302 -7386
rect 315386 -7622 315622 -7386
rect 322986 6938 323222 7174
rect 323306 6938 323542 7174
rect 322986 6618 323222 6854
rect 323306 6618 323542 6854
rect 324386 -1542 324622 -1306
rect 324706 -1542 324942 -1306
rect 324386 -1862 324622 -1626
rect 324706 -1862 324942 -1626
rect 322986 -2502 323222 -2266
rect 323306 -2502 323542 -2266
rect 322986 -2822 323222 -2586
rect 323306 -2822 323542 -2586
rect 321586 -5382 321822 -5146
rect 321906 -5382 322142 -5146
rect 321586 -5702 321822 -5466
rect 321906 -5702 322142 -5466
rect 320186 -6342 320422 -6106
rect 320506 -6342 320742 -6106
rect 320186 -6662 320422 -6426
rect 320506 -6662 320742 -6426
rect 326706 10658 326942 10894
rect 327026 10658 327262 10894
rect 326706 10338 326942 10574
rect 327026 10338 327262 10574
rect 329506 3218 329742 3454
rect 329826 3218 330062 3454
rect 329506 2898 329742 3134
rect 329826 2898 330062 3134
rect 329506 -582 329742 -346
rect 329826 -582 330062 -346
rect 329506 -902 329742 -666
rect 329826 -902 330062 -666
rect 328106 -3462 328342 -3226
rect 328426 -3462 328662 -3226
rect 328106 -3782 328342 -3546
rect 328426 -3782 328662 -3546
rect 326706 -4422 326942 -4186
rect 327026 -4422 327262 -4186
rect 326706 -4742 326942 -4506
rect 327026 -4742 327262 -4506
rect 325306 -7302 325542 -7066
rect 325626 -7302 325862 -7066
rect 325306 -7622 325542 -7386
rect 325626 -7622 325862 -7386
rect 333226 6938 333462 7174
rect 333546 6938 333782 7174
rect 333226 6618 333462 6854
rect 333546 6618 333782 6854
rect 334626 -1542 334862 -1306
rect 334946 -1542 335182 -1306
rect 334626 -1862 334862 -1626
rect 334946 -1862 335182 -1626
rect 333226 -2502 333462 -2266
rect 333546 -2502 333782 -2266
rect 333226 -2822 333462 -2586
rect 333546 -2822 333782 -2586
rect 331826 -5382 332062 -5146
rect 332146 -5382 332382 -5146
rect 331826 -5702 332062 -5466
rect 332146 -5702 332382 -5466
rect 330426 -6342 330662 -6106
rect 330746 -6342 330982 -6106
rect 330426 -6662 330662 -6426
rect 330746 -6662 330982 -6426
rect 336946 10658 337182 10894
rect 337266 10658 337502 10894
rect 336946 10338 337182 10574
rect 337266 10338 337502 10574
rect 339746 3218 339982 3454
rect 340066 3218 340302 3454
rect 339746 2898 339982 3134
rect 340066 2898 340302 3134
rect 339746 -582 339982 -346
rect 340066 -582 340302 -346
rect 339746 -902 339982 -666
rect 340066 -902 340302 -666
rect 338346 -3462 338582 -3226
rect 338666 -3462 338902 -3226
rect 338346 -3782 338582 -3546
rect 338666 -3782 338902 -3546
rect 336946 -4422 337182 -4186
rect 337266 -4422 337502 -4186
rect 336946 -4742 337182 -4506
rect 337266 -4742 337502 -4506
rect 335546 -7302 335782 -7066
rect 335866 -7302 336102 -7066
rect 335546 -7622 335782 -7386
rect 335866 -7622 336102 -7386
rect 343466 6938 343702 7174
rect 343786 6938 344022 7174
rect 343466 6618 343702 6854
rect 343786 6618 344022 6854
rect 344866 -1542 345102 -1306
rect 345186 -1542 345422 -1306
rect 344866 -1862 345102 -1626
rect 345186 -1862 345422 -1626
rect 343466 -2502 343702 -2266
rect 343786 -2502 344022 -2266
rect 343466 -2822 343702 -2586
rect 343786 -2822 344022 -2586
rect 342066 -5382 342302 -5146
rect 342386 -5382 342622 -5146
rect 342066 -5702 342302 -5466
rect 342386 -5702 342622 -5466
rect 340666 -6342 340902 -6106
rect 340986 -6342 341222 -6106
rect 340666 -6662 340902 -6426
rect 340986 -6662 341222 -6426
rect 347186 10658 347422 10894
rect 347506 10658 347742 10894
rect 347186 10338 347422 10574
rect 347506 10338 347742 10574
rect 349986 3218 350222 3454
rect 350306 3218 350542 3454
rect 349986 2898 350222 3134
rect 350306 2898 350542 3134
rect 349986 -582 350222 -346
rect 350306 -582 350542 -346
rect 349986 -902 350222 -666
rect 350306 -902 350542 -666
rect 348586 -3462 348822 -3226
rect 348906 -3462 349142 -3226
rect 348586 -3782 348822 -3546
rect 348906 -3782 349142 -3546
rect 347186 -4422 347422 -4186
rect 347506 -4422 347742 -4186
rect 347186 -4742 347422 -4506
rect 347506 -4742 347742 -4506
rect 345786 -7302 346022 -7066
rect 346106 -7302 346342 -7066
rect 345786 -7622 346022 -7386
rect 346106 -7622 346342 -7386
rect 353706 6938 353942 7174
rect 354026 6938 354262 7174
rect 353706 6618 353942 6854
rect 354026 6618 354262 6854
rect 355106 -1542 355342 -1306
rect 355426 -1542 355662 -1306
rect 355106 -1862 355342 -1626
rect 355426 -1862 355662 -1626
rect 353706 -2502 353942 -2266
rect 354026 -2502 354262 -2266
rect 353706 -2822 353942 -2586
rect 354026 -2822 354262 -2586
rect 352306 -5382 352542 -5146
rect 352626 -5382 352862 -5146
rect 352306 -5702 352542 -5466
rect 352626 -5702 352862 -5466
rect 350906 -6342 351142 -6106
rect 351226 -6342 351462 -6106
rect 350906 -6662 351142 -6426
rect 351226 -6662 351462 -6426
rect 357426 10658 357662 10894
rect 357746 10658 357982 10894
rect 357426 10338 357662 10574
rect 357746 10338 357982 10574
rect 360226 3218 360462 3454
rect 360546 3218 360782 3454
rect 360226 2898 360462 3134
rect 360546 2898 360782 3134
rect 360226 -582 360462 -346
rect 360546 -582 360782 -346
rect 360226 -902 360462 -666
rect 360546 -902 360782 -666
rect 358826 -3462 359062 -3226
rect 359146 -3462 359382 -3226
rect 358826 -3782 359062 -3546
rect 359146 -3782 359382 -3546
rect 357426 -4422 357662 -4186
rect 357746 -4422 357982 -4186
rect 357426 -4742 357662 -4506
rect 357746 -4742 357982 -4506
rect 356026 -7302 356262 -7066
rect 356346 -7302 356582 -7066
rect 356026 -7622 356262 -7386
rect 356346 -7622 356582 -7386
rect 363946 6938 364182 7174
rect 364266 6938 364502 7174
rect 363946 6618 364182 6854
rect 364266 6618 364502 6854
rect 365346 -1542 365582 -1306
rect 365666 -1542 365902 -1306
rect 365346 -1862 365582 -1626
rect 365666 -1862 365902 -1626
rect 363946 -2502 364182 -2266
rect 364266 -2502 364502 -2266
rect 363946 -2822 364182 -2586
rect 364266 -2822 364502 -2586
rect 362546 -5382 362782 -5146
rect 362866 -5382 363102 -5146
rect 362546 -5702 362782 -5466
rect 362866 -5702 363102 -5466
rect 361146 -6342 361382 -6106
rect 361466 -6342 361702 -6106
rect 361146 -6662 361382 -6426
rect 361466 -6662 361702 -6426
rect 367666 10658 367902 10894
rect 367986 10658 368222 10894
rect 367666 10338 367902 10574
rect 367986 10338 368222 10574
rect 370466 3218 370702 3454
rect 370786 3218 371022 3454
rect 370466 2898 370702 3134
rect 370786 2898 371022 3134
rect 370466 -582 370702 -346
rect 370786 -582 371022 -346
rect 370466 -902 370702 -666
rect 370786 -902 371022 -666
rect 369066 -3462 369302 -3226
rect 369386 -3462 369622 -3226
rect 369066 -3782 369302 -3546
rect 369386 -3782 369622 -3546
rect 367666 -4422 367902 -4186
rect 367986 -4422 368222 -4186
rect 367666 -4742 367902 -4506
rect 367986 -4742 368222 -4506
rect 366266 -7302 366502 -7066
rect 366586 -7302 366822 -7066
rect 366266 -7622 366502 -7386
rect 366586 -7622 366822 -7386
rect 374186 6938 374422 7174
rect 374506 6938 374742 7174
rect 374186 6618 374422 6854
rect 374506 6618 374742 6854
rect 375586 -1542 375822 -1306
rect 375906 -1542 376142 -1306
rect 375586 -1862 375822 -1626
rect 375906 -1862 376142 -1626
rect 374186 -2502 374422 -2266
rect 374506 -2502 374742 -2266
rect 374186 -2822 374422 -2586
rect 374506 -2822 374742 -2586
rect 372786 -5382 373022 -5146
rect 373106 -5382 373342 -5146
rect 372786 -5702 373022 -5466
rect 373106 -5702 373342 -5466
rect 371386 -6342 371622 -6106
rect 371706 -6342 371942 -6106
rect 371386 -6662 371622 -6426
rect 371706 -6662 371942 -6426
rect 377906 10658 378142 10894
rect 378226 10658 378462 10894
rect 377906 10338 378142 10574
rect 378226 10338 378462 10574
rect 380706 3218 380942 3454
rect 381026 3218 381262 3454
rect 380706 2898 380942 3134
rect 381026 2898 381262 3134
rect 380706 -582 380942 -346
rect 381026 -582 381262 -346
rect 380706 -902 380942 -666
rect 381026 -902 381262 -666
rect 379306 -3462 379542 -3226
rect 379626 -3462 379862 -3226
rect 379306 -3782 379542 -3546
rect 379626 -3782 379862 -3546
rect 377906 -4422 378142 -4186
rect 378226 -4422 378462 -4186
rect 377906 -4742 378142 -4506
rect 378226 -4742 378462 -4506
rect 376506 -7302 376742 -7066
rect 376826 -7302 377062 -7066
rect 376506 -7622 376742 -7386
rect 376826 -7622 377062 -7386
rect 384426 6938 384662 7174
rect 384746 6938 384982 7174
rect 384426 6618 384662 6854
rect 384746 6618 384982 6854
rect 385826 -1542 386062 -1306
rect 386146 -1542 386382 -1306
rect 385826 -1862 386062 -1626
rect 386146 -1862 386382 -1626
rect 384426 -2502 384662 -2266
rect 384746 -2502 384982 -2266
rect 384426 -2822 384662 -2586
rect 384746 -2822 384982 -2586
rect 383026 -5382 383262 -5146
rect 383346 -5382 383582 -5146
rect 383026 -5702 383262 -5466
rect 383346 -5702 383582 -5466
rect 381626 -6342 381862 -6106
rect 381946 -6342 382182 -6106
rect 381626 -6662 381862 -6426
rect 381946 -6662 382182 -6426
rect 388146 10658 388382 10894
rect 388466 10658 388702 10894
rect 388146 10338 388382 10574
rect 388466 10338 388702 10574
rect 390946 3218 391182 3454
rect 391266 3218 391502 3454
rect 390946 2898 391182 3134
rect 391266 2898 391502 3134
rect 390946 -582 391182 -346
rect 391266 -582 391502 -346
rect 390946 -902 391182 -666
rect 391266 -902 391502 -666
rect 389546 -3462 389782 -3226
rect 389866 -3462 390102 -3226
rect 389546 -3782 389782 -3546
rect 389866 -3782 390102 -3546
rect 388146 -4422 388382 -4186
rect 388466 -4422 388702 -4186
rect 388146 -4742 388382 -4506
rect 388466 -4742 388702 -4506
rect 386746 -7302 386982 -7066
rect 387066 -7302 387302 -7066
rect 386746 -7622 386982 -7386
rect 387066 -7622 387302 -7386
rect 394666 6938 394902 7174
rect 394986 6938 395222 7174
rect 394666 6618 394902 6854
rect 394986 6618 395222 6854
rect 396066 -1542 396302 -1306
rect 396386 -1542 396622 -1306
rect 396066 -1862 396302 -1626
rect 396386 -1862 396622 -1626
rect 394666 -2502 394902 -2266
rect 394986 -2502 395222 -2266
rect 394666 -2822 394902 -2586
rect 394986 -2822 395222 -2586
rect 393266 -5382 393502 -5146
rect 393586 -5382 393822 -5146
rect 393266 -5702 393502 -5466
rect 393586 -5702 393822 -5466
rect 391866 -6342 392102 -6106
rect 392186 -6342 392422 -6106
rect 391866 -6662 392102 -6426
rect 392186 -6662 392422 -6426
rect 398386 10658 398622 10894
rect 398706 10658 398942 10894
rect 398386 10338 398622 10574
rect 398706 10338 398942 10574
rect 401186 3218 401422 3454
rect 401506 3218 401742 3454
rect 401186 2898 401422 3134
rect 401506 2898 401742 3134
rect 401186 -582 401422 -346
rect 401506 -582 401742 -346
rect 401186 -902 401422 -666
rect 401506 -902 401742 -666
rect 399786 -3462 400022 -3226
rect 400106 -3462 400342 -3226
rect 399786 -3782 400022 -3546
rect 400106 -3782 400342 -3546
rect 398386 -4422 398622 -4186
rect 398706 -4422 398942 -4186
rect 398386 -4742 398622 -4506
rect 398706 -4742 398942 -4506
rect 396986 -7302 397222 -7066
rect 397306 -7302 397542 -7066
rect 396986 -7622 397222 -7386
rect 397306 -7622 397542 -7386
rect 404906 6938 405142 7174
rect 405226 6938 405462 7174
rect 404906 6618 405142 6854
rect 405226 6618 405462 6854
rect 406306 -1542 406542 -1306
rect 406626 -1542 406862 -1306
rect 406306 -1862 406542 -1626
rect 406626 -1862 406862 -1626
rect 404906 -2502 405142 -2266
rect 405226 -2502 405462 -2266
rect 404906 -2822 405142 -2586
rect 405226 -2822 405462 -2586
rect 403506 -5382 403742 -5146
rect 403826 -5382 404062 -5146
rect 403506 -5702 403742 -5466
rect 403826 -5702 404062 -5466
rect 402106 -6342 402342 -6106
rect 402426 -6342 402662 -6106
rect 402106 -6662 402342 -6426
rect 402426 -6662 402662 -6426
rect 408626 10658 408862 10894
rect 408946 10658 409182 10894
rect 408626 10338 408862 10574
rect 408946 10338 409182 10574
rect 411426 3218 411662 3454
rect 411746 3218 411982 3454
rect 411426 2898 411662 3134
rect 411746 2898 411982 3134
rect 411426 -582 411662 -346
rect 411746 -582 411982 -346
rect 411426 -902 411662 -666
rect 411746 -902 411982 -666
rect 410026 -3462 410262 -3226
rect 410346 -3462 410582 -3226
rect 410026 -3782 410262 -3546
rect 410346 -3782 410582 -3546
rect 408626 -4422 408862 -4186
rect 408946 -4422 409182 -4186
rect 408626 -4742 408862 -4506
rect 408946 -4742 409182 -4506
rect 407226 -7302 407462 -7066
rect 407546 -7302 407782 -7066
rect 407226 -7622 407462 -7386
rect 407546 -7622 407782 -7386
rect 415146 6938 415382 7174
rect 415466 6938 415702 7174
rect 415146 6618 415382 6854
rect 415466 6618 415702 6854
rect 416546 -1542 416782 -1306
rect 416866 -1542 417102 -1306
rect 416546 -1862 416782 -1626
rect 416866 -1862 417102 -1626
rect 415146 -2502 415382 -2266
rect 415466 -2502 415702 -2266
rect 415146 -2822 415382 -2586
rect 415466 -2822 415702 -2586
rect 413746 -5382 413982 -5146
rect 414066 -5382 414302 -5146
rect 413746 -5702 413982 -5466
rect 414066 -5702 414302 -5466
rect 412346 -6342 412582 -6106
rect 412666 -6342 412902 -6106
rect 412346 -6662 412582 -6426
rect 412666 -6662 412902 -6426
rect 418866 10658 419102 10894
rect 419186 10658 419422 10894
rect 418866 10338 419102 10574
rect 419186 10338 419422 10574
rect 421666 3218 421902 3454
rect 421986 3218 422222 3454
rect 421666 2898 421902 3134
rect 421986 2898 422222 3134
rect 421666 -582 421902 -346
rect 421986 -582 422222 -346
rect 421666 -902 421902 -666
rect 421986 -902 422222 -666
rect 420266 -3462 420502 -3226
rect 420586 -3462 420822 -3226
rect 420266 -3782 420502 -3546
rect 420586 -3782 420822 -3546
rect 418866 -4422 419102 -4186
rect 419186 -4422 419422 -4186
rect 418866 -4742 419102 -4506
rect 419186 -4742 419422 -4506
rect 417466 -7302 417702 -7066
rect 417786 -7302 418022 -7066
rect 417466 -7622 417702 -7386
rect 417786 -7622 418022 -7386
rect 425386 6938 425622 7174
rect 425706 6938 425942 7174
rect 425386 6618 425622 6854
rect 425706 6618 425942 6854
rect 426786 -1542 427022 -1306
rect 427106 -1542 427342 -1306
rect 426786 -1862 427022 -1626
rect 427106 -1862 427342 -1626
rect 425386 -2502 425622 -2266
rect 425706 -2502 425942 -2266
rect 425386 -2822 425622 -2586
rect 425706 -2822 425942 -2586
rect 423986 -5382 424222 -5146
rect 424306 -5382 424542 -5146
rect 423986 -5702 424222 -5466
rect 424306 -5702 424542 -5466
rect 422586 -6342 422822 -6106
rect 422906 -6342 423142 -6106
rect 422586 -6662 422822 -6426
rect 422906 -6662 423142 -6426
rect 429106 10658 429342 10894
rect 429426 10658 429662 10894
rect 429106 10338 429342 10574
rect 429426 10338 429662 10574
rect 431906 3218 432142 3454
rect 432226 3218 432462 3454
rect 431906 2898 432142 3134
rect 432226 2898 432462 3134
rect 431906 -582 432142 -346
rect 432226 -582 432462 -346
rect 431906 -902 432142 -666
rect 432226 -902 432462 -666
rect 430506 -3462 430742 -3226
rect 430826 -3462 431062 -3226
rect 430506 -3782 430742 -3546
rect 430826 -3782 431062 -3546
rect 429106 -4422 429342 -4186
rect 429426 -4422 429662 -4186
rect 429106 -4742 429342 -4506
rect 429426 -4742 429662 -4506
rect 427706 -7302 427942 -7066
rect 428026 -7302 428262 -7066
rect 427706 -7622 427942 -7386
rect 428026 -7622 428262 -7386
rect 435626 6938 435862 7174
rect 435946 6938 436182 7174
rect 435626 6618 435862 6854
rect 435946 6618 436182 6854
rect 437026 -1542 437262 -1306
rect 437346 -1542 437582 -1306
rect 437026 -1862 437262 -1626
rect 437346 -1862 437582 -1626
rect 435626 -2502 435862 -2266
rect 435946 -2502 436182 -2266
rect 435626 -2822 435862 -2586
rect 435946 -2822 436182 -2586
rect 434226 -5382 434462 -5146
rect 434546 -5382 434782 -5146
rect 434226 -5702 434462 -5466
rect 434546 -5702 434782 -5466
rect 432826 -6342 433062 -6106
rect 433146 -6342 433382 -6106
rect 432826 -6662 433062 -6426
rect 433146 -6662 433382 -6426
rect 439346 10658 439582 10894
rect 439666 10658 439902 10894
rect 439346 10338 439582 10574
rect 439666 10338 439902 10574
rect 442146 3218 442382 3454
rect 442466 3218 442702 3454
rect 442146 2898 442382 3134
rect 442466 2898 442702 3134
rect 442146 -582 442382 -346
rect 442466 -582 442702 -346
rect 442146 -902 442382 -666
rect 442466 -902 442702 -666
rect 440746 -3462 440982 -3226
rect 441066 -3462 441302 -3226
rect 440746 -3782 440982 -3546
rect 441066 -3782 441302 -3546
rect 439346 -4422 439582 -4186
rect 439666 -4422 439902 -4186
rect 439346 -4742 439582 -4506
rect 439666 -4742 439902 -4506
rect 437946 -7302 438182 -7066
rect 438266 -7302 438502 -7066
rect 437946 -7622 438182 -7386
rect 438266 -7622 438502 -7386
rect 445866 6938 446102 7174
rect 446186 6938 446422 7174
rect 445866 6618 446102 6854
rect 446186 6618 446422 6854
rect 447266 -1542 447502 -1306
rect 447586 -1542 447822 -1306
rect 447266 -1862 447502 -1626
rect 447586 -1862 447822 -1626
rect 445866 -2502 446102 -2266
rect 446186 -2502 446422 -2266
rect 445866 -2822 446102 -2586
rect 446186 -2822 446422 -2586
rect 444466 -5382 444702 -5146
rect 444786 -5382 445022 -5146
rect 444466 -5702 444702 -5466
rect 444786 -5702 445022 -5466
rect 443066 -6342 443302 -6106
rect 443386 -6342 443622 -6106
rect 443066 -6662 443302 -6426
rect 443386 -6662 443622 -6426
rect 449586 10658 449822 10894
rect 449906 10658 450142 10894
rect 449586 10338 449822 10574
rect 449906 10338 450142 10574
rect 452386 3218 452622 3454
rect 452706 3218 452942 3454
rect 452386 2898 452622 3134
rect 452706 2898 452942 3134
rect 452386 -582 452622 -346
rect 452706 -582 452942 -346
rect 452386 -902 452622 -666
rect 452706 -902 452942 -666
rect 450986 -3462 451222 -3226
rect 451306 -3462 451542 -3226
rect 450986 -3782 451222 -3546
rect 451306 -3782 451542 -3546
rect 449586 -4422 449822 -4186
rect 449906 -4422 450142 -4186
rect 449586 -4742 449822 -4506
rect 449906 -4742 450142 -4506
rect 448186 -7302 448422 -7066
rect 448506 -7302 448742 -7066
rect 448186 -7622 448422 -7386
rect 448506 -7622 448742 -7386
rect 456106 6938 456342 7174
rect 456426 6938 456662 7174
rect 456106 6618 456342 6854
rect 456426 6618 456662 6854
rect 457506 -1542 457742 -1306
rect 457826 -1542 458062 -1306
rect 457506 -1862 457742 -1626
rect 457826 -1862 458062 -1626
rect 456106 -2502 456342 -2266
rect 456426 -2502 456662 -2266
rect 456106 -2822 456342 -2586
rect 456426 -2822 456662 -2586
rect 454706 -5382 454942 -5146
rect 455026 -5382 455262 -5146
rect 454706 -5702 454942 -5466
rect 455026 -5702 455262 -5466
rect 453306 -6342 453542 -6106
rect 453626 -6342 453862 -6106
rect 453306 -6662 453542 -6426
rect 453626 -6662 453862 -6426
rect 459826 10658 460062 10894
rect 460146 10658 460382 10894
rect 459826 10338 460062 10574
rect 460146 10338 460382 10574
rect 462626 3218 462862 3454
rect 462946 3218 463182 3454
rect 462626 2898 462862 3134
rect 462946 2898 463182 3134
rect 462626 -582 462862 -346
rect 462946 -582 463182 -346
rect 462626 -902 462862 -666
rect 462946 -902 463182 -666
rect 461226 -3462 461462 -3226
rect 461546 -3462 461782 -3226
rect 461226 -3782 461462 -3546
rect 461546 -3782 461782 -3546
rect 459826 -4422 460062 -4186
rect 460146 -4422 460382 -4186
rect 459826 -4742 460062 -4506
rect 460146 -4742 460382 -4506
rect 458426 -7302 458662 -7066
rect 458746 -7302 458982 -7066
rect 458426 -7622 458662 -7386
rect 458746 -7622 458982 -7386
rect 466346 6938 466582 7174
rect 466666 6938 466902 7174
rect 466346 6618 466582 6854
rect 466666 6618 466902 6854
rect 467746 -1542 467982 -1306
rect 468066 -1542 468302 -1306
rect 467746 -1862 467982 -1626
rect 468066 -1862 468302 -1626
rect 466346 -2502 466582 -2266
rect 466666 -2502 466902 -2266
rect 466346 -2822 466582 -2586
rect 466666 -2822 466902 -2586
rect 464946 -5382 465182 -5146
rect 465266 -5382 465502 -5146
rect 464946 -5702 465182 -5466
rect 465266 -5702 465502 -5466
rect 463546 -6342 463782 -6106
rect 463866 -6342 464102 -6106
rect 463546 -6662 463782 -6426
rect 463866 -6662 464102 -6426
rect 470066 10658 470302 10894
rect 470386 10658 470622 10894
rect 470066 10338 470302 10574
rect 470386 10338 470622 10574
rect 472866 3218 473102 3454
rect 473186 3218 473422 3454
rect 472866 2898 473102 3134
rect 473186 2898 473422 3134
rect 472866 -582 473102 -346
rect 473186 -582 473422 -346
rect 472866 -902 473102 -666
rect 473186 -902 473422 -666
rect 471466 -3462 471702 -3226
rect 471786 -3462 472022 -3226
rect 471466 -3782 471702 -3546
rect 471786 -3782 472022 -3546
rect 470066 -4422 470302 -4186
rect 470386 -4422 470622 -4186
rect 470066 -4742 470302 -4506
rect 470386 -4742 470622 -4506
rect 468666 -7302 468902 -7066
rect 468986 -7302 469222 -7066
rect 468666 -7622 468902 -7386
rect 468986 -7622 469222 -7386
rect 476586 6938 476822 7174
rect 476906 6938 477142 7174
rect 476586 6618 476822 6854
rect 476906 6618 477142 6854
rect 477986 -1542 478222 -1306
rect 478306 -1542 478542 -1306
rect 477986 -1862 478222 -1626
rect 478306 -1862 478542 -1626
rect 476586 -2502 476822 -2266
rect 476906 -2502 477142 -2266
rect 476586 -2822 476822 -2586
rect 476906 -2822 477142 -2586
rect 475186 -5382 475422 -5146
rect 475506 -5382 475742 -5146
rect 475186 -5702 475422 -5466
rect 475506 -5702 475742 -5466
rect 473786 -6342 474022 -6106
rect 474106 -6342 474342 -6106
rect 473786 -6662 474022 -6426
rect 474106 -6662 474342 -6426
rect 480306 10658 480542 10894
rect 480626 10658 480862 10894
rect 480306 10338 480542 10574
rect 480626 10338 480862 10574
rect 483106 3218 483342 3454
rect 483426 3218 483662 3454
rect 483106 2898 483342 3134
rect 483426 2898 483662 3134
rect 483106 -582 483342 -346
rect 483426 -582 483662 -346
rect 483106 -902 483342 -666
rect 483426 -902 483662 -666
rect 481706 -3462 481942 -3226
rect 482026 -3462 482262 -3226
rect 481706 -3782 481942 -3546
rect 482026 -3782 482262 -3546
rect 480306 -4422 480542 -4186
rect 480626 -4422 480862 -4186
rect 480306 -4742 480542 -4506
rect 480626 -4742 480862 -4506
rect 478906 -7302 479142 -7066
rect 479226 -7302 479462 -7066
rect 478906 -7622 479142 -7386
rect 479226 -7622 479462 -7386
rect 486826 6938 487062 7174
rect 487146 6938 487382 7174
rect 486826 6618 487062 6854
rect 487146 6618 487382 6854
rect 488226 -1542 488462 -1306
rect 488546 -1542 488782 -1306
rect 488226 -1862 488462 -1626
rect 488546 -1862 488782 -1626
rect 486826 -2502 487062 -2266
rect 487146 -2502 487382 -2266
rect 486826 -2822 487062 -2586
rect 487146 -2822 487382 -2586
rect 485426 -5382 485662 -5146
rect 485746 -5382 485982 -5146
rect 485426 -5702 485662 -5466
rect 485746 -5702 485982 -5466
rect 484026 -6342 484262 -6106
rect 484346 -6342 484582 -6106
rect 484026 -6662 484262 -6426
rect 484346 -6662 484582 -6426
rect 490546 10658 490782 10894
rect 490866 10658 491102 10894
rect 490546 10338 490782 10574
rect 490866 10338 491102 10574
rect 493346 3218 493582 3454
rect 493666 3218 493902 3454
rect 493346 2898 493582 3134
rect 493666 2898 493902 3134
rect 493346 -582 493582 -346
rect 493666 -582 493902 -346
rect 493346 -902 493582 -666
rect 493666 -902 493902 -666
rect 491946 -3462 492182 -3226
rect 492266 -3462 492502 -3226
rect 491946 -3782 492182 -3546
rect 492266 -3782 492502 -3546
rect 490546 -4422 490782 -4186
rect 490866 -4422 491102 -4186
rect 490546 -4742 490782 -4506
rect 490866 -4742 491102 -4506
rect 489146 -7302 489382 -7066
rect 489466 -7302 489702 -7066
rect 489146 -7622 489382 -7386
rect 489466 -7622 489702 -7386
rect 497066 6938 497302 7174
rect 497386 6938 497622 7174
rect 497066 6618 497302 6854
rect 497386 6618 497622 6854
rect 498466 -1542 498702 -1306
rect 498786 -1542 499022 -1306
rect 498466 -1862 498702 -1626
rect 498786 -1862 499022 -1626
rect 497066 -2502 497302 -2266
rect 497386 -2502 497622 -2266
rect 497066 -2822 497302 -2586
rect 497386 -2822 497622 -2586
rect 495666 -5382 495902 -5146
rect 495986 -5382 496222 -5146
rect 495666 -5702 495902 -5466
rect 495986 -5702 496222 -5466
rect 494266 -6342 494502 -6106
rect 494586 -6342 494822 -6106
rect 494266 -6662 494502 -6426
rect 494586 -6662 494822 -6426
rect 500786 10658 501022 10894
rect 501106 10658 501342 10894
rect 500786 10338 501022 10574
rect 501106 10338 501342 10574
rect 503586 3218 503822 3454
rect 503906 3218 504142 3454
rect 503586 2898 503822 3134
rect 503906 2898 504142 3134
rect 503586 -582 503822 -346
rect 503906 -582 504142 -346
rect 503586 -902 503822 -666
rect 503906 -902 504142 -666
rect 502186 -3462 502422 -3226
rect 502506 -3462 502742 -3226
rect 502186 -3782 502422 -3546
rect 502506 -3782 502742 -3546
rect 500786 -4422 501022 -4186
rect 501106 -4422 501342 -4186
rect 500786 -4742 501022 -4506
rect 501106 -4742 501342 -4506
rect 499386 -7302 499622 -7066
rect 499706 -7302 499942 -7066
rect 499386 -7622 499622 -7386
rect 499706 -7622 499942 -7386
rect 507306 6938 507542 7174
rect 507626 6938 507862 7174
rect 507306 6618 507542 6854
rect 507626 6618 507862 6854
rect 508706 -1542 508942 -1306
rect 509026 -1542 509262 -1306
rect 508706 -1862 508942 -1626
rect 509026 -1862 509262 -1626
rect 507306 -2502 507542 -2266
rect 507626 -2502 507862 -2266
rect 507306 -2822 507542 -2586
rect 507626 -2822 507862 -2586
rect 505906 -5382 506142 -5146
rect 506226 -5382 506462 -5146
rect 505906 -5702 506142 -5466
rect 506226 -5702 506462 -5466
rect 504506 -6342 504742 -6106
rect 504826 -6342 505062 -6106
rect 504506 -6662 504742 -6426
rect 504826 -6662 505062 -6426
rect 511026 10658 511262 10894
rect 511346 10658 511582 10894
rect 511026 10338 511262 10574
rect 511346 10338 511582 10574
rect 513826 3218 514062 3454
rect 514146 3218 514382 3454
rect 513826 2898 514062 3134
rect 514146 2898 514382 3134
rect 513826 -582 514062 -346
rect 514146 -582 514382 -346
rect 513826 -902 514062 -666
rect 514146 -902 514382 -666
rect 512426 -3462 512662 -3226
rect 512746 -3462 512982 -3226
rect 512426 -3782 512662 -3546
rect 512746 -3782 512982 -3546
rect 511026 -4422 511262 -4186
rect 511346 -4422 511582 -4186
rect 511026 -4742 511262 -4506
rect 511346 -4742 511582 -4506
rect 509626 -7302 509862 -7066
rect 509946 -7302 510182 -7066
rect 509626 -7622 509862 -7386
rect 509946 -7622 510182 -7386
rect 517546 6938 517782 7174
rect 517866 6938 518102 7174
rect 517546 6618 517782 6854
rect 517866 6618 518102 6854
rect 518946 -1542 519182 -1306
rect 519266 -1542 519502 -1306
rect 518946 -1862 519182 -1626
rect 519266 -1862 519502 -1626
rect 517546 -2502 517782 -2266
rect 517866 -2502 518102 -2266
rect 517546 -2822 517782 -2586
rect 517866 -2822 518102 -2586
rect 516146 -5382 516382 -5146
rect 516466 -5382 516702 -5146
rect 516146 -5702 516382 -5466
rect 516466 -5702 516702 -5466
rect 514746 -6342 514982 -6106
rect 515066 -6342 515302 -6106
rect 514746 -6662 514982 -6426
rect 515066 -6662 515302 -6426
rect 521266 10658 521502 10894
rect 521586 10658 521822 10894
rect 521266 10338 521502 10574
rect 521586 10338 521822 10574
rect 524066 3218 524302 3454
rect 524386 3218 524622 3454
rect 524066 2898 524302 3134
rect 524386 2898 524622 3134
rect 524066 -582 524302 -346
rect 524386 -582 524622 -346
rect 524066 -902 524302 -666
rect 524386 -902 524622 -666
rect 522666 -3462 522902 -3226
rect 522986 -3462 523222 -3226
rect 522666 -3782 522902 -3546
rect 522986 -3782 523222 -3546
rect 521266 -4422 521502 -4186
rect 521586 -4422 521822 -4186
rect 521266 -4742 521502 -4506
rect 521586 -4742 521822 -4506
rect 519866 -7302 520102 -7066
rect 520186 -7302 520422 -7066
rect 519866 -7622 520102 -7386
rect 520186 -7622 520422 -7386
rect 527786 6938 528022 7174
rect 528106 6938 528342 7174
rect 527786 6618 528022 6854
rect 528106 6618 528342 6854
rect 529186 -1542 529422 -1306
rect 529506 -1542 529742 -1306
rect 529186 -1862 529422 -1626
rect 529506 -1862 529742 -1626
rect 527786 -2502 528022 -2266
rect 528106 -2502 528342 -2266
rect 527786 -2822 528022 -2586
rect 528106 -2822 528342 -2586
rect 526386 -5382 526622 -5146
rect 526706 -5382 526942 -5146
rect 526386 -5702 526622 -5466
rect 526706 -5702 526942 -5466
rect 524986 -6342 525222 -6106
rect 525306 -6342 525542 -6106
rect 524986 -6662 525222 -6426
rect 525306 -6662 525542 -6426
rect 531506 10658 531742 10894
rect 531826 10658 532062 10894
rect 531506 10338 531742 10574
rect 531826 10338 532062 10574
rect 534306 3218 534542 3454
rect 534626 3218 534862 3454
rect 534306 2898 534542 3134
rect 534626 2898 534862 3134
rect 534306 -582 534542 -346
rect 534626 -582 534862 -346
rect 534306 -902 534542 -666
rect 534626 -902 534862 -666
rect 532906 -3462 533142 -3226
rect 533226 -3462 533462 -3226
rect 532906 -3782 533142 -3546
rect 533226 -3782 533462 -3546
rect 531506 -4422 531742 -4186
rect 531826 -4422 532062 -4186
rect 531506 -4742 531742 -4506
rect 531826 -4742 532062 -4506
rect 530106 -7302 530342 -7066
rect 530426 -7302 530662 -7066
rect 530106 -7622 530342 -7386
rect 530426 -7622 530662 -7386
rect 538026 6938 538262 7174
rect 538346 6938 538582 7174
rect 538026 6618 538262 6854
rect 538346 6618 538582 6854
rect 539426 -1542 539662 -1306
rect 539746 -1542 539982 -1306
rect 539426 -1862 539662 -1626
rect 539746 -1862 539982 -1626
rect 538026 -2502 538262 -2266
rect 538346 -2502 538582 -2266
rect 538026 -2822 538262 -2586
rect 538346 -2822 538582 -2586
rect 536626 -5382 536862 -5146
rect 536946 -5382 537182 -5146
rect 536626 -5702 536862 -5466
rect 536946 -5702 537182 -5466
rect 535226 -6342 535462 -6106
rect 535546 -6342 535782 -6106
rect 535226 -6662 535462 -6426
rect 535546 -6662 535782 -6426
rect 541746 10658 541982 10894
rect 542066 10658 542302 10894
rect 541746 10338 541982 10574
rect 542066 10338 542302 10574
rect 543146 707482 543382 707718
rect 543466 707482 543702 707718
rect 543146 707162 543382 707398
rect 543466 707162 543702 707398
rect 543146 672938 543382 673174
rect 543466 672938 543702 673174
rect 543146 672618 543382 672854
rect 543466 672618 543702 672854
rect 543146 636938 543382 637174
rect 543466 636938 543702 637174
rect 543146 636618 543382 636854
rect 543466 636618 543702 636854
rect 543146 600938 543382 601174
rect 543466 600938 543702 601174
rect 543146 600618 543382 600854
rect 543466 600618 543702 600854
rect 543146 564938 543382 565174
rect 543466 564938 543702 565174
rect 543146 564618 543382 564854
rect 543466 564618 543702 564854
rect 543146 528938 543382 529174
rect 543466 528938 543702 529174
rect 543146 528618 543382 528854
rect 543466 528618 543702 528854
rect 543146 492938 543382 493174
rect 543466 492938 543702 493174
rect 543146 492618 543382 492854
rect 543466 492618 543702 492854
rect 543146 456938 543382 457174
rect 543466 456938 543702 457174
rect 543146 456618 543382 456854
rect 543466 456618 543702 456854
rect 543146 420938 543382 421174
rect 543466 420938 543702 421174
rect 543146 420618 543382 420854
rect 543466 420618 543702 420854
rect 543146 384938 543382 385174
rect 543466 384938 543702 385174
rect 543146 384618 543382 384854
rect 543466 384618 543702 384854
rect 543146 348938 543382 349174
rect 543466 348938 543702 349174
rect 543146 348618 543382 348854
rect 543466 348618 543702 348854
rect 543146 312938 543382 313174
rect 543466 312938 543702 313174
rect 543146 312618 543382 312854
rect 543466 312618 543702 312854
rect 543146 276938 543382 277174
rect 543466 276938 543702 277174
rect 543146 276618 543382 276854
rect 543466 276618 543702 276854
rect 543146 240938 543382 241174
rect 543466 240938 543702 241174
rect 543146 240618 543382 240854
rect 543466 240618 543702 240854
rect 543146 204938 543382 205174
rect 543466 204938 543702 205174
rect 543146 204618 543382 204854
rect 543466 204618 543702 204854
rect 543146 168938 543382 169174
rect 543466 168938 543702 169174
rect 543146 168618 543382 168854
rect 543466 168618 543702 168854
rect 543146 132938 543382 133174
rect 543466 132938 543702 133174
rect 543146 132618 543382 132854
rect 543466 132618 543702 132854
rect 543146 96938 543382 97174
rect 543466 96938 543702 97174
rect 543146 96618 543382 96854
rect 543466 96618 543702 96854
rect 543146 60938 543382 61174
rect 543466 60938 543702 61174
rect 543146 60618 543382 60854
rect 543466 60618 543702 60854
rect 543146 24938 543382 25174
rect 543466 24938 543702 25174
rect 543146 24618 543382 24854
rect 543466 24618 543702 24854
rect 544546 704602 544782 704838
rect 544866 704602 545102 704838
rect 544546 704282 544782 704518
rect 544866 704282 545102 704518
rect 544546 687218 544782 687454
rect 544866 687218 545102 687454
rect 544546 686898 544782 687134
rect 544866 686898 545102 687134
rect 544546 651218 544782 651454
rect 544866 651218 545102 651454
rect 544546 650898 544782 651134
rect 544866 650898 545102 651134
rect 544546 615218 544782 615454
rect 544866 615218 545102 615454
rect 544546 614898 544782 615134
rect 544866 614898 545102 615134
rect 544546 579218 544782 579454
rect 544866 579218 545102 579454
rect 544546 578898 544782 579134
rect 544866 578898 545102 579134
rect 544546 543218 544782 543454
rect 544866 543218 545102 543454
rect 544546 542898 544782 543134
rect 544866 542898 545102 543134
rect 544546 507218 544782 507454
rect 544866 507218 545102 507454
rect 544546 506898 544782 507134
rect 544866 506898 545102 507134
rect 544546 471218 544782 471454
rect 544866 471218 545102 471454
rect 544546 470898 544782 471134
rect 544866 470898 545102 471134
rect 544546 435218 544782 435454
rect 544866 435218 545102 435454
rect 544546 434898 544782 435134
rect 544866 434898 545102 435134
rect 544546 399218 544782 399454
rect 544866 399218 545102 399454
rect 544546 398898 544782 399134
rect 544866 398898 545102 399134
rect 544546 363218 544782 363454
rect 544866 363218 545102 363454
rect 544546 362898 544782 363134
rect 544866 362898 545102 363134
rect 544546 327218 544782 327454
rect 544866 327218 545102 327454
rect 544546 326898 544782 327134
rect 544866 326898 545102 327134
rect 544546 291218 544782 291454
rect 544866 291218 545102 291454
rect 544546 290898 544782 291134
rect 544866 290898 545102 291134
rect 544546 255218 544782 255454
rect 544866 255218 545102 255454
rect 544546 254898 544782 255134
rect 544866 254898 545102 255134
rect 544546 219218 544782 219454
rect 544866 219218 545102 219454
rect 544546 218898 544782 219134
rect 544866 218898 545102 219134
rect 544546 183218 544782 183454
rect 544866 183218 545102 183454
rect 544546 182898 544782 183134
rect 544866 182898 545102 183134
rect 544546 147218 544782 147454
rect 544866 147218 545102 147454
rect 544546 146898 544782 147134
rect 544866 146898 545102 147134
rect 544546 111218 544782 111454
rect 544866 111218 545102 111454
rect 544546 110898 544782 111134
rect 544866 110898 545102 111134
rect 544546 75218 544782 75454
rect 544866 75218 545102 75454
rect 544546 74898 544782 75134
rect 544866 74898 545102 75134
rect 544546 39218 544782 39454
rect 544866 39218 545102 39454
rect 544546 38898 544782 39134
rect 544866 38898 545102 39134
rect 544546 3218 544782 3454
rect 544866 3218 545102 3454
rect 544546 2898 544782 3134
rect 544866 2898 545102 3134
rect 544546 -582 544782 -346
rect 544866 -582 545102 -346
rect 544546 -902 544782 -666
rect 544866 -902 545102 -666
rect 550586 711322 550822 711558
rect 550906 711322 551142 711558
rect 550586 711002 550822 711238
rect 550906 711002 551142 711238
rect 545466 698378 545702 698614
rect 545786 698378 546022 698614
rect 545466 698058 545702 698294
rect 545786 698058 546022 698294
rect 545466 662378 545702 662614
rect 545786 662378 546022 662614
rect 545466 662058 545702 662294
rect 545786 662058 546022 662294
rect 545466 626378 545702 626614
rect 545786 626378 546022 626614
rect 545466 626058 545702 626294
rect 545786 626058 546022 626294
rect 545466 590378 545702 590614
rect 545786 590378 546022 590614
rect 545466 590058 545702 590294
rect 545786 590058 546022 590294
rect 545466 554378 545702 554614
rect 545786 554378 546022 554614
rect 545466 554058 545702 554294
rect 545786 554058 546022 554294
rect 545466 518378 545702 518614
rect 545786 518378 546022 518614
rect 545466 518058 545702 518294
rect 545786 518058 546022 518294
rect 545466 482378 545702 482614
rect 545786 482378 546022 482614
rect 545466 482058 545702 482294
rect 545786 482058 546022 482294
rect 545466 446378 545702 446614
rect 545786 446378 546022 446614
rect 545466 446058 545702 446294
rect 545786 446058 546022 446294
rect 545466 410378 545702 410614
rect 545786 410378 546022 410614
rect 545466 410058 545702 410294
rect 545786 410058 546022 410294
rect 545466 374378 545702 374614
rect 545786 374378 546022 374614
rect 545466 374058 545702 374294
rect 545786 374058 546022 374294
rect 545466 338378 545702 338614
rect 545786 338378 546022 338614
rect 545466 338058 545702 338294
rect 545786 338058 546022 338294
rect 545466 302378 545702 302614
rect 545786 302378 546022 302614
rect 545466 302058 545702 302294
rect 545786 302058 546022 302294
rect 545466 266378 545702 266614
rect 545786 266378 546022 266614
rect 545466 266058 545702 266294
rect 545786 266058 546022 266294
rect 545466 230378 545702 230614
rect 545786 230378 546022 230614
rect 545466 230058 545702 230294
rect 545786 230058 546022 230294
rect 545466 194378 545702 194614
rect 545786 194378 546022 194614
rect 545466 194058 545702 194294
rect 545786 194058 546022 194294
rect 545466 158378 545702 158614
rect 545786 158378 546022 158614
rect 545466 158058 545702 158294
rect 545786 158058 546022 158294
rect 545466 122378 545702 122614
rect 545786 122378 546022 122614
rect 545466 122058 545702 122294
rect 545786 122058 546022 122294
rect 545466 86378 545702 86614
rect 545786 86378 546022 86614
rect 545466 86058 545702 86294
rect 545786 86058 546022 86294
rect 545466 50378 545702 50614
rect 545786 50378 546022 50614
rect 545466 50058 545702 50294
rect 545786 50058 546022 50294
rect 545466 14378 545702 14614
rect 545786 14378 546022 14614
rect 545466 14058 545702 14294
rect 545786 14058 546022 14294
rect 543146 -3462 543382 -3226
rect 543466 -3462 543702 -3226
rect 543146 -3782 543382 -3546
rect 543466 -3782 543702 -3546
rect 541746 -4422 541982 -4186
rect 542066 -4422 542302 -4186
rect 541746 -4742 541982 -4506
rect 542066 -4742 542302 -4506
rect 540346 -7302 540582 -7066
rect 540666 -7302 540902 -7066
rect 540346 -7622 540582 -7386
rect 540666 -7622 540902 -7386
rect 546866 709402 547102 709638
rect 547186 709402 547422 709638
rect 546866 709082 547102 709318
rect 547186 709082 547422 709318
rect 546866 676658 547102 676894
rect 547186 676658 547422 676894
rect 546866 676338 547102 676574
rect 547186 676338 547422 676574
rect 546866 640658 547102 640894
rect 547186 640658 547422 640894
rect 546866 640338 547102 640574
rect 547186 640338 547422 640574
rect 546866 604658 547102 604894
rect 547186 604658 547422 604894
rect 546866 604338 547102 604574
rect 547186 604338 547422 604574
rect 546866 568658 547102 568894
rect 547186 568658 547422 568894
rect 546866 568338 547102 568574
rect 547186 568338 547422 568574
rect 546866 532658 547102 532894
rect 547186 532658 547422 532894
rect 546866 532338 547102 532574
rect 547186 532338 547422 532574
rect 546866 496658 547102 496894
rect 547186 496658 547422 496894
rect 546866 496338 547102 496574
rect 547186 496338 547422 496574
rect 546866 460658 547102 460894
rect 547186 460658 547422 460894
rect 546866 460338 547102 460574
rect 547186 460338 547422 460574
rect 546866 424658 547102 424894
rect 547186 424658 547422 424894
rect 546866 424338 547102 424574
rect 547186 424338 547422 424574
rect 546866 388658 547102 388894
rect 547186 388658 547422 388894
rect 546866 388338 547102 388574
rect 547186 388338 547422 388574
rect 546866 352658 547102 352894
rect 547186 352658 547422 352894
rect 546866 352338 547102 352574
rect 547186 352338 547422 352574
rect 546866 316658 547102 316894
rect 547186 316658 547422 316894
rect 546866 316338 547102 316574
rect 547186 316338 547422 316574
rect 546866 280658 547102 280894
rect 547186 280658 547422 280894
rect 546866 280338 547102 280574
rect 547186 280338 547422 280574
rect 546866 244658 547102 244894
rect 547186 244658 547422 244894
rect 546866 244338 547102 244574
rect 547186 244338 547422 244574
rect 546866 208658 547102 208894
rect 547186 208658 547422 208894
rect 546866 208338 547102 208574
rect 547186 208338 547422 208574
rect 546866 172658 547102 172894
rect 547186 172658 547422 172894
rect 546866 172338 547102 172574
rect 547186 172338 547422 172574
rect 546866 136658 547102 136894
rect 547186 136658 547422 136894
rect 546866 136338 547102 136574
rect 547186 136338 547422 136574
rect 546866 100658 547102 100894
rect 547186 100658 547422 100894
rect 546866 100338 547102 100574
rect 547186 100338 547422 100574
rect 546866 64658 547102 64894
rect 547186 64658 547422 64894
rect 546866 64338 547102 64574
rect 547186 64338 547422 64574
rect 546866 28658 547102 28894
rect 547186 28658 547422 28894
rect 546866 28338 547102 28574
rect 547186 28338 547422 28574
rect 548266 706522 548502 706758
rect 548586 706522 548822 706758
rect 548266 706202 548502 706438
rect 548586 706202 548822 706438
rect 548266 690938 548502 691174
rect 548586 690938 548822 691174
rect 548266 690618 548502 690854
rect 548586 690618 548822 690854
rect 548266 654938 548502 655174
rect 548586 654938 548822 655174
rect 548266 654618 548502 654854
rect 548586 654618 548822 654854
rect 548266 618938 548502 619174
rect 548586 618938 548822 619174
rect 548266 618618 548502 618854
rect 548586 618618 548822 618854
rect 548266 582938 548502 583174
rect 548586 582938 548822 583174
rect 548266 582618 548502 582854
rect 548586 582618 548822 582854
rect 548266 546938 548502 547174
rect 548586 546938 548822 547174
rect 548266 546618 548502 546854
rect 548586 546618 548822 546854
rect 548266 510938 548502 511174
rect 548586 510938 548822 511174
rect 548266 510618 548502 510854
rect 548586 510618 548822 510854
rect 548266 474938 548502 475174
rect 548586 474938 548822 475174
rect 548266 474618 548502 474854
rect 548586 474618 548822 474854
rect 548266 438938 548502 439174
rect 548586 438938 548822 439174
rect 548266 438618 548502 438854
rect 548586 438618 548822 438854
rect 548266 402938 548502 403174
rect 548586 402938 548822 403174
rect 548266 402618 548502 402854
rect 548586 402618 548822 402854
rect 548266 366938 548502 367174
rect 548586 366938 548822 367174
rect 548266 366618 548502 366854
rect 548586 366618 548822 366854
rect 548266 330938 548502 331174
rect 548586 330938 548822 331174
rect 548266 330618 548502 330854
rect 548586 330618 548822 330854
rect 548266 294938 548502 295174
rect 548586 294938 548822 295174
rect 548266 294618 548502 294854
rect 548586 294618 548822 294854
rect 548266 258938 548502 259174
rect 548586 258938 548822 259174
rect 548266 258618 548502 258854
rect 548586 258618 548822 258854
rect 548266 222938 548502 223174
rect 548586 222938 548822 223174
rect 548266 222618 548502 222854
rect 548586 222618 548822 222854
rect 548266 186938 548502 187174
rect 548586 186938 548822 187174
rect 548266 186618 548502 186854
rect 548586 186618 548822 186854
rect 548266 150938 548502 151174
rect 548586 150938 548822 151174
rect 548266 150618 548502 150854
rect 548586 150618 548822 150854
rect 548266 114938 548502 115174
rect 548586 114938 548822 115174
rect 548266 114618 548502 114854
rect 548586 114618 548822 114854
rect 548266 78938 548502 79174
rect 548586 78938 548822 79174
rect 548266 78618 548502 78854
rect 548586 78618 548822 78854
rect 548266 42938 548502 43174
rect 548586 42938 548822 43174
rect 548266 42618 548502 42854
rect 548586 42618 548822 42854
rect 548266 6938 548502 7174
rect 548586 6938 548822 7174
rect 548266 6618 548502 6854
rect 548586 6618 548822 6854
rect 549666 705562 549902 705798
rect 549986 705562 550222 705798
rect 549666 705242 549902 705478
rect 549986 705242 550222 705478
rect 549666 669218 549902 669454
rect 549986 669218 550222 669454
rect 549666 668898 549902 669134
rect 549986 668898 550222 669134
rect 549666 633218 549902 633454
rect 549986 633218 550222 633454
rect 549666 632898 549902 633134
rect 549986 632898 550222 633134
rect 549666 597218 549902 597454
rect 549986 597218 550222 597454
rect 549666 596898 549902 597134
rect 549986 596898 550222 597134
rect 549666 561218 549902 561454
rect 549986 561218 550222 561454
rect 549666 560898 549902 561134
rect 549986 560898 550222 561134
rect 549666 525218 549902 525454
rect 549986 525218 550222 525454
rect 549666 524898 549902 525134
rect 549986 524898 550222 525134
rect 549666 489218 549902 489454
rect 549986 489218 550222 489454
rect 549666 488898 549902 489134
rect 549986 488898 550222 489134
rect 549666 453218 549902 453454
rect 549986 453218 550222 453454
rect 549666 452898 549902 453134
rect 549986 452898 550222 453134
rect 549666 417218 549902 417454
rect 549986 417218 550222 417454
rect 549666 416898 549902 417134
rect 549986 416898 550222 417134
rect 549666 381218 549902 381454
rect 549986 381218 550222 381454
rect 549666 380898 549902 381134
rect 549986 380898 550222 381134
rect 549666 345218 549902 345454
rect 549986 345218 550222 345454
rect 549666 344898 549902 345134
rect 549986 344898 550222 345134
rect 549666 309218 549902 309454
rect 549986 309218 550222 309454
rect 549666 308898 549902 309134
rect 549986 308898 550222 309134
rect 549666 273218 549902 273454
rect 549986 273218 550222 273454
rect 549666 272898 549902 273134
rect 549986 272898 550222 273134
rect 549666 237218 549902 237454
rect 549986 237218 550222 237454
rect 549666 236898 549902 237134
rect 549986 236898 550222 237134
rect 549666 201218 549902 201454
rect 549986 201218 550222 201454
rect 549666 200898 549902 201134
rect 549986 200898 550222 201134
rect 549666 165218 549902 165454
rect 549986 165218 550222 165454
rect 549666 164898 549902 165134
rect 549986 164898 550222 165134
rect 549666 129218 549902 129454
rect 549986 129218 550222 129454
rect 549666 128898 549902 129134
rect 549986 128898 550222 129134
rect 549666 93218 549902 93454
rect 549986 93218 550222 93454
rect 549666 92898 549902 93134
rect 549986 92898 550222 93134
rect 549666 57218 549902 57454
rect 549986 57218 550222 57454
rect 549666 56898 549902 57134
rect 549986 56898 550222 57134
rect 549666 21218 549902 21454
rect 549986 21218 550222 21454
rect 549666 20898 549902 21134
rect 549986 20898 550222 21134
rect 549666 -1542 549902 -1306
rect 549986 -1542 550222 -1306
rect 549666 -1862 549902 -1626
rect 549986 -1862 550222 -1626
rect 555706 710362 555942 710598
rect 556026 710362 556262 710598
rect 555706 710042 555942 710278
rect 556026 710042 556262 710278
rect 550586 680378 550822 680614
rect 550906 680378 551142 680614
rect 550586 680058 550822 680294
rect 550906 680058 551142 680294
rect 550586 644378 550822 644614
rect 550906 644378 551142 644614
rect 550586 644058 550822 644294
rect 550906 644058 551142 644294
rect 550586 608378 550822 608614
rect 550906 608378 551142 608614
rect 550586 608058 550822 608294
rect 550906 608058 551142 608294
rect 550586 572378 550822 572614
rect 550906 572378 551142 572614
rect 550586 572058 550822 572294
rect 550906 572058 551142 572294
rect 550586 536378 550822 536614
rect 550906 536378 551142 536614
rect 550586 536058 550822 536294
rect 550906 536058 551142 536294
rect 550586 500378 550822 500614
rect 550906 500378 551142 500614
rect 550586 500058 550822 500294
rect 550906 500058 551142 500294
rect 550586 464378 550822 464614
rect 550906 464378 551142 464614
rect 550586 464058 550822 464294
rect 550906 464058 551142 464294
rect 550586 428378 550822 428614
rect 550906 428378 551142 428614
rect 550586 428058 550822 428294
rect 550906 428058 551142 428294
rect 550586 392378 550822 392614
rect 550906 392378 551142 392614
rect 550586 392058 550822 392294
rect 550906 392058 551142 392294
rect 550586 356378 550822 356614
rect 550906 356378 551142 356614
rect 550586 356058 550822 356294
rect 550906 356058 551142 356294
rect 550586 320378 550822 320614
rect 550906 320378 551142 320614
rect 550586 320058 550822 320294
rect 550906 320058 551142 320294
rect 550586 284378 550822 284614
rect 550906 284378 551142 284614
rect 550586 284058 550822 284294
rect 550906 284058 551142 284294
rect 550586 248378 550822 248614
rect 550906 248378 551142 248614
rect 550586 248058 550822 248294
rect 550906 248058 551142 248294
rect 550586 212378 550822 212614
rect 550906 212378 551142 212614
rect 550586 212058 550822 212294
rect 550906 212058 551142 212294
rect 550586 176378 550822 176614
rect 550906 176378 551142 176614
rect 550586 176058 550822 176294
rect 550906 176058 551142 176294
rect 550586 140378 550822 140614
rect 550906 140378 551142 140614
rect 550586 140058 550822 140294
rect 550906 140058 551142 140294
rect 550586 104378 550822 104614
rect 550906 104378 551142 104614
rect 550586 104058 550822 104294
rect 550906 104058 551142 104294
rect 550586 68378 550822 68614
rect 550906 68378 551142 68614
rect 550586 68058 550822 68294
rect 550906 68058 551142 68294
rect 550586 32378 550822 32614
rect 550906 32378 551142 32614
rect 550586 32058 550822 32294
rect 550906 32058 551142 32294
rect 548266 -2502 548502 -2266
rect 548586 -2502 548822 -2266
rect 548266 -2822 548502 -2586
rect 548586 -2822 548822 -2586
rect 546866 -5382 547102 -5146
rect 547186 -5382 547422 -5146
rect 546866 -5702 547102 -5466
rect 547186 -5702 547422 -5466
rect 545466 -6342 545702 -6106
rect 545786 -6342 546022 -6106
rect 545466 -6662 545702 -6426
rect 545786 -6662 546022 -6426
rect 551986 708442 552222 708678
rect 552306 708442 552542 708678
rect 551986 708122 552222 708358
rect 552306 708122 552542 708358
rect 551986 694658 552222 694894
rect 552306 694658 552542 694894
rect 551986 694338 552222 694574
rect 552306 694338 552542 694574
rect 551986 658658 552222 658894
rect 552306 658658 552542 658894
rect 551986 658338 552222 658574
rect 552306 658338 552542 658574
rect 551986 622658 552222 622894
rect 552306 622658 552542 622894
rect 551986 622338 552222 622574
rect 552306 622338 552542 622574
rect 551986 586658 552222 586894
rect 552306 586658 552542 586894
rect 551986 586338 552222 586574
rect 552306 586338 552542 586574
rect 551986 550658 552222 550894
rect 552306 550658 552542 550894
rect 551986 550338 552222 550574
rect 552306 550338 552542 550574
rect 551986 514658 552222 514894
rect 552306 514658 552542 514894
rect 551986 514338 552222 514574
rect 552306 514338 552542 514574
rect 551986 478658 552222 478894
rect 552306 478658 552542 478894
rect 551986 478338 552222 478574
rect 552306 478338 552542 478574
rect 551986 442658 552222 442894
rect 552306 442658 552542 442894
rect 551986 442338 552222 442574
rect 552306 442338 552542 442574
rect 551986 406658 552222 406894
rect 552306 406658 552542 406894
rect 551986 406338 552222 406574
rect 552306 406338 552542 406574
rect 551986 370658 552222 370894
rect 552306 370658 552542 370894
rect 551986 370338 552222 370574
rect 552306 370338 552542 370574
rect 551986 334658 552222 334894
rect 552306 334658 552542 334894
rect 551986 334338 552222 334574
rect 552306 334338 552542 334574
rect 551986 298658 552222 298894
rect 552306 298658 552542 298894
rect 551986 298338 552222 298574
rect 552306 298338 552542 298574
rect 551986 262658 552222 262894
rect 552306 262658 552542 262894
rect 551986 262338 552222 262574
rect 552306 262338 552542 262574
rect 551986 226658 552222 226894
rect 552306 226658 552542 226894
rect 551986 226338 552222 226574
rect 552306 226338 552542 226574
rect 551986 190658 552222 190894
rect 552306 190658 552542 190894
rect 551986 190338 552222 190574
rect 552306 190338 552542 190574
rect 551986 154658 552222 154894
rect 552306 154658 552542 154894
rect 551986 154338 552222 154574
rect 552306 154338 552542 154574
rect 551986 118658 552222 118894
rect 552306 118658 552542 118894
rect 551986 118338 552222 118574
rect 552306 118338 552542 118574
rect 551986 82658 552222 82894
rect 552306 82658 552542 82894
rect 551986 82338 552222 82574
rect 552306 82338 552542 82574
rect 551986 46658 552222 46894
rect 552306 46658 552542 46894
rect 551986 46338 552222 46574
rect 552306 46338 552542 46574
rect 551986 10658 552222 10894
rect 552306 10658 552542 10894
rect 551986 10338 552222 10574
rect 552306 10338 552542 10574
rect 553386 707482 553622 707718
rect 553706 707482 553942 707718
rect 553386 707162 553622 707398
rect 553706 707162 553942 707398
rect 553386 672938 553622 673174
rect 553706 672938 553942 673174
rect 553386 672618 553622 672854
rect 553706 672618 553942 672854
rect 553386 636938 553622 637174
rect 553706 636938 553942 637174
rect 553386 636618 553622 636854
rect 553706 636618 553942 636854
rect 553386 600938 553622 601174
rect 553706 600938 553942 601174
rect 553386 600618 553622 600854
rect 553706 600618 553942 600854
rect 553386 564938 553622 565174
rect 553706 564938 553942 565174
rect 553386 564618 553622 564854
rect 553706 564618 553942 564854
rect 553386 528938 553622 529174
rect 553706 528938 553942 529174
rect 553386 528618 553622 528854
rect 553706 528618 553942 528854
rect 553386 492938 553622 493174
rect 553706 492938 553942 493174
rect 553386 492618 553622 492854
rect 553706 492618 553942 492854
rect 553386 456938 553622 457174
rect 553706 456938 553942 457174
rect 553386 456618 553622 456854
rect 553706 456618 553942 456854
rect 553386 420938 553622 421174
rect 553706 420938 553942 421174
rect 553386 420618 553622 420854
rect 553706 420618 553942 420854
rect 553386 384938 553622 385174
rect 553706 384938 553942 385174
rect 553386 384618 553622 384854
rect 553706 384618 553942 384854
rect 553386 348938 553622 349174
rect 553706 348938 553942 349174
rect 553386 348618 553622 348854
rect 553706 348618 553942 348854
rect 553386 312938 553622 313174
rect 553706 312938 553942 313174
rect 553386 312618 553622 312854
rect 553706 312618 553942 312854
rect 553386 276938 553622 277174
rect 553706 276938 553942 277174
rect 553386 276618 553622 276854
rect 553706 276618 553942 276854
rect 553386 240938 553622 241174
rect 553706 240938 553942 241174
rect 553386 240618 553622 240854
rect 553706 240618 553942 240854
rect 553386 204938 553622 205174
rect 553706 204938 553942 205174
rect 553386 204618 553622 204854
rect 553706 204618 553942 204854
rect 553386 168938 553622 169174
rect 553706 168938 553942 169174
rect 553386 168618 553622 168854
rect 553706 168618 553942 168854
rect 553386 132938 553622 133174
rect 553706 132938 553942 133174
rect 553386 132618 553622 132854
rect 553706 132618 553942 132854
rect 553386 96938 553622 97174
rect 553706 96938 553942 97174
rect 553386 96618 553622 96854
rect 553706 96618 553942 96854
rect 553386 60938 553622 61174
rect 553706 60938 553942 61174
rect 553386 60618 553622 60854
rect 553706 60618 553942 60854
rect 553386 24938 553622 25174
rect 553706 24938 553942 25174
rect 553386 24618 553622 24854
rect 553706 24618 553942 24854
rect 554786 704602 555022 704838
rect 555106 704602 555342 704838
rect 554786 704282 555022 704518
rect 555106 704282 555342 704518
rect 554786 687218 555022 687454
rect 555106 687218 555342 687454
rect 554786 686898 555022 687134
rect 555106 686898 555342 687134
rect 554786 651218 555022 651454
rect 555106 651218 555342 651454
rect 554786 650898 555022 651134
rect 555106 650898 555342 651134
rect 554786 615218 555022 615454
rect 555106 615218 555342 615454
rect 554786 614898 555022 615134
rect 555106 614898 555342 615134
rect 554786 579218 555022 579454
rect 555106 579218 555342 579454
rect 554786 578898 555022 579134
rect 555106 578898 555342 579134
rect 554786 543218 555022 543454
rect 555106 543218 555342 543454
rect 554786 542898 555022 543134
rect 555106 542898 555342 543134
rect 554786 507218 555022 507454
rect 555106 507218 555342 507454
rect 554786 506898 555022 507134
rect 555106 506898 555342 507134
rect 554786 471218 555022 471454
rect 555106 471218 555342 471454
rect 554786 470898 555022 471134
rect 555106 470898 555342 471134
rect 554786 435218 555022 435454
rect 555106 435218 555342 435454
rect 554786 434898 555022 435134
rect 555106 434898 555342 435134
rect 554786 399218 555022 399454
rect 555106 399218 555342 399454
rect 554786 398898 555022 399134
rect 555106 398898 555342 399134
rect 554786 363218 555022 363454
rect 555106 363218 555342 363454
rect 554786 362898 555022 363134
rect 555106 362898 555342 363134
rect 554786 327218 555022 327454
rect 555106 327218 555342 327454
rect 554786 326898 555022 327134
rect 555106 326898 555342 327134
rect 554786 291218 555022 291454
rect 555106 291218 555342 291454
rect 554786 290898 555022 291134
rect 555106 290898 555342 291134
rect 554786 255218 555022 255454
rect 555106 255218 555342 255454
rect 554786 254898 555022 255134
rect 555106 254898 555342 255134
rect 554786 219218 555022 219454
rect 555106 219218 555342 219454
rect 554786 218898 555022 219134
rect 555106 218898 555342 219134
rect 554786 183218 555022 183454
rect 555106 183218 555342 183454
rect 554786 182898 555022 183134
rect 555106 182898 555342 183134
rect 554786 147218 555022 147454
rect 555106 147218 555342 147454
rect 554786 146898 555022 147134
rect 555106 146898 555342 147134
rect 554786 111218 555022 111454
rect 555106 111218 555342 111454
rect 554786 110898 555022 111134
rect 555106 110898 555342 111134
rect 554786 75218 555022 75454
rect 555106 75218 555342 75454
rect 554786 74898 555022 75134
rect 555106 74898 555342 75134
rect 554786 39218 555022 39454
rect 555106 39218 555342 39454
rect 554786 38898 555022 39134
rect 555106 38898 555342 39134
rect 554786 3218 555022 3454
rect 555106 3218 555342 3454
rect 554786 2898 555022 3134
rect 555106 2898 555342 3134
rect 554786 -582 555022 -346
rect 555106 -582 555342 -346
rect 554786 -902 555022 -666
rect 555106 -902 555342 -666
rect 560826 711322 561062 711558
rect 561146 711322 561382 711558
rect 560826 711002 561062 711238
rect 561146 711002 561382 711238
rect 555706 698378 555942 698614
rect 556026 698378 556262 698614
rect 555706 698058 555942 698294
rect 556026 698058 556262 698294
rect 555706 662378 555942 662614
rect 556026 662378 556262 662614
rect 555706 662058 555942 662294
rect 556026 662058 556262 662294
rect 555706 626378 555942 626614
rect 556026 626378 556262 626614
rect 555706 626058 555942 626294
rect 556026 626058 556262 626294
rect 555706 590378 555942 590614
rect 556026 590378 556262 590614
rect 555706 590058 555942 590294
rect 556026 590058 556262 590294
rect 555706 554378 555942 554614
rect 556026 554378 556262 554614
rect 555706 554058 555942 554294
rect 556026 554058 556262 554294
rect 555706 518378 555942 518614
rect 556026 518378 556262 518614
rect 555706 518058 555942 518294
rect 556026 518058 556262 518294
rect 555706 482378 555942 482614
rect 556026 482378 556262 482614
rect 555706 482058 555942 482294
rect 556026 482058 556262 482294
rect 555706 446378 555942 446614
rect 556026 446378 556262 446614
rect 555706 446058 555942 446294
rect 556026 446058 556262 446294
rect 555706 410378 555942 410614
rect 556026 410378 556262 410614
rect 555706 410058 555942 410294
rect 556026 410058 556262 410294
rect 555706 374378 555942 374614
rect 556026 374378 556262 374614
rect 555706 374058 555942 374294
rect 556026 374058 556262 374294
rect 555706 338378 555942 338614
rect 556026 338378 556262 338614
rect 555706 338058 555942 338294
rect 556026 338058 556262 338294
rect 555706 302378 555942 302614
rect 556026 302378 556262 302614
rect 555706 302058 555942 302294
rect 556026 302058 556262 302294
rect 555706 266378 555942 266614
rect 556026 266378 556262 266614
rect 555706 266058 555942 266294
rect 556026 266058 556262 266294
rect 555706 230378 555942 230614
rect 556026 230378 556262 230614
rect 555706 230058 555942 230294
rect 556026 230058 556262 230294
rect 555706 194378 555942 194614
rect 556026 194378 556262 194614
rect 555706 194058 555942 194294
rect 556026 194058 556262 194294
rect 555706 158378 555942 158614
rect 556026 158378 556262 158614
rect 555706 158058 555942 158294
rect 556026 158058 556262 158294
rect 555706 122378 555942 122614
rect 556026 122378 556262 122614
rect 555706 122058 555942 122294
rect 556026 122058 556262 122294
rect 555706 86378 555942 86614
rect 556026 86378 556262 86614
rect 555706 86058 555942 86294
rect 556026 86058 556262 86294
rect 555706 50378 555942 50614
rect 556026 50378 556262 50614
rect 555706 50058 555942 50294
rect 556026 50058 556262 50294
rect 555706 14378 555942 14614
rect 556026 14378 556262 14614
rect 555706 14058 555942 14294
rect 556026 14058 556262 14294
rect 553386 -3462 553622 -3226
rect 553706 -3462 553942 -3226
rect 553386 -3782 553622 -3546
rect 553706 -3782 553942 -3546
rect 551986 -4422 552222 -4186
rect 552306 -4422 552542 -4186
rect 551986 -4742 552222 -4506
rect 552306 -4742 552542 -4506
rect 550586 -7302 550822 -7066
rect 550906 -7302 551142 -7066
rect 550586 -7622 550822 -7386
rect 550906 -7622 551142 -7386
rect 557106 709402 557342 709638
rect 557426 709402 557662 709638
rect 557106 709082 557342 709318
rect 557426 709082 557662 709318
rect 557106 676658 557342 676894
rect 557426 676658 557662 676894
rect 557106 676338 557342 676574
rect 557426 676338 557662 676574
rect 557106 640658 557342 640894
rect 557426 640658 557662 640894
rect 557106 640338 557342 640574
rect 557426 640338 557662 640574
rect 557106 604658 557342 604894
rect 557426 604658 557662 604894
rect 557106 604338 557342 604574
rect 557426 604338 557662 604574
rect 557106 568658 557342 568894
rect 557426 568658 557662 568894
rect 557106 568338 557342 568574
rect 557426 568338 557662 568574
rect 557106 532658 557342 532894
rect 557426 532658 557662 532894
rect 557106 532338 557342 532574
rect 557426 532338 557662 532574
rect 557106 496658 557342 496894
rect 557426 496658 557662 496894
rect 557106 496338 557342 496574
rect 557426 496338 557662 496574
rect 557106 460658 557342 460894
rect 557426 460658 557662 460894
rect 557106 460338 557342 460574
rect 557426 460338 557662 460574
rect 557106 424658 557342 424894
rect 557426 424658 557662 424894
rect 557106 424338 557342 424574
rect 557426 424338 557662 424574
rect 557106 388658 557342 388894
rect 557426 388658 557662 388894
rect 557106 388338 557342 388574
rect 557426 388338 557662 388574
rect 557106 352658 557342 352894
rect 557426 352658 557662 352894
rect 557106 352338 557342 352574
rect 557426 352338 557662 352574
rect 557106 316658 557342 316894
rect 557426 316658 557662 316894
rect 557106 316338 557342 316574
rect 557426 316338 557662 316574
rect 557106 280658 557342 280894
rect 557426 280658 557662 280894
rect 557106 280338 557342 280574
rect 557426 280338 557662 280574
rect 557106 244658 557342 244894
rect 557426 244658 557662 244894
rect 557106 244338 557342 244574
rect 557426 244338 557662 244574
rect 557106 208658 557342 208894
rect 557426 208658 557662 208894
rect 557106 208338 557342 208574
rect 557426 208338 557662 208574
rect 557106 172658 557342 172894
rect 557426 172658 557662 172894
rect 557106 172338 557342 172574
rect 557426 172338 557662 172574
rect 557106 136658 557342 136894
rect 557426 136658 557662 136894
rect 557106 136338 557342 136574
rect 557426 136338 557662 136574
rect 557106 100658 557342 100894
rect 557426 100658 557662 100894
rect 557106 100338 557342 100574
rect 557426 100338 557662 100574
rect 557106 64658 557342 64894
rect 557426 64658 557662 64894
rect 557106 64338 557342 64574
rect 557426 64338 557662 64574
rect 557106 28658 557342 28894
rect 557426 28658 557662 28894
rect 557106 28338 557342 28574
rect 557426 28338 557662 28574
rect 558506 706522 558742 706758
rect 558826 706522 559062 706758
rect 558506 706202 558742 706438
rect 558826 706202 559062 706438
rect 558506 690938 558742 691174
rect 558826 690938 559062 691174
rect 558506 690618 558742 690854
rect 558826 690618 559062 690854
rect 558506 654938 558742 655174
rect 558826 654938 559062 655174
rect 558506 654618 558742 654854
rect 558826 654618 559062 654854
rect 558506 618938 558742 619174
rect 558826 618938 559062 619174
rect 558506 618618 558742 618854
rect 558826 618618 559062 618854
rect 558506 582938 558742 583174
rect 558826 582938 559062 583174
rect 558506 582618 558742 582854
rect 558826 582618 559062 582854
rect 558506 546938 558742 547174
rect 558826 546938 559062 547174
rect 558506 546618 558742 546854
rect 558826 546618 559062 546854
rect 558506 510938 558742 511174
rect 558826 510938 559062 511174
rect 558506 510618 558742 510854
rect 558826 510618 559062 510854
rect 558506 474938 558742 475174
rect 558826 474938 559062 475174
rect 558506 474618 558742 474854
rect 558826 474618 559062 474854
rect 558506 438938 558742 439174
rect 558826 438938 559062 439174
rect 558506 438618 558742 438854
rect 558826 438618 559062 438854
rect 558506 402938 558742 403174
rect 558826 402938 559062 403174
rect 558506 402618 558742 402854
rect 558826 402618 559062 402854
rect 558506 366938 558742 367174
rect 558826 366938 559062 367174
rect 558506 366618 558742 366854
rect 558826 366618 559062 366854
rect 558506 330938 558742 331174
rect 558826 330938 559062 331174
rect 558506 330618 558742 330854
rect 558826 330618 559062 330854
rect 558506 294938 558742 295174
rect 558826 294938 559062 295174
rect 558506 294618 558742 294854
rect 558826 294618 559062 294854
rect 558506 258938 558742 259174
rect 558826 258938 559062 259174
rect 558506 258618 558742 258854
rect 558826 258618 559062 258854
rect 558506 222938 558742 223174
rect 558826 222938 559062 223174
rect 558506 222618 558742 222854
rect 558826 222618 559062 222854
rect 558506 186938 558742 187174
rect 558826 186938 559062 187174
rect 558506 186618 558742 186854
rect 558826 186618 559062 186854
rect 558506 150938 558742 151174
rect 558826 150938 559062 151174
rect 558506 150618 558742 150854
rect 558826 150618 559062 150854
rect 558506 114938 558742 115174
rect 558826 114938 559062 115174
rect 558506 114618 558742 114854
rect 558826 114618 559062 114854
rect 558506 78938 558742 79174
rect 558826 78938 559062 79174
rect 558506 78618 558742 78854
rect 558826 78618 559062 78854
rect 558506 42938 558742 43174
rect 558826 42938 559062 43174
rect 558506 42618 558742 42854
rect 558826 42618 559062 42854
rect 558506 6938 558742 7174
rect 558826 6938 559062 7174
rect 558506 6618 558742 6854
rect 558826 6618 559062 6854
rect 559906 705562 560142 705798
rect 560226 705562 560462 705798
rect 559906 705242 560142 705478
rect 560226 705242 560462 705478
rect 559906 669218 560142 669454
rect 560226 669218 560462 669454
rect 559906 668898 560142 669134
rect 560226 668898 560462 669134
rect 559906 633218 560142 633454
rect 560226 633218 560462 633454
rect 559906 632898 560142 633134
rect 560226 632898 560462 633134
rect 559906 597218 560142 597454
rect 560226 597218 560462 597454
rect 559906 596898 560142 597134
rect 560226 596898 560462 597134
rect 559906 561218 560142 561454
rect 560226 561218 560462 561454
rect 559906 560898 560142 561134
rect 560226 560898 560462 561134
rect 559906 525218 560142 525454
rect 560226 525218 560462 525454
rect 559906 524898 560142 525134
rect 560226 524898 560462 525134
rect 559906 489218 560142 489454
rect 560226 489218 560462 489454
rect 559906 488898 560142 489134
rect 560226 488898 560462 489134
rect 559906 453218 560142 453454
rect 560226 453218 560462 453454
rect 559906 452898 560142 453134
rect 560226 452898 560462 453134
rect 559906 417218 560142 417454
rect 560226 417218 560462 417454
rect 559906 416898 560142 417134
rect 560226 416898 560462 417134
rect 559906 381218 560142 381454
rect 560226 381218 560462 381454
rect 559906 380898 560142 381134
rect 560226 380898 560462 381134
rect 559906 345218 560142 345454
rect 560226 345218 560462 345454
rect 559906 344898 560142 345134
rect 560226 344898 560462 345134
rect 559906 309218 560142 309454
rect 560226 309218 560462 309454
rect 559906 308898 560142 309134
rect 560226 308898 560462 309134
rect 559906 273218 560142 273454
rect 560226 273218 560462 273454
rect 559906 272898 560142 273134
rect 560226 272898 560462 273134
rect 559906 237218 560142 237454
rect 560226 237218 560462 237454
rect 559906 236898 560142 237134
rect 560226 236898 560462 237134
rect 559906 201218 560142 201454
rect 560226 201218 560462 201454
rect 559906 200898 560142 201134
rect 560226 200898 560462 201134
rect 559906 165218 560142 165454
rect 560226 165218 560462 165454
rect 559906 164898 560142 165134
rect 560226 164898 560462 165134
rect 559906 129218 560142 129454
rect 560226 129218 560462 129454
rect 559906 128898 560142 129134
rect 560226 128898 560462 129134
rect 559906 93218 560142 93454
rect 560226 93218 560462 93454
rect 559906 92898 560142 93134
rect 560226 92898 560462 93134
rect 559906 57218 560142 57454
rect 560226 57218 560462 57454
rect 559906 56898 560142 57134
rect 560226 56898 560462 57134
rect 559906 21218 560142 21454
rect 560226 21218 560462 21454
rect 559906 20898 560142 21134
rect 560226 20898 560462 21134
rect 559906 -1542 560142 -1306
rect 560226 -1542 560462 -1306
rect 559906 -1862 560142 -1626
rect 560226 -1862 560462 -1626
rect 565946 710362 566182 710598
rect 566266 710362 566502 710598
rect 565946 710042 566182 710278
rect 566266 710042 566502 710278
rect 560826 680378 561062 680614
rect 561146 680378 561382 680614
rect 560826 680058 561062 680294
rect 561146 680058 561382 680294
rect 560826 644378 561062 644614
rect 561146 644378 561382 644614
rect 560826 644058 561062 644294
rect 561146 644058 561382 644294
rect 560826 608378 561062 608614
rect 561146 608378 561382 608614
rect 560826 608058 561062 608294
rect 561146 608058 561382 608294
rect 560826 572378 561062 572614
rect 561146 572378 561382 572614
rect 560826 572058 561062 572294
rect 561146 572058 561382 572294
rect 560826 536378 561062 536614
rect 561146 536378 561382 536614
rect 560826 536058 561062 536294
rect 561146 536058 561382 536294
rect 560826 500378 561062 500614
rect 561146 500378 561382 500614
rect 560826 500058 561062 500294
rect 561146 500058 561382 500294
rect 560826 464378 561062 464614
rect 561146 464378 561382 464614
rect 560826 464058 561062 464294
rect 561146 464058 561382 464294
rect 560826 428378 561062 428614
rect 561146 428378 561382 428614
rect 560826 428058 561062 428294
rect 561146 428058 561382 428294
rect 560826 392378 561062 392614
rect 561146 392378 561382 392614
rect 560826 392058 561062 392294
rect 561146 392058 561382 392294
rect 560826 356378 561062 356614
rect 561146 356378 561382 356614
rect 560826 356058 561062 356294
rect 561146 356058 561382 356294
rect 560826 320378 561062 320614
rect 561146 320378 561382 320614
rect 560826 320058 561062 320294
rect 561146 320058 561382 320294
rect 560826 284378 561062 284614
rect 561146 284378 561382 284614
rect 560826 284058 561062 284294
rect 561146 284058 561382 284294
rect 560826 248378 561062 248614
rect 561146 248378 561382 248614
rect 560826 248058 561062 248294
rect 561146 248058 561382 248294
rect 560826 212378 561062 212614
rect 561146 212378 561382 212614
rect 560826 212058 561062 212294
rect 561146 212058 561382 212294
rect 560826 176378 561062 176614
rect 561146 176378 561382 176614
rect 560826 176058 561062 176294
rect 561146 176058 561382 176294
rect 560826 140378 561062 140614
rect 561146 140378 561382 140614
rect 560826 140058 561062 140294
rect 561146 140058 561382 140294
rect 560826 104378 561062 104614
rect 561146 104378 561382 104614
rect 560826 104058 561062 104294
rect 561146 104058 561382 104294
rect 560826 68378 561062 68614
rect 561146 68378 561382 68614
rect 560826 68058 561062 68294
rect 561146 68058 561382 68294
rect 560826 32378 561062 32614
rect 561146 32378 561382 32614
rect 560826 32058 561062 32294
rect 561146 32058 561382 32294
rect 558506 -2502 558742 -2266
rect 558826 -2502 559062 -2266
rect 558506 -2822 558742 -2586
rect 558826 -2822 559062 -2586
rect 557106 -5382 557342 -5146
rect 557426 -5382 557662 -5146
rect 557106 -5702 557342 -5466
rect 557426 -5702 557662 -5466
rect 555706 -6342 555942 -6106
rect 556026 -6342 556262 -6106
rect 555706 -6662 555942 -6426
rect 556026 -6662 556262 -6426
rect 562226 708442 562462 708678
rect 562546 708442 562782 708678
rect 562226 708122 562462 708358
rect 562546 708122 562782 708358
rect 562226 694658 562462 694894
rect 562546 694658 562782 694894
rect 562226 694338 562462 694574
rect 562546 694338 562782 694574
rect 562226 658658 562462 658894
rect 562546 658658 562782 658894
rect 562226 658338 562462 658574
rect 562546 658338 562782 658574
rect 562226 622658 562462 622894
rect 562546 622658 562782 622894
rect 562226 622338 562462 622574
rect 562546 622338 562782 622574
rect 562226 586658 562462 586894
rect 562546 586658 562782 586894
rect 562226 586338 562462 586574
rect 562546 586338 562782 586574
rect 562226 550658 562462 550894
rect 562546 550658 562782 550894
rect 562226 550338 562462 550574
rect 562546 550338 562782 550574
rect 562226 514658 562462 514894
rect 562546 514658 562782 514894
rect 562226 514338 562462 514574
rect 562546 514338 562782 514574
rect 562226 478658 562462 478894
rect 562546 478658 562782 478894
rect 562226 478338 562462 478574
rect 562546 478338 562782 478574
rect 562226 442658 562462 442894
rect 562546 442658 562782 442894
rect 562226 442338 562462 442574
rect 562546 442338 562782 442574
rect 562226 406658 562462 406894
rect 562546 406658 562782 406894
rect 562226 406338 562462 406574
rect 562546 406338 562782 406574
rect 562226 370658 562462 370894
rect 562546 370658 562782 370894
rect 562226 370338 562462 370574
rect 562546 370338 562782 370574
rect 562226 334658 562462 334894
rect 562546 334658 562782 334894
rect 562226 334338 562462 334574
rect 562546 334338 562782 334574
rect 562226 298658 562462 298894
rect 562546 298658 562782 298894
rect 562226 298338 562462 298574
rect 562546 298338 562782 298574
rect 562226 262658 562462 262894
rect 562546 262658 562782 262894
rect 562226 262338 562462 262574
rect 562546 262338 562782 262574
rect 562226 226658 562462 226894
rect 562546 226658 562782 226894
rect 562226 226338 562462 226574
rect 562546 226338 562782 226574
rect 562226 190658 562462 190894
rect 562546 190658 562782 190894
rect 562226 190338 562462 190574
rect 562546 190338 562782 190574
rect 562226 154658 562462 154894
rect 562546 154658 562782 154894
rect 562226 154338 562462 154574
rect 562546 154338 562782 154574
rect 562226 118658 562462 118894
rect 562546 118658 562782 118894
rect 562226 118338 562462 118574
rect 562546 118338 562782 118574
rect 562226 82658 562462 82894
rect 562546 82658 562782 82894
rect 562226 82338 562462 82574
rect 562546 82338 562782 82574
rect 562226 46658 562462 46894
rect 562546 46658 562782 46894
rect 562226 46338 562462 46574
rect 562546 46338 562782 46574
rect 562226 10658 562462 10894
rect 562546 10658 562782 10894
rect 562226 10338 562462 10574
rect 562546 10338 562782 10574
rect 563626 707482 563862 707718
rect 563946 707482 564182 707718
rect 563626 707162 563862 707398
rect 563946 707162 564182 707398
rect 563626 672938 563862 673174
rect 563946 672938 564182 673174
rect 563626 672618 563862 672854
rect 563946 672618 564182 672854
rect 563626 636938 563862 637174
rect 563946 636938 564182 637174
rect 563626 636618 563862 636854
rect 563946 636618 564182 636854
rect 563626 600938 563862 601174
rect 563946 600938 564182 601174
rect 563626 600618 563862 600854
rect 563946 600618 564182 600854
rect 563626 564938 563862 565174
rect 563946 564938 564182 565174
rect 563626 564618 563862 564854
rect 563946 564618 564182 564854
rect 563626 528938 563862 529174
rect 563946 528938 564182 529174
rect 563626 528618 563862 528854
rect 563946 528618 564182 528854
rect 563626 492938 563862 493174
rect 563946 492938 564182 493174
rect 563626 492618 563862 492854
rect 563946 492618 564182 492854
rect 563626 456938 563862 457174
rect 563946 456938 564182 457174
rect 563626 456618 563862 456854
rect 563946 456618 564182 456854
rect 563626 420938 563862 421174
rect 563946 420938 564182 421174
rect 563626 420618 563862 420854
rect 563946 420618 564182 420854
rect 563626 384938 563862 385174
rect 563946 384938 564182 385174
rect 563626 384618 563862 384854
rect 563946 384618 564182 384854
rect 563626 348938 563862 349174
rect 563946 348938 564182 349174
rect 563626 348618 563862 348854
rect 563946 348618 564182 348854
rect 563626 312938 563862 313174
rect 563946 312938 564182 313174
rect 563626 312618 563862 312854
rect 563946 312618 564182 312854
rect 563626 276938 563862 277174
rect 563946 276938 564182 277174
rect 563626 276618 563862 276854
rect 563946 276618 564182 276854
rect 563626 240938 563862 241174
rect 563946 240938 564182 241174
rect 563626 240618 563862 240854
rect 563946 240618 564182 240854
rect 563626 204938 563862 205174
rect 563946 204938 564182 205174
rect 563626 204618 563862 204854
rect 563946 204618 564182 204854
rect 563626 168938 563862 169174
rect 563946 168938 564182 169174
rect 563626 168618 563862 168854
rect 563946 168618 564182 168854
rect 563626 132938 563862 133174
rect 563946 132938 564182 133174
rect 563626 132618 563862 132854
rect 563946 132618 564182 132854
rect 563626 96938 563862 97174
rect 563946 96938 564182 97174
rect 563626 96618 563862 96854
rect 563946 96618 564182 96854
rect 563626 60938 563862 61174
rect 563946 60938 564182 61174
rect 563626 60618 563862 60854
rect 563946 60618 564182 60854
rect 563626 24938 563862 25174
rect 563946 24938 564182 25174
rect 563626 24618 563862 24854
rect 563946 24618 564182 24854
rect 565026 704602 565262 704838
rect 565346 704602 565582 704838
rect 565026 704282 565262 704518
rect 565346 704282 565582 704518
rect 565026 687218 565262 687454
rect 565346 687218 565582 687454
rect 565026 686898 565262 687134
rect 565346 686898 565582 687134
rect 565026 651218 565262 651454
rect 565346 651218 565582 651454
rect 565026 650898 565262 651134
rect 565346 650898 565582 651134
rect 565026 615218 565262 615454
rect 565346 615218 565582 615454
rect 565026 614898 565262 615134
rect 565346 614898 565582 615134
rect 565026 579218 565262 579454
rect 565346 579218 565582 579454
rect 565026 578898 565262 579134
rect 565346 578898 565582 579134
rect 565026 543218 565262 543454
rect 565346 543218 565582 543454
rect 565026 542898 565262 543134
rect 565346 542898 565582 543134
rect 565026 507218 565262 507454
rect 565346 507218 565582 507454
rect 565026 506898 565262 507134
rect 565346 506898 565582 507134
rect 565026 471218 565262 471454
rect 565346 471218 565582 471454
rect 565026 470898 565262 471134
rect 565346 470898 565582 471134
rect 565026 435218 565262 435454
rect 565346 435218 565582 435454
rect 565026 434898 565262 435134
rect 565346 434898 565582 435134
rect 565026 399218 565262 399454
rect 565346 399218 565582 399454
rect 565026 398898 565262 399134
rect 565346 398898 565582 399134
rect 565026 363218 565262 363454
rect 565346 363218 565582 363454
rect 565026 362898 565262 363134
rect 565346 362898 565582 363134
rect 565026 327218 565262 327454
rect 565346 327218 565582 327454
rect 565026 326898 565262 327134
rect 565346 326898 565582 327134
rect 565026 291218 565262 291454
rect 565346 291218 565582 291454
rect 565026 290898 565262 291134
rect 565346 290898 565582 291134
rect 565026 255218 565262 255454
rect 565346 255218 565582 255454
rect 565026 254898 565262 255134
rect 565346 254898 565582 255134
rect 565026 219218 565262 219454
rect 565346 219218 565582 219454
rect 565026 218898 565262 219134
rect 565346 218898 565582 219134
rect 565026 183218 565262 183454
rect 565346 183218 565582 183454
rect 565026 182898 565262 183134
rect 565346 182898 565582 183134
rect 565026 147218 565262 147454
rect 565346 147218 565582 147454
rect 565026 146898 565262 147134
rect 565346 146898 565582 147134
rect 565026 111218 565262 111454
rect 565346 111218 565582 111454
rect 565026 110898 565262 111134
rect 565346 110898 565582 111134
rect 565026 75218 565262 75454
rect 565346 75218 565582 75454
rect 565026 74898 565262 75134
rect 565346 74898 565582 75134
rect 565026 39218 565262 39454
rect 565346 39218 565582 39454
rect 565026 38898 565262 39134
rect 565346 38898 565582 39134
rect 565026 3218 565262 3454
rect 565346 3218 565582 3454
rect 565026 2898 565262 3134
rect 565346 2898 565582 3134
rect 565026 -582 565262 -346
rect 565346 -582 565582 -346
rect 565026 -902 565262 -666
rect 565346 -902 565582 -666
rect 571066 711322 571302 711558
rect 571386 711322 571622 711558
rect 571066 711002 571302 711238
rect 571386 711002 571622 711238
rect 565946 698378 566182 698614
rect 566266 698378 566502 698614
rect 565946 698058 566182 698294
rect 566266 698058 566502 698294
rect 565946 662378 566182 662614
rect 566266 662378 566502 662614
rect 565946 662058 566182 662294
rect 566266 662058 566502 662294
rect 565946 626378 566182 626614
rect 566266 626378 566502 626614
rect 565946 626058 566182 626294
rect 566266 626058 566502 626294
rect 565946 590378 566182 590614
rect 566266 590378 566502 590614
rect 565946 590058 566182 590294
rect 566266 590058 566502 590294
rect 565946 554378 566182 554614
rect 566266 554378 566502 554614
rect 565946 554058 566182 554294
rect 566266 554058 566502 554294
rect 565946 518378 566182 518614
rect 566266 518378 566502 518614
rect 565946 518058 566182 518294
rect 566266 518058 566502 518294
rect 565946 482378 566182 482614
rect 566266 482378 566502 482614
rect 565946 482058 566182 482294
rect 566266 482058 566502 482294
rect 565946 446378 566182 446614
rect 566266 446378 566502 446614
rect 565946 446058 566182 446294
rect 566266 446058 566502 446294
rect 565946 410378 566182 410614
rect 566266 410378 566502 410614
rect 565946 410058 566182 410294
rect 566266 410058 566502 410294
rect 565946 374378 566182 374614
rect 566266 374378 566502 374614
rect 565946 374058 566182 374294
rect 566266 374058 566502 374294
rect 565946 338378 566182 338614
rect 566266 338378 566502 338614
rect 565946 338058 566182 338294
rect 566266 338058 566502 338294
rect 565946 302378 566182 302614
rect 566266 302378 566502 302614
rect 565946 302058 566182 302294
rect 566266 302058 566502 302294
rect 565946 266378 566182 266614
rect 566266 266378 566502 266614
rect 565946 266058 566182 266294
rect 566266 266058 566502 266294
rect 565946 230378 566182 230614
rect 566266 230378 566502 230614
rect 565946 230058 566182 230294
rect 566266 230058 566502 230294
rect 565946 194378 566182 194614
rect 566266 194378 566502 194614
rect 565946 194058 566182 194294
rect 566266 194058 566502 194294
rect 565946 158378 566182 158614
rect 566266 158378 566502 158614
rect 565946 158058 566182 158294
rect 566266 158058 566502 158294
rect 565946 122378 566182 122614
rect 566266 122378 566502 122614
rect 565946 122058 566182 122294
rect 566266 122058 566502 122294
rect 565946 86378 566182 86614
rect 566266 86378 566502 86614
rect 565946 86058 566182 86294
rect 566266 86058 566502 86294
rect 565946 50378 566182 50614
rect 566266 50378 566502 50614
rect 565946 50058 566182 50294
rect 566266 50058 566502 50294
rect 565946 14378 566182 14614
rect 566266 14378 566502 14614
rect 565946 14058 566182 14294
rect 566266 14058 566502 14294
rect 563626 -3462 563862 -3226
rect 563946 -3462 564182 -3226
rect 563626 -3782 563862 -3546
rect 563946 -3782 564182 -3546
rect 562226 -4422 562462 -4186
rect 562546 -4422 562782 -4186
rect 562226 -4742 562462 -4506
rect 562546 -4742 562782 -4506
rect 560826 -7302 561062 -7066
rect 561146 -7302 561382 -7066
rect 560826 -7622 561062 -7386
rect 561146 -7622 561382 -7386
rect 567346 709402 567582 709638
rect 567666 709402 567902 709638
rect 567346 709082 567582 709318
rect 567666 709082 567902 709318
rect 567346 676658 567582 676894
rect 567666 676658 567902 676894
rect 567346 676338 567582 676574
rect 567666 676338 567902 676574
rect 567346 640658 567582 640894
rect 567666 640658 567902 640894
rect 567346 640338 567582 640574
rect 567666 640338 567902 640574
rect 567346 604658 567582 604894
rect 567666 604658 567902 604894
rect 567346 604338 567582 604574
rect 567666 604338 567902 604574
rect 567346 568658 567582 568894
rect 567666 568658 567902 568894
rect 567346 568338 567582 568574
rect 567666 568338 567902 568574
rect 567346 532658 567582 532894
rect 567666 532658 567902 532894
rect 567346 532338 567582 532574
rect 567666 532338 567902 532574
rect 567346 496658 567582 496894
rect 567666 496658 567902 496894
rect 567346 496338 567582 496574
rect 567666 496338 567902 496574
rect 567346 460658 567582 460894
rect 567666 460658 567902 460894
rect 567346 460338 567582 460574
rect 567666 460338 567902 460574
rect 567346 424658 567582 424894
rect 567666 424658 567902 424894
rect 567346 424338 567582 424574
rect 567666 424338 567902 424574
rect 567346 388658 567582 388894
rect 567666 388658 567902 388894
rect 567346 388338 567582 388574
rect 567666 388338 567902 388574
rect 567346 352658 567582 352894
rect 567666 352658 567902 352894
rect 567346 352338 567582 352574
rect 567666 352338 567902 352574
rect 567346 316658 567582 316894
rect 567666 316658 567902 316894
rect 567346 316338 567582 316574
rect 567666 316338 567902 316574
rect 567346 280658 567582 280894
rect 567666 280658 567902 280894
rect 567346 280338 567582 280574
rect 567666 280338 567902 280574
rect 567346 244658 567582 244894
rect 567666 244658 567902 244894
rect 567346 244338 567582 244574
rect 567666 244338 567902 244574
rect 567346 208658 567582 208894
rect 567666 208658 567902 208894
rect 567346 208338 567582 208574
rect 567666 208338 567902 208574
rect 567346 172658 567582 172894
rect 567666 172658 567902 172894
rect 567346 172338 567582 172574
rect 567666 172338 567902 172574
rect 567346 136658 567582 136894
rect 567666 136658 567902 136894
rect 567346 136338 567582 136574
rect 567666 136338 567902 136574
rect 567346 100658 567582 100894
rect 567666 100658 567902 100894
rect 567346 100338 567582 100574
rect 567666 100338 567902 100574
rect 567346 64658 567582 64894
rect 567666 64658 567902 64894
rect 567346 64338 567582 64574
rect 567666 64338 567902 64574
rect 567346 28658 567582 28894
rect 567666 28658 567902 28894
rect 567346 28338 567582 28574
rect 567666 28338 567902 28574
rect 568746 706522 568982 706758
rect 569066 706522 569302 706758
rect 568746 706202 568982 706438
rect 569066 706202 569302 706438
rect 568746 690938 568982 691174
rect 569066 690938 569302 691174
rect 568746 690618 568982 690854
rect 569066 690618 569302 690854
rect 568746 654938 568982 655174
rect 569066 654938 569302 655174
rect 568746 654618 568982 654854
rect 569066 654618 569302 654854
rect 568746 618938 568982 619174
rect 569066 618938 569302 619174
rect 568746 618618 568982 618854
rect 569066 618618 569302 618854
rect 568746 582938 568982 583174
rect 569066 582938 569302 583174
rect 568746 582618 568982 582854
rect 569066 582618 569302 582854
rect 568746 546938 568982 547174
rect 569066 546938 569302 547174
rect 568746 546618 568982 546854
rect 569066 546618 569302 546854
rect 568746 510938 568982 511174
rect 569066 510938 569302 511174
rect 568746 510618 568982 510854
rect 569066 510618 569302 510854
rect 568746 474938 568982 475174
rect 569066 474938 569302 475174
rect 568746 474618 568982 474854
rect 569066 474618 569302 474854
rect 568746 438938 568982 439174
rect 569066 438938 569302 439174
rect 568746 438618 568982 438854
rect 569066 438618 569302 438854
rect 568746 402938 568982 403174
rect 569066 402938 569302 403174
rect 568746 402618 568982 402854
rect 569066 402618 569302 402854
rect 568746 366938 568982 367174
rect 569066 366938 569302 367174
rect 568746 366618 568982 366854
rect 569066 366618 569302 366854
rect 568746 330938 568982 331174
rect 569066 330938 569302 331174
rect 568746 330618 568982 330854
rect 569066 330618 569302 330854
rect 568746 294938 568982 295174
rect 569066 294938 569302 295174
rect 568746 294618 568982 294854
rect 569066 294618 569302 294854
rect 568746 258938 568982 259174
rect 569066 258938 569302 259174
rect 568746 258618 568982 258854
rect 569066 258618 569302 258854
rect 568746 222938 568982 223174
rect 569066 222938 569302 223174
rect 568746 222618 568982 222854
rect 569066 222618 569302 222854
rect 568746 186938 568982 187174
rect 569066 186938 569302 187174
rect 568746 186618 568982 186854
rect 569066 186618 569302 186854
rect 568746 150938 568982 151174
rect 569066 150938 569302 151174
rect 568746 150618 568982 150854
rect 569066 150618 569302 150854
rect 568746 114938 568982 115174
rect 569066 114938 569302 115174
rect 568746 114618 568982 114854
rect 569066 114618 569302 114854
rect 568746 78938 568982 79174
rect 569066 78938 569302 79174
rect 568746 78618 568982 78854
rect 569066 78618 569302 78854
rect 568746 42938 568982 43174
rect 569066 42938 569302 43174
rect 568746 42618 568982 42854
rect 569066 42618 569302 42854
rect 568746 6938 568982 7174
rect 569066 6938 569302 7174
rect 568746 6618 568982 6854
rect 569066 6618 569302 6854
rect 570146 705562 570382 705798
rect 570466 705562 570702 705798
rect 570146 705242 570382 705478
rect 570466 705242 570702 705478
rect 570146 669218 570382 669454
rect 570466 669218 570702 669454
rect 570146 668898 570382 669134
rect 570466 668898 570702 669134
rect 570146 633218 570382 633454
rect 570466 633218 570702 633454
rect 570146 632898 570382 633134
rect 570466 632898 570702 633134
rect 570146 597218 570382 597454
rect 570466 597218 570702 597454
rect 570146 596898 570382 597134
rect 570466 596898 570702 597134
rect 570146 561218 570382 561454
rect 570466 561218 570702 561454
rect 570146 560898 570382 561134
rect 570466 560898 570702 561134
rect 570146 525218 570382 525454
rect 570466 525218 570702 525454
rect 570146 524898 570382 525134
rect 570466 524898 570702 525134
rect 570146 489218 570382 489454
rect 570466 489218 570702 489454
rect 570146 488898 570382 489134
rect 570466 488898 570702 489134
rect 570146 453218 570382 453454
rect 570466 453218 570702 453454
rect 570146 452898 570382 453134
rect 570466 452898 570702 453134
rect 570146 417218 570382 417454
rect 570466 417218 570702 417454
rect 570146 416898 570382 417134
rect 570466 416898 570702 417134
rect 570146 381218 570382 381454
rect 570466 381218 570702 381454
rect 570146 380898 570382 381134
rect 570466 380898 570702 381134
rect 570146 345218 570382 345454
rect 570466 345218 570702 345454
rect 570146 344898 570382 345134
rect 570466 344898 570702 345134
rect 570146 309218 570382 309454
rect 570466 309218 570702 309454
rect 570146 308898 570382 309134
rect 570466 308898 570702 309134
rect 570146 273218 570382 273454
rect 570466 273218 570702 273454
rect 570146 272898 570382 273134
rect 570466 272898 570702 273134
rect 570146 237218 570382 237454
rect 570466 237218 570702 237454
rect 570146 236898 570382 237134
rect 570466 236898 570702 237134
rect 570146 201218 570382 201454
rect 570466 201218 570702 201454
rect 570146 200898 570382 201134
rect 570466 200898 570702 201134
rect 570146 165218 570382 165454
rect 570466 165218 570702 165454
rect 570146 164898 570382 165134
rect 570466 164898 570702 165134
rect 570146 129218 570382 129454
rect 570466 129218 570702 129454
rect 570146 128898 570382 129134
rect 570466 128898 570702 129134
rect 570146 93218 570382 93454
rect 570466 93218 570702 93454
rect 570146 92898 570382 93134
rect 570466 92898 570702 93134
rect 570146 57218 570382 57454
rect 570466 57218 570702 57454
rect 570146 56898 570382 57134
rect 570466 56898 570702 57134
rect 570146 21218 570382 21454
rect 570466 21218 570702 21454
rect 570146 20898 570382 21134
rect 570466 20898 570702 21134
rect 570146 -1542 570382 -1306
rect 570466 -1542 570702 -1306
rect 570146 -1862 570382 -1626
rect 570466 -1862 570702 -1626
rect 576186 710362 576422 710598
rect 576506 710362 576742 710598
rect 576186 710042 576422 710278
rect 576506 710042 576742 710278
rect 571066 680378 571302 680614
rect 571386 680378 571622 680614
rect 571066 680058 571302 680294
rect 571386 680058 571622 680294
rect 571066 644378 571302 644614
rect 571386 644378 571622 644614
rect 571066 644058 571302 644294
rect 571386 644058 571622 644294
rect 571066 608378 571302 608614
rect 571386 608378 571622 608614
rect 571066 608058 571302 608294
rect 571386 608058 571622 608294
rect 571066 572378 571302 572614
rect 571386 572378 571622 572614
rect 571066 572058 571302 572294
rect 571386 572058 571622 572294
rect 571066 536378 571302 536614
rect 571386 536378 571622 536614
rect 571066 536058 571302 536294
rect 571386 536058 571622 536294
rect 571066 500378 571302 500614
rect 571386 500378 571622 500614
rect 571066 500058 571302 500294
rect 571386 500058 571622 500294
rect 571066 464378 571302 464614
rect 571386 464378 571622 464614
rect 571066 464058 571302 464294
rect 571386 464058 571622 464294
rect 571066 428378 571302 428614
rect 571386 428378 571622 428614
rect 571066 428058 571302 428294
rect 571386 428058 571622 428294
rect 571066 392378 571302 392614
rect 571386 392378 571622 392614
rect 571066 392058 571302 392294
rect 571386 392058 571622 392294
rect 571066 356378 571302 356614
rect 571386 356378 571622 356614
rect 571066 356058 571302 356294
rect 571386 356058 571622 356294
rect 571066 320378 571302 320614
rect 571386 320378 571622 320614
rect 571066 320058 571302 320294
rect 571386 320058 571622 320294
rect 571066 284378 571302 284614
rect 571386 284378 571622 284614
rect 571066 284058 571302 284294
rect 571386 284058 571622 284294
rect 571066 248378 571302 248614
rect 571386 248378 571622 248614
rect 571066 248058 571302 248294
rect 571386 248058 571622 248294
rect 571066 212378 571302 212614
rect 571386 212378 571622 212614
rect 571066 212058 571302 212294
rect 571386 212058 571622 212294
rect 571066 176378 571302 176614
rect 571386 176378 571622 176614
rect 571066 176058 571302 176294
rect 571386 176058 571622 176294
rect 571066 140378 571302 140614
rect 571386 140378 571622 140614
rect 571066 140058 571302 140294
rect 571386 140058 571622 140294
rect 571066 104378 571302 104614
rect 571386 104378 571622 104614
rect 571066 104058 571302 104294
rect 571386 104058 571622 104294
rect 571066 68378 571302 68614
rect 571386 68378 571622 68614
rect 571066 68058 571302 68294
rect 571386 68058 571622 68294
rect 571066 32378 571302 32614
rect 571386 32378 571622 32614
rect 571066 32058 571302 32294
rect 571386 32058 571622 32294
rect 568746 -2502 568982 -2266
rect 569066 -2502 569302 -2266
rect 568746 -2822 568982 -2586
rect 569066 -2822 569302 -2586
rect 567346 -5382 567582 -5146
rect 567666 -5382 567902 -5146
rect 567346 -5702 567582 -5466
rect 567666 -5702 567902 -5466
rect 565946 -6342 566182 -6106
rect 566266 -6342 566502 -6106
rect 565946 -6662 566182 -6426
rect 566266 -6662 566502 -6426
rect 572466 708442 572702 708678
rect 572786 708442 573022 708678
rect 572466 708122 572702 708358
rect 572786 708122 573022 708358
rect 572466 694658 572702 694894
rect 572786 694658 573022 694894
rect 572466 694338 572702 694574
rect 572786 694338 573022 694574
rect 572466 658658 572702 658894
rect 572786 658658 573022 658894
rect 572466 658338 572702 658574
rect 572786 658338 573022 658574
rect 572466 622658 572702 622894
rect 572786 622658 573022 622894
rect 572466 622338 572702 622574
rect 572786 622338 573022 622574
rect 572466 586658 572702 586894
rect 572786 586658 573022 586894
rect 572466 586338 572702 586574
rect 572786 586338 573022 586574
rect 572466 550658 572702 550894
rect 572786 550658 573022 550894
rect 572466 550338 572702 550574
rect 572786 550338 573022 550574
rect 572466 514658 572702 514894
rect 572786 514658 573022 514894
rect 572466 514338 572702 514574
rect 572786 514338 573022 514574
rect 572466 478658 572702 478894
rect 572786 478658 573022 478894
rect 572466 478338 572702 478574
rect 572786 478338 573022 478574
rect 572466 442658 572702 442894
rect 572786 442658 573022 442894
rect 572466 442338 572702 442574
rect 572786 442338 573022 442574
rect 572466 406658 572702 406894
rect 572786 406658 573022 406894
rect 572466 406338 572702 406574
rect 572786 406338 573022 406574
rect 572466 370658 572702 370894
rect 572786 370658 573022 370894
rect 572466 370338 572702 370574
rect 572786 370338 573022 370574
rect 572466 334658 572702 334894
rect 572786 334658 573022 334894
rect 572466 334338 572702 334574
rect 572786 334338 573022 334574
rect 572466 298658 572702 298894
rect 572786 298658 573022 298894
rect 572466 298338 572702 298574
rect 572786 298338 573022 298574
rect 572466 262658 572702 262894
rect 572786 262658 573022 262894
rect 572466 262338 572702 262574
rect 572786 262338 573022 262574
rect 572466 226658 572702 226894
rect 572786 226658 573022 226894
rect 572466 226338 572702 226574
rect 572786 226338 573022 226574
rect 572466 190658 572702 190894
rect 572786 190658 573022 190894
rect 572466 190338 572702 190574
rect 572786 190338 573022 190574
rect 572466 154658 572702 154894
rect 572786 154658 573022 154894
rect 572466 154338 572702 154574
rect 572786 154338 573022 154574
rect 572466 118658 572702 118894
rect 572786 118658 573022 118894
rect 572466 118338 572702 118574
rect 572786 118338 573022 118574
rect 572466 82658 572702 82894
rect 572786 82658 573022 82894
rect 572466 82338 572702 82574
rect 572786 82338 573022 82574
rect 572466 46658 572702 46894
rect 572786 46658 573022 46894
rect 572466 46338 572702 46574
rect 572786 46338 573022 46574
rect 572466 10658 572702 10894
rect 572786 10658 573022 10894
rect 572466 10338 572702 10574
rect 572786 10338 573022 10574
rect 573866 707482 574102 707718
rect 574186 707482 574422 707718
rect 573866 707162 574102 707398
rect 574186 707162 574422 707398
rect 573866 672938 574102 673174
rect 574186 672938 574422 673174
rect 573866 672618 574102 672854
rect 574186 672618 574422 672854
rect 573866 636938 574102 637174
rect 574186 636938 574422 637174
rect 573866 636618 574102 636854
rect 574186 636618 574422 636854
rect 573866 600938 574102 601174
rect 574186 600938 574422 601174
rect 573866 600618 574102 600854
rect 574186 600618 574422 600854
rect 573866 564938 574102 565174
rect 574186 564938 574422 565174
rect 573866 564618 574102 564854
rect 574186 564618 574422 564854
rect 573866 528938 574102 529174
rect 574186 528938 574422 529174
rect 573866 528618 574102 528854
rect 574186 528618 574422 528854
rect 573866 492938 574102 493174
rect 574186 492938 574422 493174
rect 573866 492618 574102 492854
rect 574186 492618 574422 492854
rect 573866 456938 574102 457174
rect 574186 456938 574422 457174
rect 573866 456618 574102 456854
rect 574186 456618 574422 456854
rect 573866 420938 574102 421174
rect 574186 420938 574422 421174
rect 573866 420618 574102 420854
rect 574186 420618 574422 420854
rect 573866 384938 574102 385174
rect 574186 384938 574422 385174
rect 573866 384618 574102 384854
rect 574186 384618 574422 384854
rect 573866 348938 574102 349174
rect 574186 348938 574422 349174
rect 573866 348618 574102 348854
rect 574186 348618 574422 348854
rect 573866 312938 574102 313174
rect 574186 312938 574422 313174
rect 573866 312618 574102 312854
rect 574186 312618 574422 312854
rect 573866 276938 574102 277174
rect 574186 276938 574422 277174
rect 573866 276618 574102 276854
rect 574186 276618 574422 276854
rect 573866 240938 574102 241174
rect 574186 240938 574422 241174
rect 573866 240618 574102 240854
rect 574186 240618 574422 240854
rect 573866 204938 574102 205174
rect 574186 204938 574422 205174
rect 573866 204618 574102 204854
rect 574186 204618 574422 204854
rect 573866 168938 574102 169174
rect 574186 168938 574422 169174
rect 573866 168618 574102 168854
rect 574186 168618 574422 168854
rect 573866 132938 574102 133174
rect 574186 132938 574422 133174
rect 573866 132618 574102 132854
rect 574186 132618 574422 132854
rect 573866 96938 574102 97174
rect 574186 96938 574422 97174
rect 573866 96618 574102 96854
rect 574186 96618 574422 96854
rect 573866 60938 574102 61174
rect 574186 60938 574422 61174
rect 573866 60618 574102 60854
rect 574186 60618 574422 60854
rect 573866 24938 574102 25174
rect 574186 24938 574422 25174
rect 573866 24618 574102 24854
rect 574186 24618 574422 24854
rect 575266 704602 575502 704838
rect 575586 704602 575822 704838
rect 575266 704282 575502 704518
rect 575586 704282 575822 704518
rect 575266 687218 575502 687454
rect 575586 687218 575822 687454
rect 575266 686898 575502 687134
rect 575586 686898 575822 687134
rect 575266 651218 575502 651454
rect 575586 651218 575822 651454
rect 575266 650898 575502 651134
rect 575586 650898 575822 651134
rect 575266 615218 575502 615454
rect 575586 615218 575822 615454
rect 575266 614898 575502 615134
rect 575586 614898 575822 615134
rect 575266 579218 575502 579454
rect 575586 579218 575822 579454
rect 575266 578898 575502 579134
rect 575586 578898 575822 579134
rect 575266 543218 575502 543454
rect 575586 543218 575822 543454
rect 575266 542898 575502 543134
rect 575586 542898 575822 543134
rect 575266 507218 575502 507454
rect 575586 507218 575822 507454
rect 575266 506898 575502 507134
rect 575586 506898 575822 507134
rect 575266 471218 575502 471454
rect 575586 471218 575822 471454
rect 575266 470898 575502 471134
rect 575586 470898 575822 471134
rect 575266 435218 575502 435454
rect 575586 435218 575822 435454
rect 575266 434898 575502 435134
rect 575586 434898 575822 435134
rect 575266 399218 575502 399454
rect 575586 399218 575822 399454
rect 575266 398898 575502 399134
rect 575586 398898 575822 399134
rect 575266 363218 575502 363454
rect 575586 363218 575822 363454
rect 575266 362898 575502 363134
rect 575586 362898 575822 363134
rect 575266 327218 575502 327454
rect 575586 327218 575822 327454
rect 575266 326898 575502 327134
rect 575586 326898 575822 327134
rect 575266 291218 575502 291454
rect 575586 291218 575822 291454
rect 575266 290898 575502 291134
rect 575586 290898 575822 291134
rect 575266 255218 575502 255454
rect 575586 255218 575822 255454
rect 575266 254898 575502 255134
rect 575586 254898 575822 255134
rect 575266 219218 575502 219454
rect 575586 219218 575822 219454
rect 575266 218898 575502 219134
rect 575586 218898 575822 219134
rect 575266 183218 575502 183454
rect 575586 183218 575822 183454
rect 575266 182898 575502 183134
rect 575586 182898 575822 183134
rect 575266 147218 575502 147454
rect 575586 147218 575822 147454
rect 575266 146898 575502 147134
rect 575586 146898 575822 147134
rect 575266 111218 575502 111454
rect 575586 111218 575822 111454
rect 575266 110898 575502 111134
rect 575586 110898 575822 111134
rect 575266 75218 575502 75454
rect 575586 75218 575822 75454
rect 575266 74898 575502 75134
rect 575586 74898 575822 75134
rect 575266 39218 575502 39454
rect 575586 39218 575822 39454
rect 575266 38898 575502 39134
rect 575586 38898 575822 39134
rect 575266 3218 575502 3454
rect 575586 3218 575822 3454
rect 575266 2898 575502 3134
rect 575586 2898 575822 3134
rect 575266 -582 575502 -346
rect 575586 -582 575822 -346
rect 575266 -902 575502 -666
rect 575586 -902 575822 -666
rect 581306 711322 581542 711558
rect 581626 711322 581862 711558
rect 581306 711002 581542 711238
rect 581626 711002 581862 711238
rect 576186 698378 576422 698614
rect 576506 698378 576742 698614
rect 576186 698058 576422 698294
rect 576506 698058 576742 698294
rect 576186 662378 576422 662614
rect 576506 662378 576742 662614
rect 576186 662058 576422 662294
rect 576506 662058 576742 662294
rect 576186 626378 576422 626614
rect 576506 626378 576742 626614
rect 576186 626058 576422 626294
rect 576506 626058 576742 626294
rect 576186 590378 576422 590614
rect 576506 590378 576742 590614
rect 576186 590058 576422 590294
rect 576506 590058 576742 590294
rect 576186 554378 576422 554614
rect 576506 554378 576742 554614
rect 576186 554058 576422 554294
rect 576506 554058 576742 554294
rect 576186 518378 576422 518614
rect 576506 518378 576742 518614
rect 576186 518058 576422 518294
rect 576506 518058 576742 518294
rect 576186 482378 576422 482614
rect 576506 482378 576742 482614
rect 576186 482058 576422 482294
rect 576506 482058 576742 482294
rect 576186 446378 576422 446614
rect 576506 446378 576742 446614
rect 576186 446058 576422 446294
rect 576506 446058 576742 446294
rect 576186 410378 576422 410614
rect 576506 410378 576742 410614
rect 576186 410058 576422 410294
rect 576506 410058 576742 410294
rect 576186 374378 576422 374614
rect 576506 374378 576742 374614
rect 576186 374058 576422 374294
rect 576506 374058 576742 374294
rect 576186 338378 576422 338614
rect 576506 338378 576742 338614
rect 576186 338058 576422 338294
rect 576506 338058 576742 338294
rect 576186 302378 576422 302614
rect 576506 302378 576742 302614
rect 576186 302058 576422 302294
rect 576506 302058 576742 302294
rect 576186 266378 576422 266614
rect 576506 266378 576742 266614
rect 576186 266058 576422 266294
rect 576506 266058 576742 266294
rect 576186 230378 576422 230614
rect 576506 230378 576742 230614
rect 576186 230058 576422 230294
rect 576506 230058 576742 230294
rect 576186 194378 576422 194614
rect 576506 194378 576742 194614
rect 576186 194058 576422 194294
rect 576506 194058 576742 194294
rect 576186 158378 576422 158614
rect 576506 158378 576742 158614
rect 576186 158058 576422 158294
rect 576506 158058 576742 158294
rect 576186 122378 576422 122614
rect 576506 122378 576742 122614
rect 576186 122058 576422 122294
rect 576506 122058 576742 122294
rect 576186 86378 576422 86614
rect 576506 86378 576742 86614
rect 576186 86058 576422 86294
rect 576506 86058 576742 86294
rect 576186 50378 576422 50614
rect 576506 50378 576742 50614
rect 576186 50058 576422 50294
rect 576506 50058 576742 50294
rect 576186 14378 576422 14614
rect 576506 14378 576742 14614
rect 576186 14058 576422 14294
rect 576506 14058 576742 14294
rect 573866 -3462 574102 -3226
rect 574186 -3462 574422 -3226
rect 573866 -3782 574102 -3546
rect 574186 -3782 574422 -3546
rect 572466 -4422 572702 -4186
rect 572786 -4422 573022 -4186
rect 572466 -4742 572702 -4506
rect 572786 -4742 573022 -4506
rect 571066 -7302 571302 -7066
rect 571386 -7302 571622 -7066
rect 571066 -7622 571302 -7386
rect 571386 -7622 571622 -7386
rect 577586 709402 577822 709638
rect 577906 709402 578142 709638
rect 577586 709082 577822 709318
rect 577906 709082 578142 709318
rect 577586 676658 577822 676894
rect 577906 676658 578142 676894
rect 577586 676338 577822 676574
rect 577906 676338 578142 676574
rect 577586 640658 577822 640894
rect 577906 640658 578142 640894
rect 577586 640338 577822 640574
rect 577906 640338 578142 640574
rect 577586 604658 577822 604894
rect 577906 604658 578142 604894
rect 577586 604338 577822 604574
rect 577906 604338 578142 604574
rect 577586 568658 577822 568894
rect 577906 568658 578142 568894
rect 577586 568338 577822 568574
rect 577906 568338 578142 568574
rect 577586 532658 577822 532894
rect 577906 532658 578142 532894
rect 577586 532338 577822 532574
rect 577906 532338 578142 532574
rect 577586 496658 577822 496894
rect 577906 496658 578142 496894
rect 577586 496338 577822 496574
rect 577906 496338 578142 496574
rect 577586 460658 577822 460894
rect 577906 460658 578142 460894
rect 577586 460338 577822 460574
rect 577906 460338 578142 460574
rect 577586 424658 577822 424894
rect 577906 424658 578142 424894
rect 577586 424338 577822 424574
rect 577906 424338 578142 424574
rect 577586 388658 577822 388894
rect 577906 388658 578142 388894
rect 577586 388338 577822 388574
rect 577906 388338 578142 388574
rect 577586 352658 577822 352894
rect 577906 352658 578142 352894
rect 577586 352338 577822 352574
rect 577906 352338 578142 352574
rect 577586 316658 577822 316894
rect 577906 316658 578142 316894
rect 577586 316338 577822 316574
rect 577906 316338 578142 316574
rect 577586 280658 577822 280894
rect 577906 280658 578142 280894
rect 577586 280338 577822 280574
rect 577906 280338 578142 280574
rect 577586 244658 577822 244894
rect 577906 244658 578142 244894
rect 577586 244338 577822 244574
rect 577906 244338 578142 244574
rect 577586 208658 577822 208894
rect 577906 208658 578142 208894
rect 577586 208338 577822 208574
rect 577906 208338 578142 208574
rect 577586 172658 577822 172894
rect 577906 172658 578142 172894
rect 577586 172338 577822 172574
rect 577906 172338 578142 172574
rect 577586 136658 577822 136894
rect 577906 136658 578142 136894
rect 577586 136338 577822 136574
rect 577906 136338 578142 136574
rect 577586 100658 577822 100894
rect 577906 100658 578142 100894
rect 577586 100338 577822 100574
rect 577906 100338 578142 100574
rect 577586 64658 577822 64894
rect 577906 64658 578142 64894
rect 577586 64338 577822 64574
rect 577906 64338 578142 64574
rect 577586 28658 577822 28894
rect 577906 28658 578142 28894
rect 577586 28338 577822 28574
rect 577906 28338 578142 28574
rect 578986 706522 579222 706758
rect 579306 706522 579542 706758
rect 578986 706202 579222 706438
rect 579306 706202 579542 706438
rect 578986 690938 579222 691174
rect 579306 690938 579542 691174
rect 578986 690618 579222 690854
rect 579306 690618 579542 690854
rect 578986 654938 579222 655174
rect 579306 654938 579542 655174
rect 578986 654618 579222 654854
rect 579306 654618 579542 654854
rect 578986 618938 579222 619174
rect 579306 618938 579542 619174
rect 578986 618618 579222 618854
rect 579306 618618 579542 618854
rect 578986 582938 579222 583174
rect 579306 582938 579542 583174
rect 578986 582618 579222 582854
rect 579306 582618 579542 582854
rect 578986 546938 579222 547174
rect 579306 546938 579542 547174
rect 578986 546618 579222 546854
rect 579306 546618 579542 546854
rect 578986 510938 579222 511174
rect 579306 510938 579542 511174
rect 578986 510618 579222 510854
rect 579306 510618 579542 510854
rect 578986 474938 579222 475174
rect 579306 474938 579542 475174
rect 578986 474618 579222 474854
rect 579306 474618 579542 474854
rect 578986 438938 579222 439174
rect 579306 438938 579542 439174
rect 578986 438618 579222 438854
rect 579306 438618 579542 438854
rect 578986 402938 579222 403174
rect 579306 402938 579542 403174
rect 578986 402618 579222 402854
rect 579306 402618 579542 402854
rect 578986 366938 579222 367174
rect 579306 366938 579542 367174
rect 578986 366618 579222 366854
rect 579306 366618 579542 366854
rect 578986 330938 579222 331174
rect 579306 330938 579542 331174
rect 578986 330618 579222 330854
rect 579306 330618 579542 330854
rect 578986 294938 579222 295174
rect 579306 294938 579542 295174
rect 578986 294618 579222 294854
rect 579306 294618 579542 294854
rect 578986 258938 579222 259174
rect 579306 258938 579542 259174
rect 578986 258618 579222 258854
rect 579306 258618 579542 258854
rect 578986 222938 579222 223174
rect 579306 222938 579542 223174
rect 578986 222618 579222 222854
rect 579306 222618 579542 222854
rect 578986 186938 579222 187174
rect 579306 186938 579542 187174
rect 578986 186618 579222 186854
rect 579306 186618 579542 186854
rect 578986 150938 579222 151174
rect 579306 150938 579542 151174
rect 578986 150618 579222 150854
rect 579306 150618 579542 150854
rect 578986 114938 579222 115174
rect 579306 114938 579542 115174
rect 578986 114618 579222 114854
rect 579306 114618 579542 114854
rect 578986 78938 579222 79174
rect 579306 78938 579542 79174
rect 578986 78618 579222 78854
rect 579306 78618 579542 78854
rect 578986 42938 579222 43174
rect 579306 42938 579542 43174
rect 578986 42618 579222 42854
rect 579306 42618 579542 42854
rect 578986 6938 579222 7174
rect 579306 6938 579542 7174
rect 578986 6618 579222 6854
rect 579306 6618 579542 6854
rect 580386 705562 580622 705798
rect 580706 705562 580942 705798
rect 580386 705242 580622 705478
rect 580706 705242 580942 705478
rect 580386 669218 580622 669454
rect 580706 669218 580942 669454
rect 580386 668898 580622 669134
rect 580706 668898 580942 669134
rect 580386 633218 580622 633454
rect 580706 633218 580942 633454
rect 580386 632898 580622 633134
rect 580706 632898 580942 633134
rect 580386 597218 580622 597454
rect 580706 597218 580942 597454
rect 580386 596898 580622 597134
rect 580706 596898 580942 597134
rect 580386 561218 580622 561454
rect 580706 561218 580942 561454
rect 580386 560898 580622 561134
rect 580706 560898 580942 561134
rect 580386 525218 580622 525454
rect 580706 525218 580942 525454
rect 580386 524898 580622 525134
rect 580706 524898 580942 525134
rect 580386 489218 580622 489454
rect 580706 489218 580942 489454
rect 580386 488898 580622 489134
rect 580706 488898 580942 489134
rect 580386 453218 580622 453454
rect 580706 453218 580942 453454
rect 580386 452898 580622 453134
rect 580706 452898 580942 453134
rect 580386 417218 580622 417454
rect 580706 417218 580942 417454
rect 580386 416898 580622 417134
rect 580706 416898 580942 417134
rect 580386 381218 580622 381454
rect 580706 381218 580942 381454
rect 580386 380898 580622 381134
rect 580706 380898 580942 381134
rect 580386 345218 580622 345454
rect 580706 345218 580942 345454
rect 580386 344898 580622 345134
rect 580706 344898 580942 345134
rect 580386 309218 580622 309454
rect 580706 309218 580942 309454
rect 580386 308898 580622 309134
rect 580706 308898 580942 309134
rect 580386 273218 580622 273454
rect 580706 273218 580942 273454
rect 580386 272898 580622 273134
rect 580706 272898 580942 273134
rect 580386 237218 580622 237454
rect 580706 237218 580942 237454
rect 580386 236898 580622 237134
rect 580706 236898 580942 237134
rect 580386 201218 580622 201454
rect 580706 201218 580942 201454
rect 580386 200898 580622 201134
rect 580706 200898 580942 201134
rect 580386 165218 580622 165454
rect 580706 165218 580942 165454
rect 580386 164898 580622 165134
rect 580706 164898 580942 165134
rect 580386 129218 580622 129454
rect 580706 129218 580942 129454
rect 580386 128898 580622 129134
rect 580706 128898 580942 129134
rect 580386 93218 580622 93454
rect 580706 93218 580942 93454
rect 580386 92898 580622 93134
rect 580706 92898 580942 93134
rect 580386 57218 580622 57454
rect 580706 57218 580942 57454
rect 580386 56898 580622 57134
rect 580706 56898 580942 57134
rect 580386 21218 580622 21454
rect 580706 21218 580942 21454
rect 580386 20898 580622 21134
rect 580706 20898 580942 21134
rect 580386 -1542 580622 -1306
rect 580706 -1542 580942 -1306
rect 580386 -1862 580622 -1626
rect 580706 -1862 580942 -1626
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581306 680378 581542 680614
rect 581626 680378 581862 680614
rect 581306 680058 581542 680294
rect 581626 680058 581862 680294
rect 581306 644378 581542 644614
rect 581626 644378 581862 644614
rect 581306 644058 581542 644294
rect 581626 644058 581862 644294
rect 581306 608378 581542 608614
rect 581626 608378 581862 608614
rect 581306 608058 581542 608294
rect 581626 608058 581862 608294
rect 581306 572378 581542 572614
rect 581626 572378 581862 572614
rect 581306 572058 581542 572294
rect 581626 572058 581862 572294
rect 581306 536378 581542 536614
rect 581626 536378 581862 536614
rect 581306 536058 581542 536294
rect 581626 536058 581862 536294
rect 581306 500378 581542 500614
rect 581626 500378 581862 500614
rect 581306 500058 581542 500294
rect 581626 500058 581862 500294
rect 581306 464378 581542 464614
rect 581626 464378 581862 464614
rect 581306 464058 581542 464294
rect 581626 464058 581862 464294
rect 581306 428378 581542 428614
rect 581626 428378 581862 428614
rect 581306 428058 581542 428294
rect 581626 428058 581862 428294
rect 581306 392378 581542 392614
rect 581626 392378 581862 392614
rect 581306 392058 581542 392294
rect 581626 392058 581862 392294
rect 581306 356378 581542 356614
rect 581626 356378 581862 356614
rect 581306 356058 581542 356294
rect 581626 356058 581862 356294
rect 581306 320378 581542 320614
rect 581626 320378 581862 320614
rect 581306 320058 581542 320294
rect 581626 320058 581862 320294
rect 581306 284378 581542 284614
rect 581626 284378 581862 284614
rect 581306 284058 581542 284294
rect 581626 284058 581862 284294
rect 581306 248378 581542 248614
rect 581626 248378 581862 248614
rect 581306 248058 581542 248294
rect 581626 248058 581862 248294
rect 581306 212378 581542 212614
rect 581626 212378 581862 212614
rect 581306 212058 581542 212294
rect 581626 212058 581862 212294
rect 581306 176378 581542 176614
rect 581626 176378 581862 176614
rect 581306 176058 581542 176294
rect 581626 176058 581862 176294
rect 581306 140378 581542 140614
rect 581626 140378 581862 140614
rect 581306 140058 581542 140294
rect 581626 140058 581862 140294
rect 581306 104378 581542 104614
rect 581626 104378 581862 104614
rect 581306 104058 581542 104294
rect 581626 104058 581862 104294
rect 581306 68378 581542 68614
rect 581626 68378 581862 68614
rect 581306 68058 581542 68294
rect 581626 68058 581862 68294
rect 581306 32378 581542 32614
rect 581626 32378 581862 32614
rect 581306 32058 581542 32294
rect 581626 32058 581862 32294
rect 578986 -2502 579222 -2266
rect 579306 -2502 579542 -2266
rect 578986 -2822 579222 -2586
rect 579306 -2822 579542 -2586
rect 577586 -5382 577822 -5146
rect 577906 -5382 578142 -5146
rect 577586 -5702 577822 -5466
rect 577906 -5702 578142 -5466
rect 576186 -6342 576422 -6106
rect 576506 -6342 576742 -6106
rect 576186 -6662 576422 -6426
rect 576506 -6662 576742 -6426
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 581306 -7302 581542 -7066
rect 581626 -7302 581862 -7066
rect 581306 -7622 581542 -7386
rect 581626 -7622 581862 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 18106 711558
rect 18342 711322 18426 711558
rect 18662 711322 28346 711558
rect 28582 711322 28666 711558
rect 28902 711322 38586 711558
rect 38822 711322 38906 711558
rect 39142 711322 48826 711558
rect 49062 711322 49146 711558
rect 49382 711322 59066 711558
rect 59302 711322 59386 711558
rect 59622 711322 69306 711558
rect 69542 711322 69626 711558
rect 69862 711322 79546 711558
rect 79782 711322 79866 711558
rect 80102 711322 89786 711558
rect 90022 711322 90106 711558
rect 90342 711322 100026 711558
rect 100262 711322 100346 711558
rect 100582 711322 110266 711558
rect 110502 711322 110586 711558
rect 110822 711322 120506 711558
rect 120742 711322 120826 711558
rect 121062 711322 130746 711558
rect 130982 711322 131066 711558
rect 131302 711322 140986 711558
rect 141222 711322 141306 711558
rect 141542 711322 151226 711558
rect 151462 711322 151546 711558
rect 151782 711322 161466 711558
rect 161702 711322 161786 711558
rect 162022 711322 171706 711558
rect 171942 711322 172026 711558
rect 172262 711322 181946 711558
rect 182182 711322 182266 711558
rect 182502 711322 192186 711558
rect 192422 711322 192506 711558
rect 192742 711322 202426 711558
rect 202662 711322 202746 711558
rect 202982 711322 212666 711558
rect 212902 711322 212986 711558
rect 213222 711322 222906 711558
rect 223142 711322 223226 711558
rect 223462 711322 233146 711558
rect 233382 711322 233466 711558
rect 233702 711322 243386 711558
rect 243622 711322 243706 711558
rect 243942 711322 253626 711558
rect 253862 711322 253946 711558
rect 254182 711322 263866 711558
rect 264102 711322 264186 711558
rect 264422 711322 274106 711558
rect 274342 711322 274426 711558
rect 274662 711322 284346 711558
rect 284582 711322 284666 711558
rect 284902 711322 294586 711558
rect 294822 711322 294906 711558
rect 295142 711322 304826 711558
rect 305062 711322 305146 711558
rect 305382 711322 315066 711558
rect 315302 711322 315386 711558
rect 315622 711322 325306 711558
rect 325542 711322 325626 711558
rect 325862 711322 335546 711558
rect 335782 711322 335866 711558
rect 336102 711322 345786 711558
rect 346022 711322 346106 711558
rect 346342 711322 356026 711558
rect 356262 711322 356346 711558
rect 356582 711322 366266 711558
rect 366502 711322 366586 711558
rect 366822 711322 376506 711558
rect 376742 711322 376826 711558
rect 377062 711322 386746 711558
rect 386982 711322 387066 711558
rect 387302 711322 396986 711558
rect 397222 711322 397306 711558
rect 397542 711322 407226 711558
rect 407462 711322 407546 711558
rect 407782 711322 417466 711558
rect 417702 711322 417786 711558
rect 418022 711322 427706 711558
rect 427942 711322 428026 711558
rect 428262 711322 437946 711558
rect 438182 711322 438266 711558
rect 438502 711322 448186 711558
rect 448422 711322 448506 711558
rect 448742 711322 458426 711558
rect 458662 711322 458746 711558
rect 458982 711322 468666 711558
rect 468902 711322 468986 711558
rect 469222 711322 478906 711558
rect 479142 711322 479226 711558
rect 479462 711322 489146 711558
rect 489382 711322 489466 711558
rect 489702 711322 499386 711558
rect 499622 711322 499706 711558
rect 499942 711322 509626 711558
rect 509862 711322 509946 711558
rect 510182 711322 519866 711558
rect 520102 711322 520186 711558
rect 520422 711322 530106 711558
rect 530342 711322 530426 711558
rect 530662 711322 540346 711558
rect 540582 711322 540666 711558
rect 540902 711322 550586 711558
rect 550822 711322 550906 711558
rect 551142 711322 560826 711558
rect 561062 711322 561146 711558
rect 561382 711322 571066 711558
rect 571302 711322 571386 711558
rect 571622 711322 581306 711558
rect 581542 711322 581626 711558
rect 581862 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 18106 711238
rect 18342 711002 18426 711238
rect 18662 711002 28346 711238
rect 28582 711002 28666 711238
rect 28902 711002 38586 711238
rect 38822 711002 38906 711238
rect 39142 711002 48826 711238
rect 49062 711002 49146 711238
rect 49382 711002 59066 711238
rect 59302 711002 59386 711238
rect 59622 711002 69306 711238
rect 69542 711002 69626 711238
rect 69862 711002 79546 711238
rect 79782 711002 79866 711238
rect 80102 711002 89786 711238
rect 90022 711002 90106 711238
rect 90342 711002 100026 711238
rect 100262 711002 100346 711238
rect 100582 711002 110266 711238
rect 110502 711002 110586 711238
rect 110822 711002 120506 711238
rect 120742 711002 120826 711238
rect 121062 711002 130746 711238
rect 130982 711002 131066 711238
rect 131302 711002 140986 711238
rect 141222 711002 141306 711238
rect 141542 711002 151226 711238
rect 151462 711002 151546 711238
rect 151782 711002 161466 711238
rect 161702 711002 161786 711238
rect 162022 711002 171706 711238
rect 171942 711002 172026 711238
rect 172262 711002 181946 711238
rect 182182 711002 182266 711238
rect 182502 711002 192186 711238
rect 192422 711002 192506 711238
rect 192742 711002 202426 711238
rect 202662 711002 202746 711238
rect 202982 711002 212666 711238
rect 212902 711002 212986 711238
rect 213222 711002 222906 711238
rect 223142 711002 223226 711238
rect 223462 711002 233146 711238
rect 233382 711002 233466 711238
rect 233702 711002 243386 711238
rect 243622 711002 243706 711238
rect 243942 711002 253626 711238
rect 253862 711002 253946 711238
rect 254182 711002 263866 711238
rect 264102 711002 264186 711238
rect 264422 711002 274106 711238
rect 274342 711002 274426 711238
rect 274662 711002 284346 711238
rect 284582 711002 284666 711238
rect 284902 711002 294586 711238
rect 294822 711002 294906 711238
rect 295142 711002 304826 711238
rect 305062 711002 305146 711238
rect 305382 711002 315066 711238
rect 315302 711002 315386 711238
rect 315622 711002 325306 711238
rect 325542 711002 325626 711238
rect 325862 711002 335546 711238
rect 335782 711002 335866 711238
rect 336102 711002 345786 711238
rect 346022 711002 346106 711238
rect 346342 711002 356026 711238
rect 356262 711002 356346 711238
rect 356582 711002 366266 711238
rect 366502 711002 366586 711238
rect 366822 711002 376506 711238
rect 376742 711002 376826 711238
rect 377062 711002 386746 711238
rect 386982 711002 387066 711238
rect 387302 711002 396986 711238
rect 397222 711002 397306 711238
rect 397542 711002 407226 711238
rect 407462 711002 407546 711238
rect 407782 711002 417466 711238
rect 417702 711002 417786 711238
rect 418022 711002 427706 711238
rect 427942 711002 428026 711238
rect 428262 711002 437946 711238
rect 438182 711002 438266 711238
rect 438502 711002 448186 711238
rect 448422 711002 448506 711238
rect 448742 711002 458426 711238
rect 458662 711002 458746 711238
rect 458982 711002 468666 711238
rect 468902 711002 468986 711238
rect 469222 711002 478906 711238
rect 479142 711002 479226 711238
rect 479462 711002 489146 711238
rect 489382 711002 489466 711238
rect 489702 711002 499386 711238
rect 499622 711002 499706 711238
rect 499942 711002 509626 711238
rect 509862 711002 509946 711238
rect 510182 711002 519866 711238
rect 520102 711002 520186 711238
rect 520422 711002 530106 711238
rect 530342 711002 530426 711238
rect 530662 711002 540346 711238
rect 540582 711002 540666 711238
rect 540902 711002 550586 711238
rect 550822 711002 550906 711238
rect 551142 711002 560826 711238
rect 561062 711002 561146 711238
rect 561382 711002 571066 711238
rect 571302 711002 571386 711238
rect 571622 711002 581306 711238
rect 581542 711002 581626 711238
rect 581862 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 23226 710598
rect 23462 710362 23546 710598
rect 23782 710362 33466 710598
rect 33702 710362 33786 710598
rect 34022 710362 43706 710598
rect 43942 710362 44026 710598
rect 44262 710362 53946 710598
rect 54182 710362 54266 710598
rect 54502 710362 64186 710598
rect 64422 710362 64506 710598
rect 64742 710362 74426 710598
rect 74662 710362 74746 710598
rect 74982 710362 84666 710598
rect 84902 710362 84986 710598
rect 85222 710362 94906 710598
rect 95142 710362 95226 710598
rect 95462 710362 105146 710598
rect 105382 710362 105466 710598
rect 105702 710362 115386 710598
rect 115622 710362 115706 710598
rect 115942 710362 125626 710598
rect 125862 710362 125946 710598
rect 126182 710362 135866 710598
rect 136102 710362 136186 710598
rect 136422 710362 146106 710598
rect 146342 710362 146426 710598
rect 146662 710362 156346 710598
rect 156582 710362 156666 710598
rect 156902 710362 166586 710598
rect 166822 710362 166906 710598
rect 167142 710362 176826 710598
rect 177062 710362 177146 710598
rect 177382 710362 187066 710598
rect 187302 710362 187386 710598
rect 187622 710362 197306 710598
rect 197542 710362 197626 710598
rect 197862 710362 207546 710598
rect 207782 710362 207866 710598
rect 208102 710362 217786 710598
rect 218022 710362 218106 710598
rect 218342 710362 228026 710598
rect 228262 710362 228346 710598
rect 228582 710362 238266 710598
rect 238502 710362 238586 710598
rect 238822 710362 248506 710598
rect 248742 710362 248826 710598
rect 249062 710362 258746 710598
rect 258982 710362 259066 710598
rect 259302 710362 268986 710598
rect 269222 710362 269306 710598
rect 269542 710362 279226 710598
rect 279462 710362 279546 710598
rect 279782 710362 289466 710598
rect 289702 710362 289786 710598
rect 290022 710362 299706 710598
rect 299942 710362 300026 710598
rect 300262 710362 309946 710598
rect 310182 710362 310266 710598
rect 310502 710362 320186 710598
rect 320422 710362 320506 710598
rect 320742 710362 330426 710598
rect 330662 710362 330746 710598
rect 330982 710362 340666 710598
rect 340902 710362 340986 710598
rect 341222 710362 350906 710598
rect 351142 710362 351226 710598
rect 351462 710362 361146 710598
rect 361382 710362 361466 710598
rect 361702 710362 371386 710598
rect 371622 710362 371706 710598
rect 371942 710362 381626 710598
rect 381862 710362 381946 710598
rect 382182 710362 391866 710598
rect 392102 710362 392186 710598
rect 392422 710362 402106 710598
rect 402342 710362 402426 710598
rect 402662 710362 412346 710598
rect 412582 710362 412666 710598
rect 412902 710362 422586 710598
rect 422822 710362 422906 710598
rect 423142 710362 432826 710598
rect 433062 710362 433146 710598
rect 433382 710362 443066 710598
rect 443302 710362 443386 710598
rect 443622 710362 453306 710598
rect 453542 710362 453626 710598
rect 453862 710362 463546 710598
rect 463782 710362 463866 710598
rect 464102 710362 473786 710598
rect 474022 710362 474106 710598
rect 474342 710362 484026 710598
rect 484262 710362 484346 710598
rect 484582 710362 494266 710598
rect 494502 710362 494586 710598
rect 494822 710362 504506 710598
rect 504742 710362 504826 710598
rect 505062 710362 514746 710598
rect 514982 710362 515066 710598
rect 515302 710362 524986 710598
rect 525222 710362 525306 710598
rect 525542 710362 535226 710598
rect 535462 710362 535546 710598
rect 535782 710362 545466 710598
rect 545702 710362 545786 710598
rect 546022 710362 555706 710598
rect 555942 710362 556026 710598
rect 556262 710362 565946 710598
rect 566182 710362 566266 710598
rect 566502 710362 576186 710598
rect 576422 710362 576506 710598
rect 576742 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 23226 710278
rect 23462 710042 23546 710278
rect 23782 710042 33466 710278
rect 33702 710042 33786 710278
rect 34022 710042 43706 710278
rect 43942 710042 44026 710278
rect 44262 710042 53946 710278
rect 54182 710042 54266 710278
rect 54502 710042 64186 710278
rect 64422 710042 64506 710278
rect 64742 710042 74426 710278
rect 74662 710042 74746 710278
rect 74982 710042 84666 710278
rect 84902 710042 84986 710278
rect 85222 710042 94906 710278
rect 95142 710042 95226 710278
rect 95462 710042 105146 710278
rect 105382 710042 105466 710278
rect 105702 710042 115386 710278
rect 115622 710042 115706 710278
rect 115942 710042 125626 710278
rect 125862 710042 125946 710278
rect 126182 710042 135866 710278
rect 136102 710042 136186 710278
rect 136422 710042 146106 710278
rect 146342 710042 146426 710278
rect 146662 710042 156346 710278
rect 156582 710042 156666 710278
rect 156902 710042 166586 710278
rect 166822 710042 166906 710278
rect 167142 710042 176826 710278
rect 177062 710042 177146 710278
rect 177382 710042 187066 710278
rect 187302 710042 187386 710278
rect 187622 710042 197306 710278
rect 197542 710042 197626 710278
rect 197862 710042 207546 710278
rect 207782 710042 207866 710278
rect 208102 710042 217786 710278
rect 218022 710042 218106 710278
rect 218342 710042 228026 710278
rect 228262 710042 228346 710278
rect 228582 710042 238266 710278
rect 238502 710042 238586 710278
rect 238822 710042 248506 710278
rect 248742 710042 248826 710278
rect 249062 710042 258746 710278
rect 258982 710042 259066 710278
rect 259302 710042 268986 710278
rect 269222 710042 269306 710278
rect 269542 710042 279226 710278
rect 279462 710042 279546 710278
rect 279782 710042 289466 710278
rect 289702 710042 289786 710278
rect 290022 710042 299706 710278
rect 299942 710042 300026 710278
rect 300262 710042 309946 710278
rect 310182 710042 310266 710278
rect 310502 710042 320186 710278
rect 320422 710042 320506 710278
rect 320742 710042 330426 710278
rect 330662 710042 330746 710278
rect 330982 710042 340666 710278
rect 340902 710042 340986 710278
rect 341222 710042 350906 710278
rect 351142 710042 351226 710278
rect 351462 710042 361146 710278
rect 361382 710042 361466 710278
rect 361702 710042 371386 710278
rect 371622 710042 371706 710278
rect 371942 710042 381626 710278
rect 381862 710042 381946 710278
rect 382182 710042 391866 710278
rect 392102 710042 392186 710278
rect 392422 710042 402106 710278
rect 402342 710042 402426 710278
rect 402662 710042 412346 710278
rect 412582 710042 412666 710278
rect 412902 710042 422586 710278
rect 422822 710042 422906 710278
rect 423142 710042 432826 710278
rect 433062 710042 433146 710278
rect 433382 710042 443066 710278
rect 443302 710042 443386 710278
rect 443622 710042 453306 710278
rect 453542 710042 453626 710278
rect 453862 710042 463546 710278
rect 463782 710042 463866 710278
rect 464102 710042 473786 710278
rect 474022 710042 474106 710278
rect 474342 710042 484026 710278
rect 484262 710042 484346 710278
rect 484582 710042 494266 710278
rect 494502 710042 494586 710278
rect 494822 710042 504506 710278
rect 504742 710042 504826 710278
rect 505062 710042 514746 710278
rect 514982 710042 515066 710278
rect 515302 710042 524986 710278
rect 525222 710042 525306 710278
rect 525542 710042 535226 710278
rect 535462 710042 535546 710278
rect 535782 710042 545466 710278
rect 545702 710042 545786 710278
rect 546022 710042 555706 710278
rect 555942 710042 556026 710278
rect 556262 710042 565946 710278
rect 566182 710042 566266 710278
rect 566502 710042 576186 710278
rect 576422 710042 576506 710278
rect 576742 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 14386 709638
rect 14622 709402 14706 709638
rect 14942 709402 24626 709638
rect 24862 709402 24946 709638
rect 25182 709402 34866 709638
rect 35102 709402 35186 709638
rect 35422 709402 45106 709638
rect 45342 709402 45426 709638
rect 45662 709402 55346 709638
rect 55582 709402 55666 709638
rect 55902 709402 65586 709638
rect 65822 709402 65906 709638
rect 66142 709402 75826 709638
rect 76062 709402 76146 709638
rect 76382 709402 86066 709638
rect 86302 709402 86386 709638
rect 86622 709402 96306 709638
rect 96542 709402 96626 709638
rect 96862 709402 106546 709638
rect 106782 709402 106866 709638
rect 107102 709402 116786 709638
rect 117022 709402 117106 709638
rect 117342 709402 127026 709638
rect 127262 709402 127346 709638
rect 127582 709402 137266 709638
rect 137502 709402 137586 709638
rect 137822 709402 147506 709638
rect 147742 709402 147826 709638
rect 148062 709402 157746 709638
rect 157982 709402 158066 709638
rect 158302 709402 167986 709638
rect 168222 709402 168306 709638
rect 168542 709402 178226 709638
rect 178462 709402 178546 709638
rect 178782 709402 188466 709638
rect 188702 709402 188786 709638
rect 189022 709402 198706 709638
rect 198942 709402 199026 709638
rect 199262 709402 208946 709638
rect 209182 709402 209266 709638
rect 209502 709402 219186 709638
rect 219422 709402 219506 709638
rect 219742 709402 229426 709638
rect 229662 709402 229746 709638
rect 229982 709402 239666 709638
rect 239902 709402 239986 709638
rect 240222 709402 249906 709638
rect 250142 709402 250226 709638
rect 250462 709402 260146 709638
rect 260382 709402 260466 709638
rect 260702 709402 270386 709638
rect 270622 709402 270706 709638
rect 270942 709402 280626 709638
rect 280862 709402 280946 709638
rect 281182 709402 290866 709638
rect 291102 709402 291186 709638
rect 291422 709402 301106 709638
rect 301342 709402 301426 709638
rect 301662 709402 311346 709638
rect 311582 709402 311666 709638
rect 311902 709402 321586 709638
rect 321822 709402 321906 709638
rect 322142 709402 331826 709638
rect 332062 709402 332146 709638
rect 332382 709402 342066 709638
rect 342302 709402 342386 709638
rect 342622 709402 352306 709638
rect 352542 709402 352626 709638
rect 352862 709402 362546 709638
rect 362782 709402 362866 709638
rect 363102 709402 372786 709638
rect 373022 709402 373106 709638
rect 373342 709402 383026 709638
rect 383262 709402 383346 709638
rect 383582 709402 393266 709638
rect 393502 709402 393586 709638
rect 393822 709402 403506 709638
rect 403742 709402 403826 709638
rect 404062 709402 413746 709638
rect 413982 709402 414066 709638
rect 414302 709402 423986 709638
rect 424222 709402 424306 709638
rect 424542 709402 434226 709638
rect 434462 709402 434546 709638
rect 434782 709402 444466 709638
rect 444702 709402 444786 709638
rect 445022 709402 454706 709638
rect 454942 709402 455026 709638
rect 455262 709402 464946 709638
rect 465182 709402 465266 709638
rect 465502 709402 475186 709638
rect 475422 709402 475506 709638
rect 475742 709402 485426 709638
rect 485662 709402 485746 709638
rect 485982 709402 495666 709638
rect 495902 709402 495986 709638
rect 496222 709402 505906 709638
rect 506142 709402 506226 709638
rect 506462 709402 516146 709638
rect 516382 709402 516466 709638
rect 516702 709402 526386 709638
rect 526622 709402 526706 709638
rect 526942 709402 536626 709638
rect 536862 709402 536946 709638
rect 537182 709402 546866 709638
rect 547102 709402 547186 709638
rect 547422 709402 557106 709638
rect 557342 709402 557426 709638
rect 557662 709402 567346 709638
rect 567582 709402 567666 709638
rect 567902 709402 577586 709638
rect 577822 709402 577906 709638
rect 578142 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 14386 709318
rect 14622 709082 14706 709318
rect 14942 709082 24626 709318
rect 24862 709082 24946 709318
rect 25182 709082 34866 709318
rect 35102 709082 35186 709318
rect 35422 709082 45106 709318
rect 45342 709082 45426 709318
rect 45662 709082 55346 709318
rect 55582 709082 55666 709318
rect 55902 709082 65586 709318
rect 65822 709082 65906 709318
rect 66142 709082 75826 709318
rect 76062 709082 76146 709318
rect 76382 709082 86066 709318
rect 86302 709082 86386 709318
rect 86622 709082 96306 709318
rect 96542 709082 96626 709318
rect 96862 709082 106546 709318
rect 106782 709082 106866 709318
rect 107102 709082 116786 709318
rect 117022 709082 117106 709318
rect 117342 709082 127026 709318
rect 127262 709082 127346 709318
rect 127582 709082 137266 709318
rect 137502 709082 137586 709318
rect 137822 709082 147506 709318
rect 147742 709082 147826 709318
rect 148062 709082 157746 709318
rect 157982 709082 158066 709318
rect 158302 709082 167986 709318
rect 168222 709082 168306 709318
rect 168542 709082 178226 709318
rect 178462 709082 178546 709318
rect 178782 709082 188466 709318
rect 188702 709082 188786 709318
rect 189022 709082 198706 709318
rect 198942 709082 199026 709318
rect 199262 709082 208946 709318
rect 209182 709082 209266 709318
rect 209502 709082 219186 709318
rect 219422 709082 219506 709318
rect 219742 709082 229426 709318
rect 229662 709082 229746 709318
rect 229982 709082 239666 709318
rect 239902 709082 239986 709318
rect 240222 709082 249906 709318
rect 250142 709082 250226 709318
rect 250462 709082 260146 709318
rect 260382 709082 260466 709318
rect 260702 709082 270386 709318
rect 270622 709082 270706 709318
rect 270942 709082 280626 709318
rect 280862 709082 280946 709318
rect 281182 709082 290866 709318
rect 291102 709082 291186 709318
rect 291422 709082 301106 709318
rect 301342 709082 301426 709318
rect 301662 709082 311346 709318
rect 311582 709082 311666 709318
rect 311902 709082 321586 709318
rect 321822 709082 321906 709318
rect 322142 709082 331826 709318
rect 332062 709082 332146 709318
rect 332382 709082 342066 709318
rect 342302 709082 342386 709318
rect 342622 709082 352306 709318
rect 352542 709082 352626 709318
rect 352862 709082 362546 709318
rect 362782 709082 362866 709318
rect 363102 709082 372786 709318
rect 373022 709082 373106 709318
rect 373342 709082 383026 709318
rect 383262 709082 383346 709318
rect 383582 709082 393266 709318
rect 393502 709082 393586 709318
rect 393822 709082 403506 709318
rect 403742 709082 403826 709318
rect 404062 709082 413746 709318
rect 413982 709082 414066 709318
rect 414302 709082 423986 709318
rect 424222 709082 424306 709318
rect 424542 709082 434226 709318
rect 434462 709082 434546 709318
rect 434782 709082 444466 709318
rect 444702 709082 444786 709318
rect 445022 709082 454706 709318
rect 454942 709082 455026 709318
rect 455262 709082 464946 709318
rect 465182 709082 465266 709318
rect 465502 709082 475186 709318
rect 475422 709082 475506 709318
rect 475742 709082 485426 709318
rect 485662 709082 485746 709318
rect 485982 709082 495666 709318
rect 495902 709082 495986 709318
rect 496222 709082 505906 709318
rect 506142 709082 506226 709318
rect 506462 709082 516146 709318
rect 516382 709082 516466 709318
rect 516702 709082 526386 709318
rect 526622 709082 526706 709318
rect 526942 709082 536626 709318
rect 536862 709082 536946 709318
rect 537182 709082 546866 709318
rect 547102 709082 547186 709318
rect 547422 709082 557106 709318
rect 557342 709082 557426 709318
rect 557662 709082 567346 709318
rect 567582 709082 567666 709318
rect 567902 709082 577586 709318
rect 577822 709082 577906 709318
rect 578142 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 19506 708678
rect 19742 708442 19826 708678
rect 20062 708442 29746 708678
rect 29982 708442 30066 708678
rect 30302 708442 39986 708678
rect 40222 708442 40306 708678
rect 40542 708442 50226 708678
rect 50462 708442 50546 708678
rect 50782 708442 60466 708678
rect 60702 708442 60786 708678
rect 61022 708442 70706 708678
rect 70942 708442 71026 708678
rect 71262 708442 80946 708678
rect 81182 708442 81266 708678
rect 81502 708442 91186 708678
rect 91422 708442 91506 708678
rect 91742 708442 101426 708678
rect 101662 708442 101746 708678
rect 101982 708442 111666 708678
rect 111902 708442 111986 708678
rect 112222 708442 121906 708678
rect 122142 708442 122226 708678
rect 122462 708442 132146 708678
rect 132382 708442 132466 708678
rect 132702 708442 142386 708678
rect 142622 708442 142706 708678
rect 142942 708442 152626 708678
rect 152862 708442 152946 708678
rect 153182 708442 162866 708678
rect 163102 708442 163186 708678
rect 163422 708442 173106 708678
rect 173342 708442 173426 708678
rect 173662 708442 183346 708678
rect 183582 708442 183666 708678
rect 183902 708442 193586 708678
rect 193822 708442 193906 708678
rect 194142 708442 203826 708678
rect 204062 708442 204146 708678
rect 204382 708442 214066 708678
rect 214302 708442 214386 708678
rect 214622 708442 224306 708678
rect 224542 708442 224626 708678
rect 224862 708442 234546 708678
rect 234782 708442 234866 708678
rect 235102 708442 244786 708678
rect 245022 708442 245106 708678
rect 245342 708442 255026 708678
rect 255262 708442 255346 708678
rect 255582 708442 265266 708678
rect 265502 708442 265586 708678
rect 265822 708442 275506 708678
rect 275742 708442 275826 708678
rect 276062 708442 285746 708678
rect 285982 708442 286066 708678
rect 286302 708442 295986 708678
rect 296222 708442 296306 708678
rect 296542 708442 306226 708678
rect 306462 708442 306546 708678
rect 306782 708442 316466 708678
rect 316702 708442 316786 708678
rect 317022 708442 326706 708678
rect 326942 708442 327026 708678
rect 327262 708442 336946 708678
rect 337182 708442 337266 708678
rect 337502 708442 347186 708678
rect 347422 708442 347506 708678
rect 347742 708442 357426 708678
rect 357662 708442 357746 708678
rect 357982 708442 367666 708678
rect 367902 708442 367986 708678
rect 368222 708442 377906 708678
rect 378142 708442 378226 708678
rect 378462 708442 388146 708678
rect 388382 708442 388466 708678
rect 388702 708442 398386 708678
rect 398622 708442 398706 708678
rect 398942 708442 408626 708678
rect 408862 708442 408946 708678
rect 409182 708442 418866 708678
rect 419102 708442 419186 708678
rect 419422 708442 429106 708678
rect 429342 708442 429426 708678
rect 429662 708442 439346 708678
rect 439582 708442 439666 708678
rect 439902 708442 449586 708678
rect 449822 708442 449906 708678
rect 450142 708442 459826 708678
rect 460062 708442 460146 708678
rect 460382 708442 470066 708678
rect 470302 708442 470386 708678
rect 470622 708442 480306 708678
rect 480542 708442 480626 708678
rect 480862 708442 490546 708678
rect 490782 708442 490866 708678
rect 491102 708442 500786 708678
rect 501022 708442 501106 708678
rect 501342 708442 511026 708678
rect 511262 708442 511346 708678
rect 511582 708442 521266 708678
rect 521502 708442 521586 708678
rect 521822 708442 531506 708678
rect 531742 708442 531826 708678
rect 532062 708442 541746 708678
rect 541982 708442 542066 708678
rect 542302 708442 551986 708678
rect 552222 708442 552306 708678
rect 552542 708442 562226 708678
rect 562462 708442 562546 708678
rect 562782 708442 572466 708678
rect 572702 708442 572786 708678
rect 573022 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 19506 708358
rect 19742 708122 19826 708358
rect 20062 708122 29746 708358
rect 29982 708122 30066 708358
rect 30302 708122 39986 708358
rect 40222 708122 40306 708358
rect 40542 708122 50226 708358
rect 50462 708122 50546 708358
rect 50782 708122 60466 708358
rect 60702 708122 60786 708358
rect 61022 708122 70706 708358
rect 70942 708122 71026 708358
rect 71262 708122 80946 708358
rect 81182 708122 81266 708358
rect 81502 708122 91186 708358
rect 91422 708122 91506 708358
rect 91742 708122 101426 708358
rect 101662 708122 101746 708358
rect 101982 708122 111666 708358
rect 111902 708122 111986 708358
rect 112222 708122 121906 708358
rect 122142 708122 122226 708358
rect 122462 708122 132146 708358
rect 132382 708122 132466 708358
rect 132702 708122 142386 708358
rect 142622 708122 142706 708358
rect 142942 708122 152626 708358
rect 152862 708122 152946 708358
rect 153182 708122 162866 708358
rect 163102 708122 163186 708358
rect 163422 708122 173106 708358
rect 173342 708122 173426 708358
rect 173662 708122 183346 708358
rect 183582 708122 183666 708358
rect 183902 708122 193586 708358
rect 193822 708122 193906 708358
rect 194142 708122 203826 708358
rect 204062 708122 204146 708358
rect 204382 708122 214066 708358
rect 214302 708122 214386 708358
rect 214622 708122 224306 708358
rect 224542 708122 224626 708358
rect 224862 708122 234546 708358
rect 234782 708122 234866 708358
rect 235102 708122 244786 708358
rect 245022 708122 245106 708358
rect 245342 708122 255026 708358
rect 255262 708122 255346 708358
rect 255582 708122 265266 708358
rect 265502 708122 265586 708358
rect 265822 708122 275506 708358
rect 275742 708122 275826 708358
rect 276062 708122 285746 708358
rect 285982 708122 286066 708358
rect 286302 708122 295986 708358
rect 296222 708122 296306 708358
rect 296542 708122 306226 708358
rect 306462 708122 306546 708358
rect 306782 708122 316466 708358
rect 316702 708122 316786 708358
rect 317022 708122 326706 708358
rect 326942 708122 327026 708358
rect 327262 708122 336946 708358
rect 337182 708122 337266 708358
rect 337502 708122 347186 708358
rect 347422 708122 347506 708358
rect 347742 708122 357426 708358
rect 357662 708122 357746 708358
rect 357982 708122 367666 708358
rect 367902 708122 367986 708358
rect 368222 708122 377906 708358
rect 378142 708122 378226 708358
rect 378462 708122 388146 708358
rect 388382 708122 388466 708358
rect 388702 708122 398386 708358
rect 398622 708122 398706 708358
rect 398942 708122 408626 708358
rect 408862 708122 408946 708358
rect 409182 708122 418866 708358
rect 419102 708122 419186 708358
rect 419422 708122 429106 708358
rect 429342 708122 429426 708358
rect 429662 708122 439346 708358
rect 439582 708122 439666 708358
rect 439902 708122 449586 708358
rect 449822 708122 449906 708358
rect 450142 708122 459826 708358
rect 460062 708122 460146 708358
rect 460382 708122 470066 708358
rect 470302 708122 470386 708358
rect 470622 708122 480306 708358
rect 480542 708122 480626 708358
rect 480862 708122 490546 708358
rect 490782 708122 490866 708358
rect 491102 708122 500786 708358
rect 501022 708122 501106 708358
rect 501342 708122 511026 708358
rect 511262 708122 511346 708358
rect 511582 708122 521266 708358
rect 521502 708122 521586 708358
rect 521822 708122 531506 708358
rect 531742 708122 531826 708358
rect 532062 708122 541746 708358
rect 541982 708122 542066 708358
rect 542302 708122 551986 708358
rect 552222 708122 552306 708358
rect 552542 708122 562226 708358
rect 562462 708122 562546 708358
rect 562782 708122 572466 708358
rect 572702 708122 572786 708358
rect 573022 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 10666 707718
rect 10902 707482 10986 707718
rect 11222 707482 20906 707718
rect 21142 707482 21226 707718
rect 21462 707482 31146 707718
rect 31382 707482 31466 707718
rect 31702 707482 41386 707718
rect 41622 707482 41706 707718
rect 41942 707482 51626 707718
rect 51862 707482 51946 707718
rect 52182 707482 61866 707718
rect 62102 707482 62186 707718
rect 62422 707482 72106 707718
rect 72342 707482 72426 707718
rect 72662 707482 82346 707718
rect 82582 707482 82666 707718
rect 82902 707482 92586 707718
rect 92822 707482 92906 707718
rect 93142 707482 102826 707718
rect 103062 707482 103146 707718
rect 103382 707482 113066 707718
rect 113302 707482 113386 707718
rect 113622 707482 123306 707718
rect 123542 707482 123626 707718
rect 123862 707482 133546 707718
rect 133782 707482 133866 707718
rect 134102 707482 143786 707718
rect 144022 707482 144106 707718
rect 144342 707482 154026 707718
rect 154262 707482 154346 707718
rect 154582 707482 164266 707718
rect 164502 707482 164586 707718
rect 164822 707482 174506 707718
rect 174742 707482 174826 707718
rect 175062 707482 184746 707718
rect 184982 707482 185066 707718
rect 185302 707482 194986 707718
rect 195222 707482 195306 707718
rect 195542 707482 205226 707718
rect 205462 707482 205546 707718
rect 205782 707482 215466 707718
rect 215702 707482 215786 707718
rect 216022 707482 225706 707718
rect 225942 707482 226026 707718
rect 226262 707482 235946 707718
rect 236182 707482 236266 707718
rect 236502 707482 246186 707718
rect 246422 707482 246506 707718
rect 246742 707482 256426 707718
rect 256662 707482 256746 707718
rect 256982 707482 266666 707718
rect 266902 707482 266986 707718
rect 267222 707482 276906 707718
rect 277142 707482 277226 707718
rect 277462 707482 287146 707718
rect 287382 707482 287466 707718
rect 287702 707482 297386 707718
rect 297622 707482 297706 707718
rect 297942 707482 307626 707718
rect 307862 707482 307946 707718
rect 308182 707482 317866 707718
rect 318102 707482 318186 707718
rect 318422 707482 328106 707718
rect 328342 707482 328426 707718
rect 328662 707482 338346 707718
rect 338582 707482 338666 707718
rect 338902 707482 348586 707718
rect 348822 707482 348906 707718
rect 349142 707482 358826 707718
rect 359062 707482 359146 707718
rect 359382 707482 369066 707718
rect 369302 707482 369386 707718
rect 369622 707482 379306 707718
rect 379542 707482 379626 707718
rect 379862 707482 389546 707718
rect 389782 707482 389866 707718
rect 390102 707482 399786 707718
rect 400022 707482 400106 707718
rect 400342 707482 410026 707718
rect 410262 707482 410346 707718
rect 410582 707482 420266 707718
rect 420502 707482 420586 707718
rect 420822 707482 430506 707718
rect 430742 707482 430826 707718
rect 431062 707482 440746 707718
rect 440982 707482 441066 707718
rect 441302 707482 450986 707718
rect 451222 707482 451306 707718
rect 451542 707482 461226 707718
rect 461462 707482 461546 707718
rect 461782 707482 471466 707718
rect 471702 707482 471786 707718
rect 472022 707482 481706 707718
rect 481942 707482 482026 707718
rect 482262 707482 491946 707718
rect 492182 707482 492266 707718
rect 492502 707482 502186 707718
rect 502422 707482 502506 707718
rect 502742 707482 512426 707718
rect 512662 707482 512746 707718
rect 512982 707482 522666 707718
rect 522902 707482 522986 707718
rect 523222 707482 532906 707718
rect 533142 707482 533226 707718
rect 533462 707482 543146 707718
rect 543382 707482 543466 707718
rect 543702 707482 553386 707718
rect 553622 707482 553706 707718
rect 553942 707482 563626 707718
rect 563862 707482 563946 707718
rect 564182 707482 573866 707718
rect 574102 707482 574186 707718
rect 574422 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 10666 707398
rect 10902 707162 10986 707398
rect 11222 707162 20906 707398
rect 21142 707162 21226 707398
rect 21462 707162 31146 707398
rect 31382 707162 31466 707398
rect 31702 707162 41386 707398
rect 41622 707162 41706 707398
rect 41942 707162 51626 707398
rect 51862 707162 51946 707398
rect 52182 707162 61866 707398
rect 62102 707162 62186 707398
rect 62422 707162 72106 707398
rect 72342 707162 72426 707398
rect 72662 707162 82346 707398
rect 82582 707162 82666 707398
rect 82902 707162 92586 707398
rect 92822 707162 92906 707398
rect 93142 707162 102826 707398
rect 103062 707162 103146 707398
rect 103382 707162 113066 707398
rect 113302 707162 113386 707398
rect 113622 707162 123306 707398
rect 123542 707162 123626 707398
rect 123862 707162 133546 707398
rect 133782 707162 133866 707398
rect 134102 707162 143786 707398
rect 144022 707162 144106 707398
rect 144342 707162 154026 707398
rect 154262 707162 154346 707398
rect 154582 707162 164266 707398
rect 164502 707162 164586 707398
rect 164822 707162 174506 707398
rect 174742 707162 174826 707398
rect 175062 707162 184746 707398
rect 184982 707162 185066 707398
rect 185302 707162 194986 707398
rect 195222 707162 195306 707398
rect 195542 707162 205226 707398
rect 205462 707162 205546 707398
rect 205782 707162 215466 707398
rect 215702 707162 215786 707398
rect 216022 707162 225706 707398
rect 225942 707162 226026 707398
rect 226262 707162 235946 707398
rect 236182 707162 236266 707398
rect 236502 707162 246186 707398
rect 246422 707162 246506 707398
rect 246742 707162 256426 707398
rect 256662 707162 256746 707398
rect 256982 707162 266666 707398
rect 266902 707162 266986 707398
rect 267222 707162 276906 707398
rect 277142 707162 277226 707398
rect 277462 707162 287146 707398
rect 287382 707162 287466 707398
rect 287702 707162 297386 707398
rect 297622 707162 297706 707398
rect 297942 707162 307626 707398
rect 307862 707162 307946 707398
rect 308182 707162 317866 707398
rect 318102 707162 318186 707398
rect 318422 707162 328106 707398
rect 328342 707162 328426 707398
rect 328662 707162 338346 707398
rect 338582 707162 338666 707398
rect 338902 707162 348586 707398
rect 348822 707162 348906 707398
rect 349142 707162 358826 707398
rect 359062 707162 359146 707398
rect 359382 707162 369066 707398
rect 369302 707162 369386 707398
rect 369622 707162 379306 707398
rect 379542 707162 379626 707398
rect 379862 707162 389546 707398
rect 389782 707162 389866 707398
rect 390102 707162 399786 707398
rect 400022 707162 400106 707398
rect 400342 707162 410026 707398
rect 410262 707162 410346 707398
rect 410582 707162 420266 707398
rect 420502 707162 420586 707398
rect 420822 707162 430506 707398
rect 430742 707162 430826 707398
rect 431062 707162 440746 707398
rect 440982 707162 441066 707398
rect 441302 707162 450986 707398
rect 451222 707162 451306 707398
rect 451542 707162 461226 707398
rect 461462 707162 461546 707398
rect 461782 707162 471466 707398
rect 471702 707162 471786 707398
rect 472022 707162 481706 707398
rect 481942 707162 482026 707398
rect 482262 707162 491946 707398
rect 492182 707162 492266 707398
rect 492502 707162 502186 707398
rect 502422 707162 502506 707398
rect 502742 707162 512426 707398
rect 512662 707162 512746 707398
rect 512982 707162 522666 707398
rect 522902 707162 522986 707398
rect 523222 707162 532906 707398
rect 533142 707162 533226 707398
rect 533462 707162 543146 707398
rect 543382 707162 543466 707398
rect 543702 707162 553386 707398
rect 553622 707162 553706 707398
rect 553942 707162 563626 707398
rect 563862 707162 563946 707398
rect 564182 707162 573866 707398
rect 574102 707162 574186 707398
rect 574422 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 15786 706758
rect 16022 706522 16106 706758
rect 16342 706522 26026 706758
rect 26262 706522 26346 706758
rect 26582 706522 36266 706758
rect 36502 706522 36586 706758
rect 36822 706522 46506 706758
rect 46742 706522 46826 706758
rect 47062 706522 56746 706758
rect 56982 706522 57066 706758
rect 57302 706522 66986 706758
rect 67222 706522 67306 706758
rect 67542 706522 77226 706758
rect 77462 706522 77546 706758
rect 77782 706522 87466 706758
rect 87702 706522 87786 706758
rect 88022 706522 97706 706758
rect 97942 706522 98026 706758
rect 98262 706522 107946 706758
rect 108182 706522 108266 706758
rect 108502 706522 118186 706758
rect 118422 706522 118506 706758
rect 118742 706522 128426 706758
rect 128662 706522 128746 706758
rect 128982 706522 138666 706758
rect 138902 706522 138986 706758
rect 139222 706522 148906 706758
rect 149142 706522 149226 706758
rect 149462 706522 159146 706758
rect 159382 706522 159466 706758
rect 159702 706522 169386 706758
rect 169622 706522 169706 706758
rect 169942 706522 179626 706758
rect 179862 706522 179946 706758
rect 180182 706522 189866 706758
rect 190102 706522 190186 706758
rect 190422 706522 200106 706758
rect 200342 706522 200426 706758
rect 200662 706522 210346 706758
rect 210582 706522 210666 706758
rect 210902 706522 220586 706758
rect 220822 706522 220906 706758
rect 221142 706522 230826 706758
rect 231062 706522 231146 706758
rect 231382 706522 241066 706758
rect 241302 706522 241386 706758
rect 241622 706522 251306 706758
rect 251542 706522 251626 706758
rect 251862 706522 261546 706758
rect 261782 706522 261866 706758
rect 262102 706522 271786 706758
rect 272022 706522 272106 706758
rect 272342 706522 282026 706758
rect 282262 706522 282346 706758
rect 282582 706522 292266 706758
rect 292502 706522 292586 706758
rect 292822 706522 302506 706758
rect 302742 706522 302826 706758
rect 303062 706522 312746 706758
rect 312982 706522 313066 706758
rect 313302 706522 322986 706758
rect 323222 706522 323306 706758
rect 323542 706522 333226 706758
rect 333462 706522 333546 706758
rect 333782 706522 343466 706758
rect 343702 706522 343786 706758
rect 344022 706522 353706 706758
rect 353942 706522 354026 706758
rect 354262 706522 363946 706758
rect 364182 706522 364266 706758
rect 364502 706522 374186 706758
rect 374422 706522 374506 706758
rect 374742 706522 384426 706758
rect 384662 706522 384746 706758
rect 384982 706522 394666 706758
rect 394902 706522 394986 706758
rect 395222 706522 404906 706758
rect 405142 706522 405226 706758
rect 405462 706522 415146 706758
rect 415382 706522 415466 706758
rect 415702 706522 425386 706758
rect 425622 706522 425706 706758
rect 425942 706522 435626 706758
rect 435862 706522 435946 706758
rect 436182 706522 445866 706758
rect 446102 706522 446186 706758
rect 446422 706522 456106 706758
rect 456342 706522 456426 706758
rect 456662 706522 466346 706758
rect 466582 706522 466666 706758
rect 466902 706522 476586 706758
rect 476822 706522 476906 706758
rect 477142 706522 486826 706758
rect 487062 706522 487146 706758
rect 487382 706522 497066 706758
rect 497302 706522 497386 706758
rect 497622 706522 507306 706758
rect 507542 706522 507626 706758
rect 507862 706522 517546 706758
rect 517782 706522 517866 706758
rect 518102 706522 527786 706758
rect 528022 706522 528106 706758
rect 528342 706522 538026 706758
rect 538262 706522 538346 706758
rect 538582 706522 548266 706758
rect 548502 706522 548586 706758
rect 548822 706522 558506 706758
rect 558742 706522 558826 706758
rect 559062 706522 568746 706758
rect 568982 706522 569066 706758
rect 569302 706522 578986 706758
rect 579222 706522 579306 706758
rect 579542 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 15786 706438
rect 16022 706202 16106 706438
rect 16342 706202 26026 706438
rect 26262 706202 26346 706438
rect 26582 706202 36266 706438
rect 36502 706202 36586 706438
rect 36822 706202 46506 706438
rect 46742 706202 46826 706438
rect 47062 706202 56746 706438
rect 56982 706202 57066 706438
rect 57302 706202 66986 706438
rect 67222 706202 67306 706438
rect 67542 706202 77226 706438
rect 77462 706202 77546 706438
rect 77782 706202 87466 706438
rect 87702 706202 87786 706438
rect 88022 706202 97706 706438
rect 97942 706202 98026 706438
rect 98262 706202 107946 706438
rect 108182 706202 108266 706438
rect 108502 706202 118186 706438
rect 118422 706202 118506 706438
rect 118742 706202 128426 706438
rect 128662 706202 128746 706438
rect 128982 706202 138666 706438
rect 138902 706202 138986 706438
rect 139222 706202 148906 706438
rect 149142 706202 149226 706438
rect 149462 706202 159146 706438
rect 159382 706202 159466 706438
rect 159702 706202 169386 706438
rect 169622 706202 169706 706438
rect 169942 706202 179626 706438
rect 179862 706202 179946 706438
rect 180182 706202 189866 706438
rect 190102 706202 190186 706438
rect 190422 706202 200106 706438
rect 200342 706202 200426 706438
rect 200662 706202 210346 706438
rect 210582 706202 210666 706438
rect 210902 706202 220586 706438
rect 220822 706202 220906 706438
rect 221142 706202 230826 706438
rect 231062 706202 231146 706438
rect 231382 706202 241066 706438
rect 241302 706202 241386 706438
rect 241622 706202 251306 706438
rect 251542 706202 251626 706438
rect 251862 706202 261546 706438
rect 261782 706202 261866 706438
rect 262102 706202 271786 706438
rect 272022 706202 272106 706438
rect 272342 706202 282026 706438
rect 282262 706202 282346 706438
rect 282582 706202 292266 706438
rect 292502 706202 292586 706438
rect 292822 706202 302506 706438
rect 302742 706202 302826 706438
rect 303062 706202 312746 706438
rect 312982 706202 313066 706438
rect 313302 706202 322986 706438
rect 323222 706202 323306 706438
rect 323542 706202 333226 706438
rect 333462 706202 333546 706438
rect 333782 706202 343466 706438
rect 343702 706202 343786 706438
rect 344022 706202 353706 706438
rect 353942 706202 354026 706438
rect 354262 706202 363946 706438
rect 364182 706202 364266 706438
rect 364502 706202 374186 706438
rect 374422 706202 374506 706438
rect 374742 706202 384426 706438
rect 384662 706202 384746 706438
rect 384982 706202 394666 706438
rect 394902 706202 394986 706438
rect 395222 706202 404906 706438
rect 405142 706202 405226 706438
rect 405462 706202 415146 706438
rect 415382 706202 415466 706438
rect 415702 706202 425386 706438
rect 425622 706202 425706 706438
rect 425942 706202 435626 706438
rect 435862 706202 435946 706438
rect 436182 706202 445866 706438
rect 446102 706202 446186 706438
rect 446422 706202 456106 706438
rect 456342 706202 456426 706438
rect 456662 706202 466346 706438
rect 466582 706202 466666 706438
rect 466902 706202 476586 706438
rect 476822 706202 476906 706438
rect 477142 706202 486826 706438
rect 487062 706202 487146 706438
rect 487382 706202 497066 706438
rect 497302 706202 497386 706438
rect 497622 706202 507306 706438
rect 507542 706202 507626 706438
rect 507862 706202 517546 706438
rect 517782 706202 517866 706438
rect 518102 706202 527786 706438
rect 528022 706202 528106 706438
rect 528342 706202 538026 706438
rect 538262 706202 538346 706438
rect 538582 706202 548266 706438
rect 548502 706202 548586 706438
rect 548822 706202 558506 706438
rect 558742 706202 558826 706438
rect 559062 706202 568746 706438
rect 568982 706202 569066 706438
rect 569302 706202 578986 706438
rect 579222 706202 579306 706438
rect 579542 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6946 705798
rect 7182 705562 7266 705798
rect 7502 705562 17186 705798
rect 17422 705562 17506 705798
rect 17742 705562 27426 705798
rect 27662 705562 27746 705798
rect 27982 705562 37666 705798
rect 37902 705562 37986 705798
rect 38222 705562 47906 705798
rect 48142 705562 48226 705798
rect 48462 705562 58146 705798
rect 58382 705562 58466 705798
rect 58702 705562 68386 705798
rect 68622 705562 68706 705798
rect 68942 705562 78626 705798
rect 78862 705562 78946 705798
rect 79182 705562 88866 705798
rect 89102 705562 89186 705798
rect 89422 705562 99106 705798
rect 99342 705562 99426 705798
rect 99662 705562 109346 705798
rect 109582 705562 109666 705798
rect 109902 705562 119586 705798
rect 119822 705562 119906 705798
rect 120142 705562 129826 705798
rect 130062 705562 130146 705798
rect 130382 705562 140066 705798
rect 140302 705562 140386 705798
rect 140622 705562 150306 705798
rect 150542 705562 150626 705798
rect 150862 705562 160546 705798
rect 160782 705562 160866 705798
rect 161102 705562 170786 705798
rect 171022 705562 171106 705798
rect 171342 705562 181026 705798
rect 181262 705562 181346 705798
rect 181582 705562 191266 705798
rect 191502 705562 191586 705798
rect 191822 705562 201506 705798
rect 201742 705562 201826 705798
rect 202062 705562 211746 705798
rect 211982 705562 212066 705798
rect 212302 705562 221986 705798
rect 222222 705562 222306 705798
rect 222542 705562 232226 705798
rect 232462 705562 232546 705798
rect 232782 705562 242466 705798
rect 242702 705562 242786 705798
rect 243022 705562 252706 705798
rect 252942 705562 253026 705798
rect 253262 705562 262946 705798
rect 263182 705562 263266 705798
rect 263502 705562 273186 705798
rect 273422 705562 273506 705798
rect 273742 705562 283426 705798
rect 283662 705562 283746 705798
rect 283982 705562 293666 705798
rect 293902 705562 293986 705798
rect 294222 705562 303906 705798
rect 304142 705562 304226 705798
rect 304462 705562 314146 705798
rect 314382 705562 314466 705798
rect 314702 705562 324386 705798
rect 324622 705562 324706 705798
rect 324942 705562 334626 705798
rect 334862 705562 334946 705798
rect 335182 705562 344866 705798
rect 345102 705562 345186 705798
rect 345422 705562 355106 705798
rect 355342 705562 355426 705798
rect 355662 705562 365346 705798
rect 365582 705562 365666 705798
rect 365902 705562 375586 705798
rect 375822 705562 375906 705798
rect 376142 705562 385826 705798
rect 386062 705562 386146 705798
rect 386382 705562 396066 705798
rect 396302 705562 396386 705798
rect 396622 705562 406306 705798
rect 406542 705562 406626 705798
rect 406862 705562 416546 705798
rect 416782 705562 416866 705798
rect 417102 705562 426786 705798
rect 427022 705562 427106 705798
rect 427342 705562 437026 705798
rect 437262 705562 437346 705798
rect 437582 705562 447266 705798
rect 447502 705562 447586 705798
rect 447822 705562 457506 705798
rect 457742 705562 457826 705798
rect 458062 705562 467746 705798
rect 467982 705562 468066 705798
rect 468302 705562 477986 705798
rect 478222 705562 478306 705798
rect 478542 705562 488226 705798
rect 488462 705562 488546 705798
rect 488782 705562 498466 705798
rect 498702 705562 498786 705798
rect 499022 705562 508706 705798
rect 508942 705562 509026 705798
rect 509262 705562 518946 705798
rect 519182 705562 519266 705798
rect 519502 705562 529186 705798
rect 529422 705562 529506 705798
rect 529742 705562 539426 705798
rect 539662 705562 539746 705798
rect 539982 705562 549666 705798
rect 549902 705562 549986 705798
rect 550222 705562 559906 705798
rect 560142 705562 560226 705798
rect 560462 705562 570146 705798
rect 570382 705562 570466 705798
rect 570702 705562 580386 705798
rect 580622 705562 580706 705798
rect 580942 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6946 705478
rect 7182 705242 7266 705478
rect 7502 705242 17186 705478
rect 17422 705242 17506 705478
rect 17742 705242 27426 705478
rect 27662 705242 27746 705478
rect 27982 705242 37666 705478
rect 37902 705242 37986 705478
rect 38222 705242 47906 705478
rect 48142 705242 48226 705478
rect 48462 705242 58146 705478
rect 58382 705242 58466 705478
rect 58702 705242 68386 705478
rect 68622 705242 68706 705478
rect 68942 705242 78626 705478
rect 78862 705242 78946 705478
rect 79182 705242 88866 705478
rect 89102 705242 89186 705478
rect 89422 705242 99106 705478
rect 99342 705242 99426 705478
rect 99662 705242 109346 705478
rect 109582 705242 109666 705478
rect 109902 705242 119586 705478
rect 119822 705242 119906 705478
rect 120142 705242 129826 705478
rect 130062 705242 130146 705478
rect 130382 705242 140066 705478
rect 140302 705242 140386 705478
rect 140622 705242 150306 705478
rect 150542 705242 150626 705478
rect 150862 705242 160546 705478
rect 160782 705242 160866 705478
rect 161102 705242 170786 705478
rect 171022 705242 171106 705478
rect 171342 705242 181026 705478
rect 181262 705242 181346 705478
rect 181582 705242 191266 705478
rect 191502 705242 191586 705478
rect 191822 705242 201506 705478
rect 201742 705242 201826 705478
rect 202062 705242 211746 705478
rect 211982 705242 212066 705478
rect 212302 705242 221986 705478
rect 222222 705242 222306 705478
rect 222542 705242 232226 705478
rect 232462 705242 232546 705478
rect 232782 705242 242466 705478
rect 242702 705242 242786 705478
rect 243022 705242 252706 705478
rect 252942 705242 253026 705478
rect 253262 705242 262946 705478
rect 263182 705242 263266 705478
rect 263502 705242 273186 705478
rect 273422 705242 273506 705478
rect 273742 705242 283426 705478
rect 283662 705242 283746 705478
rect 283982 705242 293666 705478
rect 293902 705242 293986 705478
rect 294222 705242 303906 705478
rect 304142 705242 304226 705478
rect 304462 705242 314146 705478
rect 314382 705242 314466 705478
rect 314702 705242 324386 705478
rect 324622 705242 324706 705478
rect 324942 705242 334626 705478
rect 334862 705242 334946 705478
rect 335182 705242 344866 705478
rect 345102 705242 345186 705478
rect 345422 705242 355106 705478
rect 355342 705242 355426 705478
rect 355662 705242 365346 705478
rect 365582 705242 365666 705478
rect 365902 705242 375586 705478
rect 375822 705242 375906 705478
rect 376142 705242 385826 705478
rect 386062 705242 386146 705478
rect 386382 705242 396066 705478
rect 396302 705242 396386 705478
rect 396622 705242 406306 705478
rect 406542 705242 406626 705478
rect 406862 705242 416546 705478
rect 416782 705242 416866 705478
rect 417102 705242 426786 705478
rect 427022 705242 427106 705478
rect 427342 705242 437026 705478
rect 437262 705242 437346 705478
rect 437582 705242 447266 705478
rect 447502 705242 447586 705478
rect 447822 705242 457506 705478
rect 457742 705242 457826 705478
rect 458062 705242 467746 705478
rect 467982 705242 468066 705478
rect 468302 705242 477986 705478
rect 478222 705242 478306 705478
rect 478542 705242 488226 705478
rect 488462 705242 488546 705478
rect 488782 705242 498466 705478
rect 498702 705242 498786 705478
rect 499022 705242 508706 705478
rect 508942 705242 509026 705478
rect 509262 705242 518946 705478
rect 519182 705242 519266 705478
rect 519502 705242 529186 705478
rect 529422 705242 529506 705478
rect 529742 705242 539426 705478
rect 539662 705242 539746 705478
rect 539982 705242 549666 705478
rect 549902 705242 549986 705478
rect 550222 705242 559906 705478
rect 560142 705242 560226 705478
rect 560462 705242 570146 705478
rect 570382 705242 570466 705478
rect 570702 705242 580386 705478
rect 580622 705242 580706 705478
rect 580942 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 12066 704838
rect 12302 704602 12386 704838
rect 12622 704602 22306 704838
rect 22542 704602 22626 704838
rect 22862 704602 32546 704838
rect 32782 704602 32866 704838
rect 33102 704602 42786 704838
rect 43022 704602 43106 704838
rect 43342 704602 53026 704838
rect 53262 704602 53346 704838
rect 53582 704602 63266 704838
rect 63502 704602 63586 704838
rect 63822 704602 73506 704838
rect 73742 704602 73826 704838
rect 74062 704602 83746 704838
rect 83982 704602 84066 704838
rect 84302 704602 93986 704838
rect 94222 704602 94306 704838
rect 94542 704602 104226 704838
rect 104462 704602 104546 704838
rect 104782 704602 114466 704838
rect 114702 704602 114786 704838
rect 115022 704602 124706 704838
rect 124942 704602 125026 704838
rect 125262 704602 134946 704838
rect 135182 704602 135266 704838
rect 135502 704602 145186 704838
rect 145422 704602 145506 704838
rect 145742 704602 155426 704838
rect 155662 704602 155746 704838
rect 155982 704602 165666 704838
rect 165902 704602 165986 704838
rect 166222 704602 175906 704838
rect 176142 704602 176226 704838
rect 176462 704602 186146 704838
rect 186382 704602 186466 704838
rect 186702 704602 196386 704838
rect 196622 704602 196706 704838
rect 196942 704602 206626 704838
rect 206862 704602 206946 704838
rect 207182 704602 216866 704838
rect 217102 704602 217186 704838
rect 217422 704602 227106 704838
rect 227342 704602 227426 704838
rect 227662 704602 237346 704838
rect 237582 704602 237666 704838
rect 237902 704602 247586 704838
rect 247822 704602 247906 704838
rect 248142 704602 257826 704838
rect 258062 704602 258146 704838
rect 258382 704602 268066 704838
rect 268302 704602 268386 704838
rect 268622 704602 278306 704838
rect 278542 704602 278626 704838
rect 278862 704602 288546 704838
rect 288782 704602 288866 704838
rect 289102 704602 298786 704838
rect 299022 704602 299106 704838
rect 299342 704602 309026 704838
rect 309262 704602 309346 704838
rect 309582 704602 319266 704838
rect 319502 704602 319586 704838
rect 319822 704602 329506 704838
rect 329742 704602 329826 704838
rect 330062 704602 339746 704838
rect 339982 704602 340066 704838
rect 340302 704602 349986 704838
rect 350222 704602 350306 704838
rect 350542 704602 360226 704838
rect 360462 704602 360546 704838
rect 360782 704602 370466 704838
rect 370702 704602 370786 704838
rect 371022 704602 380706 704838
rect 380942 704602 381026 704838
rect 381262 704602 390946 704838
rect 391182 704602 391266 704838
rect 391502 704602 401186 704838
rect 401422 704602 401506 704838
rect 401742 704602 411426 704838
rect 411662 704602 411746 704838
rect 411982 704602 421666 704838
rect 421902 704602 421986 704838
rect 422222 704602 431906 704838
rect 432142 704602 432226 704838
rect 432462 704602 442146 704838
rect 442382 704602 442466 704838
rect 442702 704602 452386 704838
rect 452622 704602 452706 704838
rect 452942 704602 462626 704838
rect 462862 704602 462946 704838
rect 463182 704602 472866 704838
rect 473102 704602 473186 704838
rect 473422 704602 483106 704838
rect 483342 704602 483426 704838
rect 483662 704602 493346 704838
rect 493582 704602 493666 704838
rect 493902 704602 503586 704838
rect 503822 704602 503906 704838
rect 504142 704602 513826 704838
rect 514062 704602 514146 704838
rect 514382 704602 524066 704838
rect 524302 704602 524386 704838
rect 524622 704602 534306 704838
rect 534542 704602 534626 704838
rect 534862 704602 544546 704838
rect 544782 704602 544866 704838
rect 545102 704602 554786 704838
rect 555022 704602 555106 704838
rect 555342 704602 565026 704838
rect 565262 704602 565346 704838
rect 565582 704602 575266 704838
rect 575502 704602 575586 704838
rect 575822 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 12066 704518
rect 12302 704282 12386 704518
rect 12622 704282 22306 704518
rect 22542 704282 22626 704518
rect 22862 704282 32546 704518
rect 32782 704282 32866 704518
rect 33102 704282 42786 704518
rect 43022 704282 43106 704518
rect 43342 704282 53026 704518
rect 53262 704282 53346 704518
rect 53582 704282 63266 704518
rect 63502 704282 63586 704518
rect 63822 704282 73506 704518
rect 73742 704282 73826 704518
rect 74062 704282 83746 704518
rect 83982 704282 84066 704518
rect 84302 704282 93986 704518
rect 94222 704282 94306 704518
rect 94542 704282 104226 704518
rect 104462 704282 104546 704518
rect 104782 704282 114466 704518
rect 114702 704282 114786 704518
rect 115022 704282 124706 704518
rect 124942 704282 125026 704518
rect 125262 704282 134946 704518
rect 135182 704282 135266 704518
rect 135502 704282 145186 704518
rect 145422 704282 145506 704518
rect 145742 704282 155426 704518
rect 155662 704282 155746 704518
rect 155982 704282 165666 704518
rect 165902 704282 165986 704518
rect 166222 704282 175906 704518
rect 176142 704282 176226 704518
rect 176462 704282 186146 704518
rect 186382 704282 186466 704518
rect 186702 704282 196386 704518
rect 196622 704282 196706 704518
rect 196942 704282 206626 704518
rect 206862 704282 206946 704518
rect 207182 704282 216866 704518
rect 217102 704282 217186 704518
rect 217422 704282 227106 704518
rect 227342 704282 227426 704518
rect 227662 704282 237346 704518
rect 237582 704282 237666 704518
rect 237902 704282 247586 704518
rect 247822 704282 247906 704518
rect 248142 704282 257826 704518
rect 258062 704282 258146 704518
rect 258382 704282 268066 704518
rect 268302 704282 268386 704518
rect 268622 704282 278306 704518
rect 278542 704282 278626 704518
rect 278862 704282 288546 704518
rect 288782 704282 288866 704518
rect 289102 704282 298786 704518
rect 299022 704282 299106 704518
rect 299342 704282 309026 704518
rect 309262 704282 309346 704518
rect 309582 704282 319266 704518
rect 319502 704282 319586 704518
rect 319822 704282 329506 704518
rect 329742 704282 329826 704518
rect 330062 704282 339746 704518
rect 339982 704282 340066 704518
rect 340302 704282 349986 704518
rect 350222 704282 350306 704518
rect 350542 704282 360226 704518
rect 360462 704282 360546 704518
rect 360782 704282 370466 704518
rect 370702 704282 370786 704518
rect 371022 704282 380706 704518
rect 380942 704282 381026 704518
rect 381262 704282 390946 704518
rect 391182 704282 391266 704518
rect 391502 704282 401186 704518
rect 401422 704282 401506 704518
rect 401742 704282 411426 704518
rect 411662 704282 411746 704518
rect 411982 704282 421666 704518
rect 421902 704282 421986 704518
rect 422222 704282 431906 704518
rect 432142 704282 432226 704518
rect 432462 704282 442146 704518
rect 442382 704282 442466 704518
rect 442702 704282 452386 704518
rect 452622 704282 452706 704518
rect 452942 704282 462626 704518
rect 462862 704282 462946 704518
rect 463182 704282 472866 704518
rect 473102 704282 473186 704518
rect 473422 704282 483106 704518
rect 483342 704282 483426 704518
rect 483662 704282 493346 704518
rect 493582 704282 493666 704518
rect 493902 704282 503586 704518
rect 503822 704282 503906 704518
rect 504142 704282 513826 704518
rect 514062 704282 514146 704518
rect 514382 704282 524066 704518
rect 524302 704282 524386 704518
rect 524622 704282 534306 704518
rect 534542 704282 534626 704518
rect 534862 704282 544546 704518
rect 544782 704282 544866 704518
rect 545102 704282 554786 704518
rect 555022 704282 555106 704518
rect 555342 704282 565026 704518
rect 565262 704282 565346 704518
rect 565582 704282 575266 704518
rect 575502 704282 575586 704518
rect 575822 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 23226 698614
rect 23462 698378 23546 698614
rect 23782 698378 33466 698614
rect 33702 698378 33786 698614
rect 34022 698378 43706 698614
rect 43942 698378 44026 698614
rect 44262 698378 53946 698614
rect 54182 698378 54266 698614
rect 54502 698378 64186 698614
rect 64422 698378 64506 698614
rect 64742 698378 74426 698614
rect 74662 698378 74746 698614
rect 74982 698378 84666 698614
rect 84902 698378 84986 698614
rect 85222 698378 94906 698614
rect 95142 698378 95226 698614
rect 95462 698378 105146 698614
rect 105382 698378 105466 698614
rect 105702 698378 115386 698614
rect 115622 698378 115706 698614
rect 115942 698378 125626 698614
rect 125862 698378 125946 698614
rect 126182 698378 135866 698614
rect 136102 698378 136186 698614
rect 136422 698378 146106 698614
rect 146342 698378 146426 698614
rect 146662 698378 156346 698614
rect 156582 698378 156666 698614
rect 156902 698378 166586 698614
rect 166822 698378 166906 698614
rect 167142 698378 176826 698614
rect 177062 698378 177146 698614
rect 177382 698378 187066 698614
rect 187302 698378 187386 698614
rect 187622 698378 197306 698614
rect 197542 698378 197626 698614
rect 197862 698378 207546 698614
rect 207782 698378 207866 698614
rect 208102 698378 217786 698614
rect 218022 698378 218106 698614
rect 218342 698378 228026 698614
rect 228262 698378 228346 698614
rect 228582 698378 238266 698614
rect 238502 698378 238586 698614
rect 238822 698378 248506 698614
rect 248742 698378 248826 698614
rect 249062 698378 258746 698614
rect 258982 698378 259066 698614
rect 259302 698378 268986 698614
rect 269222 698378 269306 698614
rect 269542 698378 279226 698614
rect 279462 698378 279546 698614
rect 279782 698378 289466 698614
rect 289702 698378 289786 698614
rect 290022 698378 299706 698614
rect 299942 698378 300026 698614
rect 300262 698378 309946 698614
rect 310182 698378 310266 698614
rect 310502 698378 320186 698614
rect 320422 698378 320506 698614
rect 320742 698378 330426 698614
rect 330662 698378 330746 698614
rect 330982 698378 340666 698614
rect 340902 698378 340986 698614
rect 341222 698378 350906 698614
rect 351142 698378 351226 698614
rect 351462 698378 361146 698614
rect 361382 698378 361466 698614
rect 361702 698378 371386 698614
rect 371622 698378 371706 698614
rect 371942 698378 381626 698614
rect 381862 698378 381946 698614
rect 382182 698378 391866 698614
rect 392102 698378 392186 698614
rect 392422 698378 402106 698614
rect 402342 698378 402426 698614
rect 402662 698378 412346 698614
rect 412582 698378 412666 698614
rect 412902 698378 422586 698614
rect 422822 698378 422906 698614
rect 423142 698378 432826 698614
rect 433062 698378 433146 698614
rect 433382 698378 443066 698614
rect 443302 698378 443386 698614
rect 443622 698378 453306 698614
rect 453542 698378 453626 698614
rect 453862 698378 463546 698614
rect 463782 698378 463866 698614
rect 464102 698378 473786 698614
rect 474022 698378 474106 698614
rect 474342 698378 484026 698614
rect 484262 698378 484346 698614
rect 484582 698378 494266 698614
rect 494502 698378 494586 698614
rect 494822 698378 504506 698614
rect 504742 698378 504826 698614
rect 505062 698378 514746 698614
rect 514982 698378 515066 698614
rect 515302 698378 524986 698614
rect 525222 698378 525306 698614
rect 525542 698378 535226 698614
rect 535462 698378 535546 698614
rect 535782 698378 545466 698614
rect 545702 698378 545786 698614
rect 546022 698378 555706 698614
rect 555942 698378 556026 698614
rect 556262 698378 565946 698614
rect 566182 698378 566266 698614
rect 566502 698378 576186 698614
rect 576422 698378 576506 698614
rect 576742 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 23226 698294
rect 23462 698058 23546 698294
rect 23782 698058 33466 698294
rect 33702 698058 33786 698294
rect 34022 698058 43706 698294
rect 43942 698058 44026 698294
rect 44262 698058 53946 698294
rect 54182 698058 54266 698294
rect 54502 698058 64186 698294
rect 64422 698058 64506 698294
rect 64742 698058 74426 698294
rect 74662 698058 74746 698294
rect 74982 698058 84666 698294
rect 84902 698058 84986 698294
rect 85222 698058 94906 698294
rect 95142 698058 95226 698294
rect 95462 698058 105146 698294
rect 105382 698058 105466 698294
rect 105702 698058 115386 698294
rect 115622 698058 115706 698294
rect 115942 698058 125626 698294
rect 125862 698058 125946 698294
rect 126182 698058 135866 698294
rect 136102 698058 136186 698294
rect 136422 698058 146106 698294
rect 146342 698058 146426 698294
rect 146662 698058 156346 698294
rect 156582 698058 156666 698294
rect 156902 698058 166586 698294
rect 166822 698058 166906 698294
rect 167142 698058 176826 698294
rect 177062 698058 177146 698294
rect 177382 698058 187066 698294
rect 187302 698058 187386 698294
rect 187622 698058 197306 698294
rect 197542 698058 197626 698294
rect 197862 698058 207546 698294
rect 207782 698058 207866 698294
rect 208102 698058 217786 698294
rect 218022 698058 218106 698294
rect 218342 698058 228026 698294
rect 228262 698058 228346 698294
rect 228582 698058 238266 698294
rect 238502 698058 238586 698294
rect 238822 698058 248506 698294
rect 248742 698058 248826 698294
rect 249062 698058 258746 698294
rect 258982 698058 259066 698294
rect 259302 698058 268986 698294
rect 269222 698058 269306 698294
rect 269542 698058 279226 698294
rect 279462 698058 279546 698294
rect 279782 698058 289466 698294
rect 289702 698058 289786 698294
rect 290022 698058 299706 698294
rect 299942 698058 300026 698294
rect 300262 698058 309946 698294
rect 310182 698058 310266 698294
rect 310502 698058 320186 698294
rect 320422 698058 320506 698294
rect 320742 698058 330426 698294
rect 330662 698058 330746 698294
rect 330982 698058 340666 698294
rect 340902 698058 340986 698294
rect 341222 698058 350906 698294
rect 351142 698058 351226 698294
rect 351462 698058 361146 698294
rect 361382 698058 361466 698294
rect 361702 698058 371386 698294
rect 371622 698058 371706 698294
rect 371942 698058 381626 698294
rect 381862 698058 381946 698294
rect 382182 698058 391866 698294
rect 392102 698058 392186 698294
rect 392422 698058 402106 698294
rect 402342 698058 402426 698294
rect 402662 698058 412346 698294
rect 412582 698058 412666 698294
rect 412902 698058 422586 698294
rect 422822 698058 422906 698294
rect 423142 698058 432826 698294
rect 433062 698058 433146 698294
rect 433382 698058 443066 698294
rect 443302 698058 443386 698294
rect 443622 698058 453306 698294
rect 453542 698058 453626 698294
rect 453862 698058 463546 698294
rect 463782 698058 463866 698294
rect 464102 698058 473786 698294
rect 474022 698058 474106 698294
rect 474342 698058 484026 698294
rect 484262 698058 484346 698294
rect 484582 698058 494266 698294
rect 494502 698058 494586 698294
rect 494822 698058 504506 698294
rect 504742 698058 504826 698294
rect 505062 698058 514746 698294
rect 514982 698058 515066 698294
rect 515302 698058 524986 698294
rect 525222 698058 525306 698294
rect 525542 698058 535226 698294
rect 535462 698058 535546 698294
rect 535782 698058 545466 698294
rect 545702 698058 545786 698294
rect 546022 698058 555706 698294
rect 555942 698058 556026 698294
rect 556262 698058 565946 698294
rect 566182 698058 566266 698294
rect 566502 698058 576186 698294
rect 576422 698058 576506 698294
rect 576742 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 19506 694894
rect 19742 694658 19826 694894
rect 20062 694658 29746 694894
rect 29982 694658 30066 694894
rect 30302 694658 39986 694894
rect 40222 694658 40306 694894
rect 40542 694658 50226 694894
rect 50462 694658 50546 694894
rect 50782 694658 60466 694894
rect 60702 694658 60786 694894
rect 61022 694658 70706 694894
rect 70942 694658 71026 694894
rect 71262 694658 80946 694894
rect 81182 694658 81266 694894
rect 81502 694658 91186 694894
rect 91422 694658 91506 694894
rect 91742 694658 101426 694894
rect 101662 694658 101746 694894
rect 101982 694658 111666 694894
rect 111902 694658 111986 694894
rect 112222 694658 121906 694894
rect 122142 694658 122226 694894
rect 122462 694658 132146 694894
rect 132382 694658 132466 694894
rect 132702 694658 142386 694894
rect 142622 694658 142706 694894
rect 142942 694658 152626 694894
rect 152862 694658 152946 694894
rect 153182 694658 162866 694894
rect 163102 694658 163186 694894
rect 163422 694658 173106 694894
rect 173342 694658 173426 694894
rect 173662 694658 183346 694894
rect 183582 694658 183666 694894
rect 183902 694658 193586 694894
rect 193822 694658 193906 694894
rect 194142 694658 203826 694894
rect 204062 694658 204146 694894
rect 204382 694658 214066 694894
rect 214302 694658 214386 694894
rect 214622 694658 224306 694894
rect 224542 694658 224626 694894
rect 224862 694658 234546 694894
rect 234782 694658 234866 694894
rect 235102 694658 244786 694894
rect 245022 694658 245106 694894
rect 245342 694658 255026 694894
rect 255262 694658 255346 694894
rect 255582 694658 265266 694894
rect 265502 694658 265586 694894
rect 265822 694658 275506 694894
rect 275742 694658 275826 694894
rect 276062 694658 285746 694894
rect 285982 694658 286066 694894
rect 286302 694658 295986 694894
rect 296222 694658 296306 694894
rect 296542 694658 306226 694894
rect 306462 694658 306546 694894
rect 306782 694658 316466 694894
rect 316702 694658 316786 694894
rect 317022 694658 326706 694894
rect 326942 694658 327026 694894
rect 327262 694658 336946 694894
rect 337182 694658 337266 694894
rect 337502 694658 347186 694894
rect 347422 694658 347506 694894
rect 347742 694658 357426 694894
rect 357662 694658 357746 694894
rect 357982 694658 367666 694894
rect 367902 694658 367986 694894
rect 368222 694658 377906 694894
rect 378142 694658 378226 694894
rect 378462 694658 388146 694894
rect 388382 694658 388466 694894
rect 388702 694658 398386 694894
rect 398622 694658 398706 694894
rect 398942 694658 408626 694894
rect 408862 694658 408946 694894
rect 409182 694658 418866 694894
rect 419102 694658 419186 694894
rect 419422 694658 429106 694894
rect 429342 694658 429426 694894
rect 429662 694658 439346 694894
rect 439582 694658 439666 694894
rect 439902 694658 449586 694894
rect 449822 694658 449906 694894
rect 450142 694658 459826 694894
rect 460062 694658 460146 694894
rect 460382 694658 470066 694894
rect 470302 694658 470386 694894
rect 470622 694658 480306 694894
rect 480542 694658 480626 694894
rect 480862 694658 490546 694894
rect 490782 694658 490866 694894
rect 491102 694658 500786 694894
rect 501022 694658 501106 694894
rect 501342 694658 511026 694894
rect 511262 694658 511346 694894
rect 511582 694658 521266 694894
rect 521502 694658 521586 694894
rect 521822 694658 531506 694894
rect 531742 694658 531826 694894
rect 532062 694658 541746 694894
rect 541982 694658 542066 694894
rect 542302 694658 551986 694894
rect 552222 694658 552306 694894
rect 552542 694658 562226 694894
rect 562462 694658 562546 694894
rect 562782 694658 572466 694894
rect 572702 694658 572786 694894
rect 573022 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 19506 694574
rect 19742 694338 19826 694574
rect 20062 694338 29746 694574
rect 29982 694338 30066 694574
rect 30302 694338 39986 694574
rect 40222 694338 40306 694574
rect 40542 694338 50226 694574
rect 50462 694338 50546 694574
rect 50782 694338 60466 694574
rect 60702 694338 60786 694574
rect 61022 694338 70706 694574
rect 70942 694338 71026 694574
rect 71262 694338 80946 694574
rect 81182 694338 81266 694574
rect 81502 694338 91186 694574
rect 91422 694338 91506 694574
rect 91742 694338 101426 694574
rect 101662 694338 101746 694574
rect 101982 694338 111666 694574
rect 111902 694338 111986 694574
rect 112222 694338 121906 694574
rect 122142 694338 122226 694574
rect 122462 694338 132146 694574
rect 132382 694338 132466 694574
rect 132702 694338 142386 694574
rect 142622 694338 142706 694574
rect 142942 694338 152626 694574
rect 152862 694338 152946 694574
rect 153182 694338 162866 694574
rect 163102 694338 163186 694574
rect 163422 694338 173106 694574
rect 173342 694338 173426 694574
rect 173662 694338 183346 694574
rect 183582 694338 183666 694574
rect 183902 694338 193586 694574
rect 193822 694338 193906 694574
rect 194142 694338 203826 694574
rect 204062 694338 204146 694574
rect 204382 694338 214066 694574
rect 214302 694338 214386 694574
rect 214622 694338 224306 694574
rect 224542 694338 224626 694574
rect 224862 694338 234546 694574
rect 234782 694338 234866 694574
rect 235102 694338 244786 694574
rect 245022 694338 245106 694574
rect 245342 694338 255026 694574
rect 255262 694338 255346 694574
rect 255582 694338 265266 694574
rect 265502 694338 265586 694574
rect 265822 694338 275506 694574
rect 275742 694338 275826 694574
rect 276062 694338 285746 694574
rect 285982 694338 286066 694574
rect 286302 694338 295986 694574
rect 296222 694338 296306 694574
rect 296542 694338 306226 694574
rect 306462 694338 306546 694574
rect 306782 694338 316466 694574
rect 316702 694338 316786 694574
rect 317022 694338 326706 694574
rect 326942 694338 327026 694574
rect 327262 694338 336946 694574
rect 337182 694338 337266 694574
rect 337502 694338 347186 694574
rect 347422 694338 347506 694574
rect 347742 694338 357426 694574
rect 357662 694338 357746 694574
rect 357982 694338 367666 694574
rect 367902 694338 367986 694574
rect 368222 694338 377906 694574
rect 378142 694338 378226 694574
rect 378462 694338 388146 694574
rect 388382 694338 388466 694574
rect 388702 694338 398386 694574
rect 398622 694338 398706 694574
rect 398942 694338 408626 694574
rect 408862 694338 408946 694574
rect 409182 694338 418866 694574
rect 419102 694338 419186 694574
rect 419422 694338 429106 694574
rect 429342 694338 429426 694574
rect 429662 694338 439346 694574
rect 439582 694338 439666 694574
rect 439902 694338 449586 694574
rect 449822 694338 449906 694574
rect 450142 694338 459826 694574
rect 460062 694338 460146 694574
rect 460382 694338 470066 694574
rect 470302 694338 470386 694574
rect 470622 694338 480306 694574
rect 480542 694338 480626 694574
rect 480862 694338 490546 694574
rect 490782 694338 490866 694574
rect 491102 694338 500786 694574
rect 501022 694338 501106 694574
rect 501342 694338 511026 694574
rect 511262 694338 511346 694574
rect 511582 694338 521266 694574
rect 521502 694338 521586 694574
rect 521822 694338 531506 694574
rect 531742 694338 531826 694574
rect 532062 694338 541746 694574
rect 541982 694338 542066 694574
rect 542302 694338 551986 694574
rect 552222 694338 552306 694574
rect 552542 694338 562226 694574
rect 562462 694338 562546 694574
rect 562782 694338 572466 694574
rect 572702 694338 572786 694574
rect 573022 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 15786 691174
rect 16022 690938 16106 691174
rect 16342 690938 26026 691174
rect 26262 690938 26346 691174
rect 26582 690938 36266 691174
rect 36502 690938 36586 691174
rect 36822 690938 46506 691174
rect 46742 690938 46826 691174
rect 47062 690938 56746 691174
rect 56982 690938 57066 691174
rect 57302 690938 66986 691174
rect 67222 690938 67306 691174
rect 67542 690938 77226 691174
rect 77462 690938 77546 691174
rect 77782 690938 87466 691174
rect 87702 690938 87786 691174
rect 88022 690938 97706 691174
rect 97942 690938 98026 691174
rect 98262 690938 107946 691174
rect 108182 690938 108266 691174
rect 108502 690938 118186 691174
rect 118422 690938 118506 691174
rect 118742 690938 128426 691174
rect 128662 690938 128746 691174
rect 128982 690938 138666 691174
rect 138902 690938 138986 691174
rect 139222 690938 148906 691174
rect 149142 690938 149226 691174
rect 149462 690938 159146 691174
rect 159382 690938 159466 691174
rect 159702 690938 169386 691174
rect 169622 690938 169706 691174
rect 169942 690938 179626 691174
rect 179862 690938 179946 691174
rect 180182 690938 189866 691174
rect 190102 690938 190186 691174
rect 190422 690938 200106 691174
rect 200342 690938 200426 691174
rect 200662 690938 210346 691174
rect 210582 690938 210666 691174
rect 210902 690938 220586 691174
rect 220822 690938 220906 691174
rect 221142 690938 230826 691174
rect 231062 690938 231146 691174
rect 231382 690938 241066 691174
rect 241302 690938 241386 691174
rect 241622 690938 251306 691174
rect 251542 690938 251626 691174
rect 251862 690938 261546 691174
rect 261782 690938 261866 691174
rect 262102 690938 271786 691174
rect 272022 690938 272106 691174
rect 272342 690938 282026 691174
rect 282262 690938 282346 691174
rect 282582 690938 292266 691174
rect 292502 690938 292586 691174
rect 292822 690938 302506 691174
rect 302742 690938 302826 691174
rect 303062 690938 312746 691174
rect 312982 690938 313066 691174
rect 313302 690938 322986 691174
rect 323222 690938 323306 691174
rect 323542 690938 333226 691174
rect 333462 690938 333546 691174
rect 333782 690938 343466 691174
rect 343702 690938 343786 691174
rect 344022 690938 353706 691174
rect 353942 690938 354026 691174
rect 354262 690938 363946 691174
rect 364182 690938 364266 691174
rect 364502 690938 374186 691174
rect 374422 690938 374506 691174
rect 374742 690938 384426 691174
rect 384662 690938 384746 691174
rect 384982 690938 394666 691174
rect 394902 690938 394986 691174
rect 395222 690938 404906 691174
rect 405142 690938 405226 691174
rect 405462 690938 415146 691174
rect 415382 690938 415466 691174
rect 415702 690938 425386 691174
rect 425622 690938 425706 691174
rect 425942 690938 435626 691174
rect 435862 690938 435946 691174
rect 436182 690938 445866 691174
rect 446102 690938 446186 691174
rect 446422 690938 456106 691174
rect 456342 690938 456426 691174
rect 456662 690938 466346 691174
rect 466582 690938 466666 691174
rect 466902 690938 476586 691174
rect 476822 690938 476906 691174
rect 477142 690938 486826 691174
rect 487062 690938 487146 691174
rect 487382 690938 497066 691174
rect 497302 690938 497386 691174
rect 497622 690938 507306 691174
rect 507542 690938 507626 691174
rect 507862 690938 517546 691174
rect 517782 690938 517866 691174
rect 518102 690938 527786 691174
rect 528022 690938 528106 691174
rect 528342 690938 538026 691174
rect 538262 690938 538346 691174
rect 538582 690938 548266 691174
rect 548502 690938 548586 691174
rect 548822 690938 558506 691174
rect 558742 690938 558826 691174
rect 559062 690938 568746 691174
rect 568982 690938 569066 691174
rect 569302 690938 578986 691174
rect 579222 690938 579306 691174
rect 579542 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 15786 690854
rect 16022 690618 16106 690854
rect 16342 690618 26026 690854
rect 26262 690618 26346 690854
rect 26582 690618 36266 690854
rect 36502 690618 36586 690854
rect 36822 690618 46506 690854
rect 46742 690618 46826 690854
rect 47062 690618 56746 690854
rect 56982 690618 57066 690854
rect 57302 690618 66986 690854
rect 67222 690618 67306 690854
rect 67542 690618 77226 690854
rect 77462 690618 77546 690854
rect 77782 690618 87466 690854
rect 87702 690618 87786 690854
rect 88022 690618 97706 690854
rect 97942 690618 98026 690854
rect 98262 690618 107946 690854
rect 108182 690618 108266 690854
rect 108502 690618 118186 690854
rect 118422 690618 118506 690854
rect 118742 690618 128426 690854
rect 128662 690618 128746 690854
rect 128982 690618 138666 690854
rect 138902 690618 138986 690854
rect 139222 690618 148906 690854
rect 149142 690618 149226 690854
rect 149462 690618 159146 690854
rect 159382 690618 159466 690854
rect 159702 690618 169386 690854
rect 169622 690618 169706 690854
rect 169942 690618 179626 690854
rect 179862 690618 179946 690854
rect 180182 690618 189866 690854
rect 190102 690618 190186 690854
rect 190422 690618 200106 690854
rect 200342 690618 200426 690854
rect 200662 690618 210346 690854
rect 210582 690618 210666 690854
rect 210902 690618 220586 690854
rect 220822 690618 220906 690854
rect 221142 690618 230826 690854
rect 231062 690618 231146 690854
rect 231382 690618 241066 690854
rect 241302 690618 241386 690854
rect 241622 690618 251306 690854
rect 251542 690618 251626 690854
rect 251862 690618 261546 690854
rect 261782 690618 261866 690854
rect 262102 690618 271786 690854
rect 272022 690618 272106 690854
rect 272342 690618 282026 690854
rect 282262 690618 282346 690854
rect 282582 690618 292266 690854
rect 292502 690618 292586 690854
rect 292822 690618 302506 690854
rect 302742 690618 302826 690854
rect 303062 690618 312746 690854
rect 312982 690618 313066 690854
rect 313302 690618 322986 690854
rect 323222 690618 323306 690854
rect 323542 690618 333226 690854
rect 333462 690618 333546 690854
rect 333782 690618 343466 690854
rect 343702 690618 343786 690854
rect 344022 690618 353706 690854
rect 353942 690618 354026 690854
rect 354262 690618 363946 690854
rect 364182 690618 364266 690854
rect 364502 690618 374186 690854
rect 374422 690618 374506 690854
rect 374742 690618 384426 690854
rect 384662 690618 384746 690854
rect 384982 690618 394666 690854
rect 394902 690618 394986 690854
rect 395222 690618 404906 690854
rect 405142 690618 405226 690854
rect 405462 690618 415146 690854
rect 415382 690618 415466 690854
rect 415702 690618 425386 690854
rect 425622 690618 425706 690854
rect 425942 690618 435626 690854
rect 435862 690618 435946 690854
rect 436182 690618 445866 690854
rect 446102 690618 446186 690854
rect 446422 690618 456106 690854
rect 456342 690618 456426 690854
rect 456662 690618 466346 690854
rect 466582 690618 466666 690854
rect 466902 690618 476586 690854
rect 476822 690618 476906 690854
rect 477142 690618 486826 690854
rect 487062 690618 487146 690854
rect 487382 690618 497066 690854
rect 497302 690618 497386 690854
rect 497622 690618 507306 690854
rect 507542 690618 507626 690854
rect 507862 690618 517546 690854
rect 517782 690618 517866 690854
rect 518102 690618 527786 690854
rect 528022 690618 528106 690854
rect 528342 690618 538026 690854
rect 538262 690618 538346 690854
rect 538582 690618 548266 690854
rect 548502 690618 548586 690854
rect 548822 690618 558506 690854
rect 558742 690618 558826 690854
rect 559062 690618 568746 690854
rect 568982 690618 569066 690854
rect 569302 690618 578986 690854
rect 579222 690618 579306 690854
rect 579542 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 12066 687454
rect 12302 687218 12386 687454
rect 12622 687218 22306 687454
rect 22542 687218 22626 687454
rect 22862 687218 32546 687454
rect 32782 687218 32866 687454
rect 33102 687218 42786 687454
rect 43022 687218 43106 687454
rect 43342 687218 53026 687454
rect 53262 687218 53346 687454
rect 53582 687218 63266 687454
rect 63502 687218 63586 687454
rect 63822 687218 73506 687454
rect 73742 687218 73826 687454
rect 74062 687218 83746 687454
rect 83982 687218 84066 687454
rect 84302 687218 93986 687454
rect 94222 687218 94306 687454
rect 94542 687218 104226 687454
rect 104462 687218 104546 687454
rect 104782 687218 114466 687454
rect 114702 687218 114786 687454
rect 115022 687218 124706 687454
rect 124942 687218 125026 687454
rect 125262 687218 134946 687454
rect 135182 687218 135266 687454
rect 135502 687218 145186 687454
rect 145422 687218 145506 687454
rect 145742 687218 155426 687454
rect 155662 687218 155746 687454
rect 155982 687218 165666 687454
rect 165902 687218 165986 687454
rect 166222 687218 175906 687454
rect 176142 687218 176226 687454
rect 176462 687218 186146 687454
rect 186382 687218 186466 687454
rect 186702 687218 196386 687454
rect 196622 687218 196706 687454
rect 196942 687218 206626 687454
rect 206862 687218 206946 687454
rect 207182 687218 216866 687454
rect 217102 687218 217186 687454
rect 217422 687218 227106 687454
rect 227342 687218 227426 687454
rect 227662 687218 237346 687454
rect 237582 687218 237666 687454
rect 237902 687218 247586 687454
rect 247822 687218 247906 687454
rect 248142 687218 257826 687454
rect 258062 687218 258146 687454
rect 258382 687218 268066 687454
rect 268302 687218 268386 687454
rect 268622 687218 278306 687454
rect 278542 687218 278626 687454
rect 278862 687218 288546 687454
rect 288782 687218 288866 687454
rect 289102 687218 298786 687454
rect 299022 687218 299106 687454
rect 299342 687218 309026 687454
rect 309262 687218 309346 687454
rect 309582 687218 319266 687454
rect 319502 687218 319586 687454
rect 319822 687218 329506 687454
rect 329742 687218 329826 687454
rect 330062 687218 339746 687454
rect 339982 687218 340066 687454
rect 340302 687218 349986 687454
rect 350222 687218 350306 687454
rect 350542 687218 360226 687454
rect 360462 687218 360546 687454
rect 360782 687218 370466 687454
rect 370702 687218 370786 687454
rect 371022 687218 380706 687454
rect 380942 687218 381026 687454
rect 381262 687218 390946 687454
rect 391182 687218 391266 687454
rect 391502 687218 401186 687454
rect 401422 687218 401506 687454
rect 401742 687218 411426 687454
rect 411662 687218 411746 687454
rect 411982 687218 421666 687454
rect 421902 687218 421986 687454
rect 422222 687218 431906 687454
rect 432142 687218 432226 687454
rect 432462 687218 442146 687454
rect 442382 687218 442466 687454
rect 442702 687218 452386 687454
rect 452622 687218 452706 687454
rect 452942 687218 462626 687454
rect 462862 687218 462946 687454
rect 463182 687218 472866 687454
rect 473102 687218 473186 687454
rect 473422 687218 483106 687454
rect 483342 687218 483426 687454
rect 483662 687218 493346 687454
rect 493582 687218 493666 687454
rect 493902 687218 503586 687454
rect 503822 687218 503906 687454
rect 504142 687218 513826 687454
rect 514062 687218 514146 687454
rect 514382 687218 524066 687454
rect 524302 687218 524386 687454
rect 524622 687218 534306 687454
rect 534542 687218 534626 687454
rect 534862 687218 544546 687454
rect 544782 687218 544866 687454
rect 545102 687218 554786 687454
rect 555022 687218 555106 687454
rect 555342 687218 565026 687454
rect 565262 687218 565346 687454
rect 565582 687218 575266 687454
rect 575502 687218 575586 687454
rect 575822 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 12066 687134
rect 12302 686898 12386 687134
rect 12622 686898 22306 687134
rect 22542 686898 22626 687134
rect 22862 686898 32546 687134
rect 32782 686898 32866 687134
rect 33102 686898 42786 687134
rect 43022 686898 43106 687134
rect 43342 686898 53026 687134
rect 53262 686898 53346 687134
rect 53582 686898 63266 687134
rect 63502 686898 63586 687134
rect 63822 686898 73506 687134
rect 73742 686898 73826 687134
rect 74062 686898 83746 687134
rect 83982 686898 84066 687134
rect 84302 686898 93986 687134
rect 94222 686898 94306 687134
rect 94542 686898 104226 687134
rect 104462 686898 104546 687134
rect 104782 686898 114466 687134
rect 114702 686898 114786 687134
rect 115022 686898 124706 687134
rect 124942 686898 125026 687134
rect 125262 686898 134946 687134
rect 135182 686898 135266 687134
rect 135502 686898 145186 687134
rect 145422 686898 145506 687134
rect 145742 686898 155426 687134
rect 155662 686898 155746 687134
rect 155982 686898 165666 687134
rect 165902 686898 165986 687134
rect 166222 686898 175906 687134
rect 176142 686898 176226 687134
rect 176462 686898 186146 687134
rect 186382 686898 186466 687134
rect 186702 686898 196386 687134
rect 196622 686898 196706 687134
rect 196942 686898 206626 687134
rect 206862 686898 206946 687134
rect 207182 686898 216866 687134
rect 217102 686898 217186 687134
rect 217422 686898 227106 687134
rect 227342 686898 227426 687134
rect 227662 686898 237346 687134
rect 237582 686898 237666 687134
rect 237902 686898 247586 687134
rect 247822 686898 247906 687134
rect 248142 686898 257826 687134
rect 258062 686898 258146 687134
rect 258382 686898 268066 687134
rect 268302 686898 268386 687134
rect 268622 686898 278306 687134
rect 278542 686898 278626 687134
rect 278862 686898 288546 687134
rect 288782 686898 288866 687134
rect 289102 686898 298786 687134
rect 299022 686898 299106 687134
rect 299342 686898 309026 687134
rect 309262 686898 309346 687134
rect 309582 686898 319266 687134
rect 319502 686898 319586 687134
rect 319822 686898 329506 687134
rect 329742 686898 329826 687134
rect 330062 686898 339746 687134
rect 339982 686898 340066 687134
rect 340302 686898 349986 687134
rect 350222 686898 350306 687134
rect 350542 686898 360226 687134
rect 360462 686898 360546 687134
rect 360782 686898 370466 687134
rect 370702 686898 370786 687134
rect 371022 686898 380706 687134
rect 380942 686898 381026 687134
rect 381262 686898 390946 687134
rect 391182 686898 391266 687134
rect 391502 686898 401186 687134
rect 401422 686898 401506 687134
rect 401742 686898 411426 687134
rect 411662 686898 411746 687134
rect 411982 686898 421666 687134
rect 421902 686898 421986 687134
rect 422222 686898 431906 687134
rect 432142 686898 432226 687134
rect 432462 686898 442146 687134
rect 442382 686898 442466 687134
rect 442702 686898 452386 687134
rect 452622 686898 452706 687134
rect 452942 686898 462626 687134
rect 462862 686898 462946 687134
rect 463182 686898 472866 687134
rect 473102 686898 473186 687134
rect 473422 686898 483106 687134
rect 483342 686898 483426 687134
rect 483662 686898 493346 687134
rect 493582 686898 493666 687134
rect 493902 686898 503586 687134
rect 503822 686898 503906 687134
rect 504142 686898 513826 687134
rect 514062 686898 514146 687134
rect 514382 686898 524066 687134
rect 524302 686898 524386 687134
rect 524622 686898 534306 687134
rect 534542 686898 534626 687134
rect 534862 686898 544546 687134
rect 544782 686898 544866 687134
rect 545102 686898 554786 687134
rect 555022 686898 555106 687134
rect 555342 686898 565026 687134
rect 565262 686898 565346 687134
rect 565582 686898 575266 687134
rect 575502 686898 575586 687134
rect 575822 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 18106 680614
rect 18342 680378 18426 680614
rect 18662 680378 28346 680614
rect 28582 680378 28666 680614
rect 28902 680378 38586 680614
rect 38822 680378 38906 680614
rect 39142 680378 48826 680614
rect 49062 680378 49146 680614
rect 49382 680378 59066 680614
rect 59302 680378 59386 680614
rect 59622 680378 69306 680614
rect 69542 680378 69626 680614
rect 69862 680378 79546 680614
rect 79782 680378 79866 680614
rect 80102 680378 89786 680614
rect 90022 680378 90106 680614
rect 90342 680378 100026 680614
rect 100262 680378 100346 680614
rect 100582 680378 110266 680614
rect 110502 680378 110586 680614
rect 110822 680378 120506 680614
rect 120742 680378 120826 680614
rect 121062 680378 130746 680614
rect 130982 680378 131066 680614
rect 131302 680378 140986 680614
rect 141222 680378 141306 680614
rect 141542 680378 151226 680614
rect 151462 680378 151546 680614
rect 151782 680378 161466 680614
rect 161702 680378 161786 680614
rect 162022 680378 171706 680614
rect 171942 680378 172026 680614
rect 172262 680378 181946 680614
rect 182182 680378 182266 680614
rect 182502 680378 192186 680614
rect 192422 680378 192506 680614
rect 192742 680378 202426 680614
rect 202662 680378 202746 680614
rect 202982 680378 212666 680614
rect 212902 680378 212986 680614
rect 213222 680378 222906 680614
rect 223142 680378 223226 680614
rect 223462 680378 233146 680614
rect 233382 680378 233466 680614
rect 233702 680378 243386 680614
rect 243622 680378 243706 680614
rect 243942 680378 253626 680614
rect 253862 680378 253946 680614
rect 254182 680378 263866 680614
rect 264102 680378 264186 680614
rect 264422 680378 274106 680614
rect 274342 680378 274426 680614
rect 274662 680378 284346 680614
rect 284582 680378 284666 680614
rect 284902 680378 294586 680614
rect 294822 680378 294906 680614
rect 295142 680378 304826 680614
rect 305062 680378 305146 680614
rect 305382 680378 315066 680614
rect 315302 680378 315386 680614
rect 315622 680378 325306 680614
rect 325542 680378 325626 680614
rect 325862 680378 335546 680614
rect 335782 680378 335866 680614
rect 336102 680378 345786 680614
rect 346022 680378 346106 680614
rect 346342 680378 356026 680614
rect 356262 680378 356346 680614
rect 356582 680378 366266 680614
rect 366502 680378 366586 680614
rect 366822 680378 376506 680614
rect 376742 680378 376826 680614
rect 377062 680378 386746 680614
rect 386982 680378 387066 680614
rect 387302 680378 396986 680614
rect 397222 680378 397306 680614
rect 397542 680378 407226 680614
rect 407462 680378 407546 680614
rect 407782 680378 417466 680614
rect 417702 680378 417786 680614
rect 418022 680378 427706 680614
rect 427942 680378 428026 680614
rect 428262 680378 437946 680614
rect 438182 680378 438266 680614
rect 438502 680378 448186 680614
rect 448422 680378 448506 680614
rect 448742 680378 458426 680614
rect 458662 680378 458746 680614
rect 458982 680378 468666 680614
rect 468902 680378 468986 680614
rect 469222 680378 478906 680614
rect 479142 680378 479226 680614
rect 479462 680378 489146 680614
rect 489382 680378 489466 680614
rect 489702 680378 499386 680614
rect 499622 680378 499706 680614
rect 499942 680378 509626 680614
rect 509862 680378 509946 680614
rect 510182 680378 519866 680614
rect 520102 680378 520186 680614
rect 520422 680378 530106 680614
rect 530342 680378 530426 680614
rect 530662 680378 540346 680614
rect 540582 680378 540666 680614
rect 540902 680378 550586 680614
rect 550822 680378 550906 680614
rect 551142 680378 560826 680614
rect 561062 680378 561146 680614
rect 561382 680378 571066 680614
rect 571302 680378 571386 680614
rect 571622 680378 581306 680614
rect 581542 680378 581626 680614
rect 581862 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 18106 680294
rect 18342 680058 18426 680294
rect 18662 680058 28346 680294
rect 28582 680058 28666 680294
rect 28902 680058 38586 680294
rect 38822 680058 38906 680294
rect 39142 680058 48826 680294
rect 49062 680058 49146 680294
rect 49382 680058 59066 680294
rect 59302 680058 59386 680294
rect 59622 680058 69306 680294
rect 69542 680058 69626 680294
rect 69862 680058 79546 680294
rect 79782 680058 79866 680294
rect 80102 680058 89786 680294
rect 90022 680058 90106 680294
rect 90342 680058 100026 680294
rect 100262 680058 100346 680294
rect 100582 680058 110266 680294
rect 110502 680058 110586 680294
rect 110822 680058 120506 680294
rect 120742 680058 120826 680294
rect 121062 680058 130746 680294
rect 130982 680058 131066 680294
rect 131302 680058 140986 680294
rect 141222 680058 141306 680294
rect 141542 680058 151226 680294
rect 151462 680058 151546 680294
rect 151782 680058 161466 680294
rect 161702 680058 161786 680294
rect 162022 680058 171706 680294
rect 171942 680058 172026 680294
rect 172262 680058 181946 680294
rect 182182 680058 182266 680294
rect 182502 680058 192186 680294
rect 192422 680058 192506 680294
rect 192742 680058 202426 680294
rect 202662 680058 202746 680294
rect 202982 680058 212666 680294
rect 212902 680058 212986 680294
rect 213222 680058 222906 680294
rect 223142 680058 223226 680294
rect 223462 680058 233146 680294
rect 233382 680058 233466 680294
rect 233702 680058 243386 680294
rect 243622 680058 243706 680294
rect 243942 680058 253626 680294
rect 253862 680058 253946 680294
rect 254182 680058 263866 680294
rect 264102 680058 264186 680294
rect 264422 680058 274106 680294
rect 274342 680058 274426 680294
rect 274662 680058 284346 680294
rect 284582 680058 284666 680294
rect 284902 680058 294586 680294
rect 294822 680058 294906 680294
rect 295142 680058 304826 680294
rect 305062 680058 305146 680294
rect 305382 680058 315066 680294
rect 315302 680058 315386 680294
rect 315622 680058 325306 680294
rect 325542 680058 325626 680294
rect 325862 680058 335546 680294
rect 335782 680058 335866 680294
rect 336102 680058 345786 680294
rect 346022 680058 346106 680294
rect 346342 680058 356026 680294
rect 356262 680058 356346 680294
rect 356582 680058 366266 680294
rect 366502 680058 366586 680294
rect 366822 680058 376506 680294
rect 376742 680058 376826 680294
rect 377062 680058 386746 680294
rect 386982 680058 387066 680294
rect 387302 680058 396986 680294
rect 397222 680058 397306 680294
rect 397542 680058 407226 680294
rect 407462 680058 407546 680294
rect 407782 680058 417466 680294
rect 417702 680058 417786 680294
rect 418022 680058 427706 680294
rect 427942 680058 428026 680294
rect 428262 680058 437946 680294
rect 438182 680058 438266 680294
rect 438502 680058 448186 680294
rect 448422 680058 448506 680294
rect 448742 680058 458426 680294
rect 458662 680058 458746 680294
rect 458982 680058 468666 680294
rect 468902 680058 468986 680294
rect 469222 680058 478906 680294
rect 479142 680058 479226 680294
rect 479462 680058 489146 680294
rect 489382 680058 489466 680294
rect 489702 680058 499386 680294
rect 499622 680058 499706 680294
rect 499942 680058 509626 680294
rect 509862 680058 509946 680294
rect 510182 680058 519866 680294
rect 520102 680058 520186 680294
rect 520422 680058 530106 680294
rect 530342 680058 530426 680294
rect 530662 680058 540346 680294
rect 540582 680058 540666 680294
rect 540902 680058 550586 680294
rect 550822 680058 550906 680294
rect 551142 680058 560826 680294
rect 561062 680058 561146 680294
rect 561382 680058 571066 680294
rect 571302 680058 571386 680294
rect 571622 680058 581306 680294
rect 581542 680058 581626 680294
rect 581862 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 14386 676894
rect 14622 676658 14706 676894
rect 14942 676658 24626 676894
rect 24862 676658 24946 676894
rect 25182 676658 34866 676894
rect 35102 676658 35186 676894
rect 35422 676658 45106 676894
rect 45342 676658 45426 676894
rect 45662 676658 55346 676894
rect 55582 676658 55666 676894
rect 55902 676658 65586 676894
rect 65822 676658 65906 676894
rect 66142 676658 75826 676894
rect 76062 676658 76146 676894
rect 76382 676658 86066 676894
rect 86302 676658 86386 676894
rect 86622 676658 96306 676894
rect 96542 676658 96626 676894
rect 96862 676658 106546 676894
rect 106782 676658 106866 676894
rect 107102 676658 116786 676894
rect 117022 676658 117106 676894
rect 117342 676658 127026 676894
rect 127262 676658 127346 676894
rect 127582 676658 137266 676894
rect 137502 676658 137586 676894
rect 137822 676658 147506 676894
rect 147742 676658 147826 676894
rect 148062 676658 157746 676894
rect 157982 676658 158066 676894
rect 158302 676658 167986 676894
rect 168222 676658 168306 676894
rect 168542 676658 178226 676894
rect 178462 676658 178546 676894
rect 178782 676658 188466 676894
rect 188702 676658 188786 676894
rect 189022 676658 198706 676894
rect 198942 676658 199026 676894
rect 199262 676658 208946 676894
rect 209182 676658 209266 676894
rect 209502 676658 219186 676894
rect 219422 676658 219506 676894
rect 219742 676658 229426 676894
rect 229662 676658 229746 676894
rect 229982 676658 239666 676894
rect 239902 676658 239986 676894
rect 240222 676658 249906 676894
rect 250142 676658 250226 676894
rect 250462 676658 260146 676894
rect 260382 676658 260466 676894
rect 260702 676658 270386 676894
rect 270622 676658 270706 676894
rect 270942 676658 280626 676894
rect 280862 676658 280946 676894
rect 281182 676658 290866 676894
rect 291102 676658 291186 676894
rect 291422 676658 301106 676894
rect 301342 676658 301426 676894
rect 301662 676658 311346 676894
rect 311582 676658 311666 676894
rect 311902 676658 321586 676894
rect 321822 676658 321906 676894
rect 322142 676658 331826 676894
rect 332062 676658 332146 676894
rect 332382 676658 342066 676894
rect 342302 676658 342386 676894
rect 342622 676658 352306 676894
rect 352542 676658 352626 676894
rect 352862 676658 362546 676894
rect 362782 676658 362866 676894
rect 363102 676658 372786 676894
rect 373022 676658 373106 676894
rect 373342 676658 383026 676894
rect 383262 676658 383346 676894
rect 383582 676658 393266 676894
rect 393502 676658 393586 676894
rect 393822 676658 403506 676894
rect 403742 676658 403826 676894
rect 404062 676658 413746 676894
rect 413982 676658 414066 676894
rect 414302 676658 423986 676894
rect 424222 676658 424306 676894
rect 424542 676658 434226 676894
rect 434462 676658 434546 676894
rect 434782 676658 444466 676894
rect 444702 676658 444786 676894
rect 445022 676658 454706 676894
rect 454942 676658 455026 676894
rect 455262 676658 464946 676894
rect 465182 676658 465266 676894
rect 465502 676658 475186 676894
rect 475422 676658 475506 676894
rect 475742 676658 485426 676894
rect 485662 676658 485746 676894
rect 485982 676658 495666 676894
rect 495902 676658 495986 676894
rect 496222 676658 505906 676894
rect 506142 676658 506226 676894
rect 506462 676658 516146 676894
rect 516382 676658 516466 676894
rect 516702 676658 526386 676894
rect 526622 676658 526706 676894
rect 526942 676658 536626 676894
rect 536862 676658 536946 676894
rect 537182 676658 546866 676894
rect 547102 676658 547186 676894
rect 547422 676658 557106 676894
rect 557342 676658 557426 676894
rect 557662 676658 567346 676894
rect 567582 676658 567666 676894
rect 567902 676658 577586 676894
rect 577822 676658 577906 676894
rect 578142 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 14386 676574
rect 14622 676338 14706 676574
rect 14942 676338 24626 676574
rect 24862 676338 24946 676574
rect 25182 676338 34866 676574
rect 35102 676338 35186 676574
rect 35422 676338 45106 676574
rect 45342 676338 45426 676574
rect 45662 676338 55346 676574
rect 55582 676338 55666 676574
rect 55902 676338 65586 676574
rect 65822 676338 65906 676574
rect 66142 676338 75826 676574
rect 76062 676338 76146 676574
rect 76382 676338 86066 676574
rect 86302 676338 86386 676574
rect 86622 676338 96306 676574
rect 96542 676338 96626 676574
rect 96862 676338 106546 676574
rect 106782 676338 106866 676574
rect 107102 676338 116786 676574
rect 117022 676338 117106 676574
rect 117342 676338 127026 676574
rect 127262 676338 127346 676574
rect 127582 676338 137266 676574
rect 137502 676338 137586 676574
rect 137822 676338 147506 676574
rect 147742 676338 147826 676574
rect 148062 676338 157746 676574
rect 157982 676338 158066 676574
rect 158302 676338 167986 676574
rect 168222 676338 168306 676574
rect 168542 676338 178226 676574
rect 178462 676338 178546 676574
rect 178782 676338 188466 676574
rect 188702 676338 188786 676574
rect 189022 676338 198706 676574
rect 198942 676338 199026 676574
rect 199262 676338 208946 676574
rect 209182 676338 209266 676574
rect 209502 676338 219186 676574
rect 219422 676338 219506 676574
rect 219742 676338 229426 676574
rect 229662 676338 229746 676574
rect 229982 676338 239666 676574
rect 239902 676338 239986 676574
rect 240222 676338 249906 676574
rect 250142 676338 250226 676574
rect 250462 676338 260146 676574
rect 260382 676338 260466 676574
rect 260702 676338 270386 676574
rect 270622 676338 270706 676574
rect 270942 676338 280626 676574
rect 280862 676338 280946 676574
rect 281182 676338 290866 676574
rect 291102 676338 291186 676574
rect 291422 676338 301106 676574
rect 301342 676338 301426 676574
rect 301662 676338 311346 676574
rect 311582 676338 311666 676574
rect 311902 676338 321586 676574
rect 321822 676338 321906 676574
rect 322142 676338 331826 676574
rect 332062 676338 332146 676574
rect 332382 676338 342066 676574
rect 342302 676338 342386 676574
rect 342622 676338 352306 676574
rect 352542 676338 352626 676574
rect 352862 676338 362546 676574
rect 362782 676338 362866 676574
rect 363102 676338 372786 676574
rect 373022 676338 373106 676574
rect 373342 676338 383026 676574
rect 383262 676338 383346 676574
rect 383582 676338 393266 676574
rect 393502 676338 393586 676574
rect 393822 676338 403506 676574
rect 403742 676338 403826 676574
rect 404062 676338 413746 676574
rect 413982 676338 414066 676574
rect 414302 676338 423986 676574
rect 424222 676338 424306 676574
rect 424542 676338 434226 676574
rect 434462 676338 434546 676574
rect 434782 676338 444466 676574
rect 444702 676338 444786 676574
rect 445022 676338 454706 676574
rect 454942 676338 455026 676574
rect 455262 676338 464946 676574
rect 465182 676338 465266 676574
rect 465502 676338 475186 676574
rect 475422 676338 475506 676574
rect 475742 676338 485426 676574
rect 485662 676338 485746 676574
rect 485982 676338 495666 676574
rect 495902 676338 495986 676574
rect 496222 676338 505906 676574
rect 506142 676338 506226 676574
rect 506462 676338 516146 676574
rect 516382 676338 516466 676574
rect 516702 676338 526386 676574
rect 526622 676338 526706 676574
rect 526942 676338 536626 676574
rect 536862 676338 536946 676574
rect 537182 676338 546866 676574
rect 547102 676338 547186 676574
rect 547422 676338 557106 676574
rect 557342 676338 557426 676574
rect 557662 676338 567346 676574
rect 567582 676338 567666 676574
rect 567902 676338 577586 676574
rect 577822 676338 577906 676574
rect 578142 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 10666 673174
rect 10902 672938 10986 673174
rect 11222 672938 20906 673174
rect 21142 672938 21226 673174
rect 21462 672938 31146 673174
rect 31382 672938 31466 673174
rect 31702 672938 41386 673174
rect 41622 672938 41706 673174
rect 41942 672938 51626 673174
rect 51862 672938 51946 673174
rect 52182 672938 61866 673174
rect 62102 672938 62186 673174
rect 62422 672938 72106 673174
rect 72342 672938 72426 673174
rect 72662 672938 82346 673174
rect 82582 672938 82666 673174
rect 82902 672938 92586 673174
rect 92822 672938 92906 673174
rect 93142 672938 102826 673174
rect 103062 672938 103146 673174
rect 103382 672938 113066 673174
rect 113302 672938 113386 673174
rect 113622 672938 123306 673174
rect 123542 672938 123626 673174
rect 123862 672938 133546 673174
rect 133782 672938 133866 673174
rect 134102 672938 143786 673174
rect 144022 672938 144106 673174
rect 144342 672938 154026 673174
rect 154262 672938 154346 673174
rect 154582 672938 164266 673174
rect 164502 672938 164586 673174
rect 164822 672938 174506 673174
rect 174742 672938 174826 673174
rect 175062 672938 184746 673174
rect 184982 672938 185066 673174
rect 185302 672938 194986 673174
rect 195222 672938 195306 673174
rect 195542 672938 205226 673174
rect 205462 672938 205546 673174
rect 205782 672938 215466 673174
rect 215702 672938 215786 673174
rect 216022 672938 225706 673174
rect 225942 672938 226026 673174
rect 226262 672938 235946 673174
rect 236182 672938 236266 673174
rect 236502 672938 246186 673174
rect 246422 672938 246506 673174
rect 246742 672938 256426 673174
rect 256662 672938 256746 673174
rect 256982 672938 266666 673174
rect 266902 672938 266986 673174
rect 267222 672938 276906 673174
rect 277142 672938 277226 673174
rect 277462 672938 287146 673174
rect 287382 672938 287466 673174
rect 287702 672938 297386 673174
rect 297622 672938 297706 673174
rect 297942 672938 307626 673174
rect 307862 672938 307946 673174
rect 308182 672938 317866 673174
rect 318102 672938 318186 673174
rect 318422 672938 328106 673174
rect 328342 672938 328426 673174
rect 328662 672938 338346 673174
rect 338582 672938 338666 673174
rect 338902 672938 348586 673174
rect 348822 672938 348906 673174
rect 349142 672938 358826 673174
rect 359062 672938 359146 673174
rect 359382 672938 369066 673174
rect 369302 672938 369386 673174
rect 369622 672938 379306 673174
rect 379542 672938 379626 673174
rect 379862 672938 389546 673174
rect 389782 672938 389866 673174
rect 390102 672938 399786 673174
rect 400022 672938 400106 673174
rect 400342 672938 410026 673174
rect 410262 672938 410346 673174
rect 410582 672938 420266 673174
rect 420502 672938 420586 673174
rect 420822 672938 430506 673174
rect 430742 672938 430826 673174
rect 431062 672938 440746 673174
rect 440982 672938 441066 673174
rect 441302 672938 450986 673174
rect 451222 672938 451306 673174
rect 451542 672938 461226 673174
rect 461462 672938 461546 673174
rect 461782 672938 471466 673174
rect 471702 672938 471786 673174
rect 472022 672938 481706 673174
rect 481942 672938 482026 673174
rect 482262 672938 491946 673174
rect 492182 672938 492266 673174
rect 492502 672938 502186 673174
rect 502422 672938 502506 673174
rect 502742 672938 512426 673174
rect 512662 672938 512746 673174
rect 512982 672938 522666 673174
rect 522902 672938 522986 673174
rect 523222 672938 532906 673174
rect 533142 672938 533226 673174
rect 533462 672938 543146 673174
rect 543382 672938 543466 673174
rect 543702 672938 553386 673174
rect 553622 672938 553706 673174
rect 553942 672938 563626 673174
rect 563862 672938 563946 673174
rect 564182 672938 573866 673174
rect 574102 672938 574186 673174
rect 574422 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 10666 672854
rect 10902 672618 10986 672854
rect 11222 672618 20906 672854
rect 21142 672618 21226 672854
rect 21462 672618 31146 672854
rect 31382 672618 31466 672854
rect 31702 672618 41386 672854
rect 41622 672618 41706 672854
rect 41942 672618 51626 672854
rect 51862 672618 51946 672854
rect 52182 672618 61866 672854
rect 62102 672618 62186 672854
rect 62422 672618 72106 672854
rect 72342 672618 72426 672854
rect 72662 672618 82346 672854
rect 82582 672618 82666 672854
rect 82902 672618 92586 672854
rect 92822 672618 92906 672854
rect 93142 672618 102826 672854
rect 103062 672618 103146 672854
rect 103382 672618 113066 672854
rect 113302 672618 113386 672854
rect 113622 672618 123306 672854
rect 123542 672618 123626 672854
rect 123862 672618 133546 672854
rect 133782 672618 133866 672854
rect 134102 672618 143786 672854
rect 144022 672618 144106 672854
rect 144342 672618 154026 672854
rect 154262 672618 154346 672854
rect 154582 672618 164266 672854
rect 164502 672618 164586 672854
rect 164822 672618 174506 672854
rect 174742 672618 174826 672854
rect 175062 672618 184746 672854
rect 184982 672618 185066 672854
rect 185302 672618 194986 672854
rect 195222 672618 195306 672854
rect 195542 672618 205226 672854
rect 205462 672618 205546 672854
rect 205782 672618 215466 672854
rect 215702 672618 215786 672854
rect 216022 672618 225706 672854
rect 225942 672618 226026 672854
rect 226262 672618 235946 672854
rect 236182 672618 236266 672854
rect 236502 672618 246186 672854
rect 246422 672618 246506 672854
rect 246742 672618 256426 672854
rect 256662 672618 256746 672854
rect 256982 672618 266666 672854
rect 266902 672618 266986 672854
rect 267222 672618 276906 672854
rect 277142 672618 277226 672854
rect 277462 672618 287146 672854
rect 287382 672618 287466 672854
rect 287702 672618 297386 672854
rect 297622 672618 297706 672854
rect 297942 672618 307626 672854
rect 307862 672618 307946 672854
rect 308182 672618 317866 672854
rect 318102 672618 318186 672854
rect 318422 672618 328106 672854
rect 328342 672618 328426 672854
rect 328662 672618 338346 672854
rect 338582 672618 338666 672854
rect 338902 672618 348586 672854
rect 348822 672618 348906 672854
rect 349142 672618 358826 672854
rect 359062 672618 359146 672854
rect 359382 672618 369066 672854
rect 369302 672618 369386 672854
rect 369622 672618 379306 672854
rect 379542 672618 379626 672854
rect 379862 672618 389546 672854
rect 389782 672618 389866 672854
rect 390102 672618 399786 672854
rect 400022 672618 400106 672854
rect 400342 672618 410026 672854
rect 410262 672618 410346 672854
rect 410582 672618 420266 672854
rect 420502 672618 420586 672854
rect 420822 672618 430506 672854
rect 430742 672618 430826 672854
rect 431062 672618 440746 672854
rect 440982 672618 441066 672854
rect 441302 672618 450986 672854
rect 451222 672618 451306 672854
rect 451542 672618 461226 672854
rect 461462 672618 461546 672854
rect 461782 672618 471466 672854
rect 471702 672618 471786 672854
rect 472022 672618 481706 672854
rect 481942 672618 482026 672854
rect 482262 672618 491946 672854
rect 492182 672618 492266 672854
rect 492502 672618 502186 672854
rect 502422 672618 502506 672854
rect 502742 672618 512426 672854
rect 512662 672618 512746 672854
rect 512982 672618 522666 672854
rect 522902 672618 522986 672854
rect 523222 672618 532906 672854
rect 533142 672618 533226 672854
rect 533462 672618 543146 672854
rect 543382 672618 543466 672854
rect 543702 672618 553386 672854
rect 553622 672618 553706 672854
rect 553942 672618 563626 672854
rect 563862 672618 563946 672854
rect 564182 672618 573866 672854
rect 574102 672618 574186 672854
rect 574422 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 6946 669454
rect 7182 669218 7266 669454
rect 7502 669218 17186 669454
rect 17422 669218 17506 669454
rect 17742 669218 27426 669454
rect 27662 669218 27746 669454
rect 27982 669218 37666 669454
rect 37902 669218 37986 669454
rect 38222 669218 47906 669454
rect 48142 669218 48226 669454
rect 48462 669218 58146 669454
rect 58382 669218 58466 669454
rect 58702 669218 68386 669454
rect 68622 669218 68706 669454
rect 68942 669218 78626 669454
rect 78862 669218 78946 669454
rect 79182 669218 88866 669454
rect 89102 669218 89186 669454
rect 89422 669218 99106 669454
rect 99342 669218 99426 669454
rect 99662 669218 109346 669454
rect 109582 669218 109666 669454
rect 109902 669218 119586 669454
rect 119822 669218 119906 669454
rect 120142 669218 129826 669454
rect 130062 669218 130146 669454
rect 130382 669218 140066 669454
rect 140302 669218 140386 669454
rect 140622 669218 150306 669454
rect 150542 669218 150626 669454
rect 150862 669218 160546 669454
rect 160782 669218 160866 669454
rect 161102 669218 170786 669454
rect 171022 669218 171106 669454
rect 171342 669218 181026 669454
rect 181262 669218 181346 669454
rect 181582 669218 191266 669454
rect 191502 669218 191586 669454
rect 191822 669218 201506 669454
rect 201742 669218 201826 669454
rect 202062 669218 211746 669454
rect 211982 669218 212066 669454
rect 212302 669218 221986 669454
rect 222222 669218 222306 669454
rect 222542 669218 232226 669454
rect 232462 669218 232546 669454
rect 232782 669218 242466 669454
rect 242702 669218 242786 669454
rect 243022 669218 252706 669454
rect 252942 669218 253026 669454
rect 253262 669218 262946 669454
rect 263182 669218 263266 669454
rect 263502 669218 273186 669454
rect 273422 669218 273506 669454
rect 273742 669218 283426 669454
rect 283662 669218 283746 669454
rect 283982 669218 293666 669454
rect 293902 669218 293986 669454
rect 294222 669218 303906 669454
rect 304142 669218 304226 669454
rect 304462 669218 314146 669454
rect 314382 669218 314466 669454
rect 314702 669218 324386 669454
rect 324622 669218 324706 669454
rect 324942 669218 334626 669454
rect 334862 669218 334946 669454
rect 335182 669218 344866 669454
rect 345102 669218 345186 669454
rect 345422 669218 355106 669454
rect 355342 669218 355426 669454
rect 355662 669218 365346 669454
rect 365582 669218 365666 669454
rect 365902 669218 375586 669454
rect 375822 669218 375906 669454
rect 376142 669218 385826 669454
rect 386062 669218 386146 669454
rect 386382 669218 396066 669454
rect 396302 669218 396386 669454
rect 396622 669218 406306 669454
rect 406542 669218 406626 669454
rect 406862 669218 416546 669454
rect 416782 669218 416866 669454
rect 417102 669218 426786 669454
rect 427022 669218 427106 669454
rect 427342 669218 437026 669454
rect 437262 669218 437346 669454
rect 437582 669218 447266 669454
rect 447502 669218 447586 669454
rect 447822 669218 457506 669454
rect 457742 669218 457826 669454
rect 458062 669218 467746 669454
rect 467982 669218 468066 669454
rect 468302 669218 477986 669454
rect 478222 669218 478306 669454
rect 478542 669218 488226 669454
rect 488462 669218 488546 669454
rect 488782 669218 498466 669454
rect 498702 669218 498786 669454
rect 499022 669218 508706 669454
rect 508942 669218 509026 669454
rect 509262 669218 518946 669454
rect 519182 669218 519266 669454
rect 519502 669218 529186 669454
rect 529422 669218 529506 669454
rect 529742 669218 539426 669454
rect 539662 669218 539746 669454
rect 539982 669218 549666 669454
rect 549902 669218 549986 669454
rect 550222 669218 559906 669454
rect 560142 669218 560226 669454
rect 560462 669218 570146 669454
rect 570382 669218 570466 669454
rect 570702 669218 580386 669454
rect 580622 669218 580706 669454
rect 580942 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 6946 669134
rect 7182 668898 7266 669134
rect 7502 668898 17186 669134
rect 17422 668898 17506 669134
rect 17742 668898 27426 669134
rect 27662 668898 27746 669134
rect 27982 668898 37666 669134
rect 37902 668898 37986 669134
rect 38222 668898 47906 669134
rect 48142 668898 48226 669134
rect 48462 668898 58146 669134
rect 58382 668898 58466 669134
rect 58702 668898 68386 669134
rect 68622 668898 68706 669134
rect 68942 668898 78626 669134
rect 78862 668898 78946 669134
rect 79182 668898 88866 669134
rect 89102 668898 89186 669134
rect 89422 668898 99106 669134
rect 99342 668898 99426 669134
rect 99662 668898 109346 669134
rect 109582 668898 109666 669134
rect 109902 668898 119586 669134
rect 119822 668898 119906 669134
rect 120142 668898 129826 669134
rect 130062 668898 130146 669134
rect 130382 668898 140066 669134
rect 140302 668898 140386 669134
rect 140622 668898 150306 669134
rect 150542 668898 150626 669134
rect 150862 668898 160546 669134
rect 160782 668898 160866 669134
rect 161102 668898 170786 669134
rect 171022 668898 171106 669134
rect 171342 668898 181026 669134
rect 181262 668898 181346 669134
rect 181582 668898 191266 669134
rect 191502 668898 191586 669134
rect 191822 668898 201506 669134
rect 201742 668898 201826 669134
rect 202062 668898 211746 669134
rect 211982 668898 212066 669134
rect 212302 668898 221986 669134
rect 222222 668898 222306 669134
rect 222542 668898 232226 669134
rect 232462 668898 232546 669134
rect 232782 668898 242466 669134
rect 242702 668898 242786 669134
rect 243022 668898 252706 669134
rect 252942 668898 253026 669134
rect 253262 668898 262946 669134
rect 263182 668898 263266 669134
rect 263502 668898 273186 669134
rect 273422 668898 273506 669134
rect 273742 668898 283426 669134
rect 283662 668898 283746 669134
rect 283982 668898 293666 669134
rect 293902 668898 293986 669134
rect 294222 668898 303906 669134
rect 304142 668898 304226 669134
rect 304462 668898 314146 669134
rect 314382 668898 314466 669134
rect 314702 668898 324386 669134
rect 324622 668898 324706 669134
rect 324942 668898 334626 669134
rect 334862 668898 334946 669134
rect 335182 668898 344866 669134
rect 345102 668898 345186 669134
rect 345422 668898 355106 669134
rect 355342 668898 355426 669134
rect 355662 668898 365346 669134
rect 365582 668898 365666 669134
rect 365902 668898 375586 669134
rect 375822 668898 375906 669134
rect 376142 668898 385826 669134
rect 386062 668898 386146 669134
rect 386382 668898 396066 669134
rect 396302 668898 396386 669134
rect 396622 668898 406306 669134
rect 406542 668898 406626 669134
rect 406862 668898 416546 669134
rect 416782 668898 416866 669134
rect 417102 668898 426786 669134
rect 427022 668898 427106 669134
rect 427342 668898 437026 669134
rect 437262 668898 437346 669134
rect 437582 668898 447266 669134
rect 447502 668898 447586 669134
rect 447822 668898 457506 669134
rect 457742 668898 457826 669134
rect 458062 668898 467746 669134
rect 467982 668898 468066 669134
rect 468302 668898 477986 669134
rect 478222 668898 478306 669134
rect 478542 668898 488226 669134
rect 488462 668898 488546 669134
rect 488782 668898 498466 669134
rect 498702 668898 498786 669134
rect 499022 668898 508706 669134
rect 508942 668898 509026 669134
rect 509262 668898 518946 669134
rect 519182 668898 519266 669134
rect 519502 668898 529186 669134
rect 529422 668898 529506 669134
rect 529742 668898 539426 669134
rect 539662 668898 539746 669134
rect 539982 668898 549666 669134
rect 549902 668898 549986 669134
rect 550222 668898 559906 669134
rect 560142 668898 560226 669134
rect 560462 668898 570146 669134
rect 570382 668898 570466 669134
rect 570702 668898 580386 669134
rect 580622 668898 580706 669134
rect 580942 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 23226 662614
rect 23462 662378 23546 662614
rect 23782 662378 33466 662614
rect 33702 662378 33786 662614
rect 34022 662378 43706 662614
rect 43942 662378 44026 662614
rect 44262 662378 53946 662614
rect 54182 662378 54266 662614
rect 54502 662378 64186 662614
rect 64422 662378 64506 662614
rect 64742 662378 74426 662614
rect 74662 662378 74746 662614
rect 74982 662378 84666 662614
rect 84902 662378 84986 662614
rect 85222 662378 94906 662614
rect 95142 662378 95226 662614
rect 95462 662378 105146 662614
rect 105382 662378 105466 662614
rect 105702 662378 115386 662614
rect 115622 662378 115706 662614
rect 115942 662378 125626 662614
rect 125862 662378 125946 662614
rect 126182 662378 135866 662614
rect 136102 662378 136186 662614
rect 136422 662378 146106 662614
rect 146342 662378 146426 662614
rect 146662 662378 156346 662614
rect 156582 662378 156666 662614
rect 156902 662378 166586 662614
rect 166822 662378 166906 662614
rect 167142 662378 176826 662614
rect 177062 662378 177146 662614
rect 177382 662378 187066 662614
rect 187302 662378 187386 662614
rect 187622 662378 197306 662614
rect 197542 662378 197626 662614
rect 197862 662378 207546 662614
rect 207782 662378 207866 662614
rect 208102 662378 217786 662614
rect 218022 662378 218106 662614
rect 218342 662378 228026 662614
rect 228262 662378 228346 662614
rect 228582 662378 238266 662614
rect 238502 662378 238586 662614
rect 238822 662378 248506 662614
rect 248742 662378 248826 662614
rect 249062 662378 258746 662614
rect 258982 662378 259066 662614
rect 259302 662378 268986 662614
rect 269222 662378 269306 662614
rect 269542 662378 279226 662614
rect 279462 662378 279546 662614
rect 279782 662378 289466 662614
rect 289702 662378 289786 662614
rect 290022 662378 299706 662614
rect 299942 662378 300026 662614
rect 300262 662378 309946 662614
rect 310182 662378 310266 662614
rect 310502 662378 320186 662614
rect 320422 662378 320506 662614
rect 320742 662378 330426 662614
rect 330662 662378 330746 662614
rect 330982 662378 340666 662614
rect 340902 662378 340986 662614
rect 341222 662378 350906 662614
rect 351142 662378 351226 662614
rect 351462 662378 361146 662614
rect 361382 662378 361466 662614
rect 361702 662378 371386 662614
rect 371622 662378 371706 662614
rect 371942 662378 381626 662614
rect 381862 662378 381946 662614
rect 382182 662378 391866 662614
rect 392102 662378 392186 662614
rect 392422 662378 402106 662614
rect 402342 662378 402426 662614
rect 402662 662378 412346 662614
rect 412582 662378 412666 662614
rect 412902 662378 422586 662614
rect 422822 662378 422906 662614
rect 423142 662378 432826 662614
rect 433062 662378 433146 662614
rect 433382 662378 443066 662614
rect 443302 662378 443386 662614
rect 443622 662378 453306 662614
rect 453542 662378 453626 662614
rect 453862 662378 463546 662614
rect 463782 662378 463866 662614
rect 464102 662378 473786 662614
rect 474022 662378 474106 662614
rect 474342 662378 484026 662614
rect 484262 662378 484346 662614
rect 484582 662378 494266 662614
rect 494502 662378 494586 662614
rect 494822 662378 504506 662614
rect 504742 662378 504826 662614
rect 505062 662378 514746 662614
rect 514982 662378 515066 662614
rect 515302 662378 524986 662614
rect 525222 662378 525306 662614
rect 525542 662378 535226 662614
rect 535462 662378 535546 662614
rect 535782 662378 545466 662614
rect 545702 662378 545786 662614
rect 546022 662378 555706 662614
rect 555942 662378 556026 662614
rect 556262 662378 565946 662614
rect 566182 662378 566266 662614
rect 566502 662378 576186 662614
rect 576422 662378 576506 662614
rect 576742 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 23226 662294
rect 23462 662058 23546 662294
rect 23782 662058 33466 662294
rect 33702 662058 33786 662294
rect 34022 662058 43706 662294
rect 43942 662058 44026 662294
rect 44262 662058 53946 662294
rect 54182 662058 54266 662294
rect 54502 662058 64186 662294
rect 64422 662058 64506 662294
rect 64742 662058 74426 662294
rect 74662 662058 74746 662294
rect 74982 662058 84666 662294
rect 84902 662058 84986 662294
rect 85222 662058 94906 662294
rect 95142 662058 95226 662294
rect 95462 662058 105146 662294
rect 105382 662058 105466 662294
rect 105702 662058 115386 662294
rect 115622 662058 115706 662294
rect 115942 662058 125626 662294
rect 125862 662058 125946 662294
rect 126182 662058 135866 662294
rect 136102 662058 136186 662294
rect 136422 662058 146106 662294
rect 146342 662058 146426 662294
rect 146662 662058 156346 662294
rect 156582 662058 156666 662294
rect 156902 662058 166586 662294
rect 166822 662058 166906 662294
rect 167142 662058 176826 662294
rect 177062 662058 177146 662294
rect 177382 662058 187066 662294
rect 187302 662058 187386 662294
rect 187622 662058 197306 662294
rect 197542 662058 197626 662294
rect 197862 662058 207546 662294
rect 207782 662058 207866 662294
rect 208102 662058 217786 662294
rect 218022 662058 218106 662294
rect 218342 662058 228026 662294
rect 228262 662058 228346 662294
rect 228582 662058 238266 662294
rect 238502 662058 238586 662294
rect 238822 662058 248506 662294
rect 248742 662058 248826 662294
rect 249062 662058 258746 662294
rect 258982 662058 259066 662294
rect 259302 662058 268986 662294
rect 269222 662058 269306 662294
rect 269542 662058 279226 662294
rect 279462 662058 279546 662294
rect 279782 662058 289466 662294
rect 289702 662058 289786 662294
rect 290022 662058 299706 662294
rect 299942 662058 300026 662294
rect 300262 662058 309946 662294
rect 310182 662058 310266 662294
rect 310502 662058 320186 662294
rect 320422 662058 320506 662294
rect 320742 662058 330426 662294
rect 330662 662058 330746 662294
rect 330982 662058 340666 662294
rect 340902 662058 340986 662294
rect 341222 662058 350906 662294
rect 351142 662058 351226 662294
rect 351462 662058 361146 662294
rect 361382 662058 361466 662294
rect 361702 662058 371386 662294
rect 371622 662058 371706 662294
rect 371942 662058 381626 662294
rect 381862 662058 381946 662294
rect 382182 662058 391866 662294
rect 392102 662058 392186 662294
rect 392422 662058 402106 662294
rect 402342 662058 402426 662294
rect 402662 662058 412346 662294
rect 412582 662058 412666 662294
rect 412902 662058 422586 662294
rect 422822 662058 422906 662294
rect 423142 662058 432826 662294
rect 433062 662058 433146 662294
rect 433382 662058 443066 662294
rect 443302 662058 443386 662294
rect 443622 662058 453306 662294
rect 453542 662058 453626 662294
rect 453862 662058 463546 662294
rect 463782 662058 463866 662294
rect 464102 662058 473786 662294
rect 474022 662058 474106 662294
rect 474342 662058 484026 662294
rect 484262 662058 484346 662294
rect 484582 662058 494266 662294
rect 494502 662058 494586 662294
rect 494822 662058 504506 662294
rect 504742 662058 504826 662294
rect 505062 662058 514746 662294
rect 514982 662058 515066 662294
rect 515302 662058 524986 662294
rect 525222 662058 525306 662294
rect 525542 662058 535226 662294
rect 535462 662058 535546 662294
rect 535782 662058 545466 662294
rect 545702 662058 545786 662294
rect 546022 662058 555706 662294
rect 555942 662058 556026 662294
rect 556262 662058 565946 662294
rect 566182 662058 566266 662294
rect 566502 662058 576186 662294
rect 576422 662058 576506 662294
rect 576742 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 19506 658894
rect 19742 658658 19826 658894
rect 20062 658658 29746 658894
rect 29982 658658 30066 658894
rect 30302 658658 39986 658894
rect 40222 658658 40306 658894
rect 40542 658658 50226 658894
rect 50462 658658 50546 658894
rect 50782 658658 60466 658894
rect 60702 658658 60786 658894
rect 61022 658658 70706 658894
rect 70942 658658 71026 658894
rect 71262 658658 80946 658894
rect 81182 658658 81266 658894
rect 81502 658658 91186 658894
rect 91422 658658 91506 658894
rect 91742 658658 101426 658894
rect 101662 658658 101746 658894
rect 101982 658658 111666 658894
rect 111902 658658 111986 658894
rect 112222 658658 121906 658894
rect 122142 658658 122226 658894
rect 122462 658658 132146 658894
rect 132382 658658 132466 658894
rect 132702 658658 142386 658894
rect 142622 658658 142706 658894
rect 142942 658658 152626 658894
rect 152862 658658 152946 658894
rect 153182 658658 162866 658894
rect 163102 658658 163186 658894
rect 163422 658658 173106 658894
rect 173342 658658 173426 658894
rect 173662 658658 183346 658894
rect 183582 658658 183666 658894
rect 183902 658658 193586 658894
rect 193822 658658 193906 658894
rect 194142 658658 203826 658894
rect 204062 658658 204146 658894
rect 204382 658658 214066 658894
rect 214302 658658 214386 658894
rect 214622 658658 224306 658894
rect 224542 658658 224626 658894
rect 224862 658658 234546 658894
rect 234782 658658 234866 658894
rect 235102 658658 244786 658894
rect 245022 658658 245106 658894
rect 245342 658658 255026 658894
rect 255262 658658 255346 658894
rect 255582 658658 265266 658894
rect 265502 658658 265586 658894
rect 265822 658658 275506 658894
rect 275742 658658 275826 658894
rect 276062 658658 285746 658894
rect 285982 658658 286066 658894
rect 286302 658658 295986 658894
rect 296222 658658 296306 658894
rect 296542 658658 306226 658894
rect 306462 658658 306546 658894
rect 306782 658658 316466 658894
rect 316702 658658 316786 658894
rect 317022 658658 326706 658894
rect 326942 658658 327026 658894
rect 327262 658658 336946 658894
rect 337182 658658 337266 658894
rect 337502 658658 347186 658894
rect 347422 658658 347506 658894
rect 347742 658658 357426 658894
rect 357662 658658 357746 658894
rect 357982 658658 367666 658894
rect 367902 658658 367986 658894
rect 368222 658658 377906 658894
rect 378142 658658 378226 658894
rect 378462 658658 388146 658894
rect 388382 658658 388466 658894
rect 388702 658658 398386 658894
rect 398622 658658 398706 658894
rect 398942 658658 408626 658894
rect 408862 658658 408946 658894
rect 409182 658658 418866 658894
rect 419102 658658 419186 658894
rect 419422 658658 429106 658894
rect 429342 658658 429426 658894
rect 429662 658658 439346 658894
rect 439582 658658 439666 658894
rect 439902 658658 449586 658894
rect 449822 658658 449906 658894
rect 450142 658658 459826 658894
rect 460062 658658 460146 658894
rect 460382 658658 470066 658894
rect 470302 658658 470386 658894
rect 470622 658658 480306 658894
rect 480542 658658 480626 658894
rect 480862 658658 490546 658894
rect 490782 658658 490866 658894
rect 491102 658658 500786 658894
rect 501022 658658 501106 658894
rect 501342 658658 511026 658894
rect 511262 658658 511346 658894
rect 511582 658658 521266 658894
rect 521502 658658 521586 658894
rect 521822 658658 531506 658894
rect 531742 658658 531826 658894
rect 532062 658658 541746 658894
rect 541982 658658 542066 658894
rect 542302 658658 551986 658894
rect 552222 658658 552306 658894
rect 552542 658658 562226 658894
rect 562462 658658 562546 658894
rect 562782 658658 572466 658894
rect 572702 658658 572786 658894
rect 573022 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 19506 658574
rect 19742 658338 19826 658574
rect 20062 658338 29746 658574
rect 29982 658338 30066 658574
rect 30302 658338 39986 658574
rect 40222 658338 40306 658574
rect 40542 658338 50226 658574
rect 50462 658338 50546 658574
rect 50782 658338 60466 658574
rect 60702 658338 60786 658574
rect 61022 658338 70706 658574
rect 70942 658338 71026 658574
rect 71262 658338 80946 658574
rect 81182 658338 81266 658574
rect 81502 658338 91186 658574
rect 91422 658338 91506 658574
rect 91742 658338 101426 658574
rect 101662 658338 101746 658574
rect 101982 658338 111666 658574
rect 111902 658338 111986 658574
rect 112222 658338 121906 658574
rect 122142 658338 122226 658574
rect 122462 658338 132146 658574
rect 132382 658338 132466 658574
rect 132702 658338 142386 658574
rect 142622 658338 142706 658574
rect 142942 658338 152626 658574
rect 152862 658338 152946 658574
rect 153182 658338 162866 658574
rect 163102 658338 163186 658574
rect 163422 658338 173106 658574
rect 173342 658338 173426 658574
rect 173662 658338 183346 658574
rect 183582 658338 183666 658574
rect 183902 658338 193586 658574
rect 193822 658338 193906 658574
rect 194142 658338 203826 658574
rect 204062 658338 204146 658574
rect 204382 658338 214066 658574
rect 214302 658338 214386 658574
rect 214622 658338 224306 658574
rect 224542 658338 224626 658574
rect 224862 658338 234546 658574
rect 234782 658338 234866 658574
rect 235102 658338 244786 658574
rect 245022 658338 245106 658574
rect 245342 658338 255026 658574
rect 255262 658338 255346 658574
rect 255582 658338 265266 658574
rect 265502 658338 265586 658574
rect 265822 658338 275506 658574
rect 275742 658338 275826 658574
rect 276062 658338 285746 658574
rect 285982 658338 286066 658574
rect 286302 658338 295986 658574
rect 296222 658338 296306 658574
rect 296542 658338 306226 658574
rect 306462 658338 306546 658574
rect 306782 658338 316466 658574
rect 316702 658338 316786 658574
rect 317022 658338 326706 658574
rect 326942 658338 327026 658574
rect 327262 658338 336946 658574
rect 337182 658338 337266 658574
rect 337502 658338 347186 658574
rect 347422 658338 347506 658574
rect 347742 658338 357426 658574
rect 357662 658338 357746 658574
rect 357982 658338 367666 658574
rect 367902 658338 367986 658574
rect 368222 658338 377906 658574
rect 378142 658338 378226 658574
rect 378462 658338 388146 658574
rect 388382 658338 388466 658574
rect 388702 658338 398386 658574
rect 398622 658338 398706 658574
rect 398942 658338 408626 658574
rect 408862 658338 408946 658574
rect 409182 658338 418866 658574
rect 419102 658338 419186 658574
rect 419422 658338 429106 658574
rect 429342 658338 429426 658574
rect 429662 658338 439346 658574
rect 439582 658338 439666 658574
rect 439902 658338 449586 658574
rect 449822 658338 449906 658574
rect 450142 658338 459826 658574
rect 460062 658338 460146 658574
rect 460382 658338 470066 658574
rect 470302 658338 470386 658574
rect 470622 658338 480306 658574
rect 480542 658338 480626 658574
rect 480862 658338 490546 658574
rect 490782 658338 490866 658574
rect 491102 658338 500786 658574
rect 501022 658338 501106 658574
rect 501342 658338 511026 658574
rect 511262 658338 511346 658574
rect 511582 658338 521266 658574
rect 521502 658338 521586 658574
rect 521822 658338 531506 658574
rect 531742 658338 531826 658574
rect 532062 658338 541746 658574
rect 541982 658338 542066 658574
rect 542302 658338 551986 658574
rect 552222 658338 552306 658574
rect 552542 658338 562226 658574
rect 562462 658338 562546 658574
rect 562782 658338 572466 658574
rect 572702 658338 572786 658574
rect 573022 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 15786 655174
rect 16022 654938 16106 655174
rect 16342 654938 548266 655174
rect 548502 654938 548586 655174
rect 548822 654938 558506 655174
rect 558742 654938 558826 655174
rect 559062 654938 568746 655174
rect 568982 654938 569066 655174
rect 569302 654938 578986 655174
rect 579222 654938 579306 655174
rect 579542 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 15786 654854
rect 16022 654618 16106 654854
rect 16342 654618 548266 654854
rect 548502 654618 548586 654854
rect 548822 654618 558506 654854
rect 558742 654618 558826 654854
rect 559062 654618 568746 654854
rect 568982 654618 569066 654854
rect 569302 654618 578986 654854
rect 579222 654618 579306 654854
rect 579542 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 12066 651454
rect 12302 651218 12386 651454
rect 12622 651218 23330 651454
rect 23566 651218 33570 651454
rect 33806 651218 43810 651454
rect 44046 651218 54050 651454
rect 54286 651218 64290 651454
rect 64526 651218 74530 651454
rect 74766 651218 84770 651454
rect 85006 651218 95010 651454
rect 95246 651218 105250 651454
rect 105486 651218 115490 651454
rect 115726 651218 125730 651454
rect 125966 651218 135970 651454
rect 136206 651218 146210 651454
rect 146446 651218 156450 651454
rect 156686 651218 166690 651454
rect 166926 651218 176930 651454
rect 177166 651218 187170 651454
rect 187406 651218 197410 651454
rect 197646 651218 207650 651454
rect 207886 651218 217890 651454
rect 218126 651218 228130 651454
rect 228366 651218 238370 651454
rect 238606 651218 248610 651454
rect 248846 651218 258850 651454
rect 259086 651218 269090 651454
rect 269326 651218 279330 651454
rect 279566 651218 289570 651454
rect 289806 651218 299810 651454
rect 300046 651218 310050 651454
rect 310286 651218 320290 651454
rect 320526 651218 330530 651454
rect 330766 651218 340770 651454
rect 341006 651218 351010 651454
rect 351246 651218 361250 651454
rect 361486 651218 371490 651454
rect 371726 651218 381730 651454
rect 381966 651218 391970 651454
rect 392206 651218 402210 651454
rect 402446 651218 412450 651454
rect 412686 651218 422690 651454
rect 422926 651218 432930 651454
rect 433166 651218 443170 651454
rect 443406 651218 453410 651454
rect 453646 651218 463650 651454
rect 463886 651218 473890 651454
rect 474126 651218 484130 651454
rect 484366 651218 494370 651454
rect 494606 651218 504610 651454
rect 504846 651218 514850 651454
rect 515086 651218 525090 651454
rect 525326 651218 535330 651454
rect 535566 651218 544546 651454
rect 544782 651218 544866 651454
rect 545102 651218 554786 651454
rect 555022 651218 555106 651454
rect 555342 651218 565026 651454
rect 565262 651218 565346 651454
rect 565582 651218 575266 651454
rect 575502 651218 575586 651454
rect 575822 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 12066 651134
rect 12302 650898 12386 651134
rect 12622 650898 23330 651134
rect 23566 650898 33570 651134
rect 33806 650898 43810 651134
rect 44046 650898 54050 651134
rect 54286 650898 64290 651134
rect 64526 650898 74530 651134
rect 74766 650898 84770 651134
rect 85006 650898 95010 651134
rect 95246 650898 105250 651134
rect 105486 650898 115490 651134
rect 115726 650898 125730 651134
rect 125966 650898 135970 651134
rect 136206 650898 146210 651134
rect 146446 650898 156450 651134
rect 156686 650898 166690 651134
rect 166926 650898 176930 651134
rect 177166 650898 187170 651134
rect 187406 650898 197410 651134
rect 197646 650898 207650 651134
rect 207886 650898 217890 651134
rect 218126 650898 228130 651134
rect 228366 650898 238370 651134
rect 238606 650898 248610 651134
rect 248846 650898 258850 651134
rect 259086 650898 269090 651134
rect 269326 650898 279330 651134
rect 279566 650898 289570 651134
rect 289806 650898 299810 651134
rect 300046 650898 310050 651134
rect 310286 650898 320290 651134
rect 320526 650898 330530 651134
rect 330766 650898 340770 651134
rect 341006 650898 351010 651134
rect 351246 650898 361250 651134
rect 361486 650898 371490 651134
rect 371726 650898 381730 651134
rect 381966 650898 391970 651134
rect 392206 650898 402210 651134
rect 402446 650898 412450 651134
rect 412686 650898 422690 651134
rect 422926 650898 432930 651134
rect 433166 650898 443170 651134
rect 443406 650898 453410 651134
rect 453646 650898 463650 651134
rect 463886 650898 473890 651134
rect 474126 650898 484130 651134
rect 484366 650898 494370 651134
rect 494606 650898 504610 651134
rect 504846 650898 514850 651134
rect 515086 650898 525090 651134
rect 525326 650898 535330 651134
rect 535566 650898 544546 651134
rect 544782 650898 544866 651134
rect 545102 650898 554786 651134
rect 555022 650898 555106 651134
rect 555342 650898 565026 651134
rect 565262 650898 565346 651134
rect 565582 650898 575266 651134
rect 575502 650898 575586 651134
rect 575822 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 550586 644614
rect 550822 644378 550906 644614
rect 551142 644378 560826 644614
rect 561062 644378 561146 644614
rect 561382 644378 571066 644614
rect 571302 644378 571386 644614
rect 571622 644378 581306 644614
rect 581542 644378 581626 644614
rect 581862 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 550586 644294
rect 550822 644058 550906 644294
rect 551142 644058 560826 644294
rect 561062 644058 561146 644294
rect 561382 644058 571066 644294
rect 571302 644058 571386 644294
rect 571622 644058 581306 644294
rect 581542 644058 581626 644294
rect 581862 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 14386 640894
rect 14622 640658 14706 640894
rect 14942 640658 546866 640894
rect 547102 640658 547186 640894
rect 547422 640658 557106 640894
rect 557342 640658 557426 640894
rect 557662 640658 567346 640894
rect 567582 640658 567666 640894
rect 567902 640658 577586 640894
rect 577822 640658 577906 640894
rect 578142 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 14386 640574
rect 14622 640338 14706 640574
rect 14942 640338 546866 640574
rect 547102 640338 547186 640574
rect 547422 640338 557106 640574
rect 557342 640338 557426 640574
rect 557662 640338 567346 640574
rect 567582 640338 567666 640574
rect 567902 640338 577586 640574
rect 577822 640338 577906 640574
rect 578142 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 10666 637174
rect 10902 636938 10986 637174
rect 11222 636938 543146 637174
rect 543382 636938 543466 637174
rect 543702 636938 553386 637174
rect 553622 636938 553706 637174
rect 553942 636938 563626 637174
rect 563862 636938 563946 637174
rect 564182 636938 573866 637174
rect 574102 636938 574186 637174
rect 574422 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 10666 636854
rect 10902 636618 10986 636854
rect 11222 636618 543146 636854
rect 543382 636618 543466 636854
rect 543702 636618 553386 636854
rect 553622 636618 553706 636854
rect 553942 636618 563626 636854
rect 563862 636618 563946 636854
rect 564182 636618 573866 636854
rect 574102 636618 574186 636854
rect 574422 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 6946 633454
rect 7182 633218 7266 633454
rect 7502 633218 28450 633454
rect 28686 633218 38690 633454
rect 38926 633218 48930 633454
rect 49166 633218 59170 633454
rect 59406 633218 69410 633454
rect 69646 633218 79650 633454
rect 79886 633218 89890 633454
rect 90126 633218 100130 633454
rect 100366 633218 110370 633454
rect 110606 633218 120610 633454
rect 120846 633218 130850 633454
rect 131086 633218 141090 633454
rect 141326 633218 151330 633454
rect 151566 633218 161570 633454
rect 161806 633218 171810 633454
rect 172046 633218 182050 633454
rect 182286 633218 192290 633454
rect 192526 633218 202530 633454
rect 202766 633218 212770 633454
rect 213006 633218 223010 633454
rect 223246 633218 233250 633454
rect 233486 633218 243490 633454
rect 243726 633218 253730 633454
rect 253966 633218 263970 633454
rect 264206 633218 274210 633454
rect 274446 633218 284450 633454
rect 284686 633218 294690 633454
rect 294926 633218 304930 633454
rect 305166 633218 315170 633454
rect 315406 633218 325410 633454
rect 325646 633218 335650 633454
rect 335886 633218 345890 633454
rect 346126 633218 356130 633454
rect 356366 633218 366370 633454
rect 366606 633218 376610 633454
rect 376846 633218 386850 633454
rect 387086 633218 397090 633454
rect 397326 633218 407330 633454
rect 407566 633218 417570 633454
rect 417806 633218 427810 633454
rect 428046 633218 438050 633454
rect 438286 633218 448290 633454
rect 448526 633218 458530 633454
rect 458766 633218 468770 633454
rect 469006 633218 479010 633454
rect 479246 633218 489250 633454
rect 489486 633218 499490 633454
rect 499726 633218 509730 633454
rect 509966 633218 519970 633454
rect 520206 633218 530210 633454
rect 530446 633218 549666 633454
rect 549902 633218 549986 633454
rect 550222 633218 559906 633454
rect 560142 633218 560226 633454
rect 560462 633218 570146 633454
rect 570382 633218 570466 633454
rect 570702 633218 580386 633454
rect 580622 633218 580706 633454
rect 580942 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 6946 633134
rect 7182 632898 7266 633134
rect 7502 632898 28450 633134
rect 28686 632898 38690 633134
rect 38926 632898 48930 633134
rect 49166 632898 59170 633134
rect 59406 632898 69410 633134
rect 69646 632898 79650 633134
rect 79886 632898 89890 633134
rect 90126 632898 100130 633134
rect 100366 632898 110370 633134
rect 110606 632898 120610 633134
rect 120846 632898 130850 633134
rect 131086 632898 141090 633134
rect 141326 632898 151330 633134
rect 151566 632898 161570 633134
rect 161806 632898 171810 633134
rect 172046 632898 182050 633134
rect 182286 632898 192290 633134
rect 192526 632898 202530 633134
rect 202766 632898 212770 633134
rect 213006 632898 223010 633134
rect 223246 632898 233250 633134
rect 233486 632898 243490 633134
rect 243726 632898 253730 633134
rect 253966 632898 263970 633134
rect 264206 632898 274210 633134
rect 274446 632898 284450 633134
rect 284686 632898 294690 633134
rect 294926 632898 304930 633134
rect 305166 632898 315170 633134
rect 315406 632898 325410 633134
rect 325646 632898 335650 633134
rect 335886 632898 345890 633134
rect 346126 632898 356130 633134
rect 356366 632898 366370 633134
rect 366606 632898 376610 633134
rect 376846 632898 386850 633134
rect 387086 632898 397090 633134
rect 397326 632898 407330 633134
rect 407566 632898 417570 633134
rect 417806 632898 427810 633134
rect 428046 632898 438050 633134
rect 438286 632898 448290 633134
rect 448526 632898 458530 633134
rect 458766 632898 468770 633134
rect 469006 632898 479010 633134
rect 479246 632898 489250 633134
rect 489486 632898 499490 633134
rect 499726 632898 509730 633134
rect 509966 632898 519970 633134
rect 520206 632898 530210 633134
rect 530446 632898 549666 633134
rect 549902 632898 549986 633134
rect 550222 632898 559906 633134
rect 560142 632898 560226 633134
rect 560462 632898 570146 633134
rect 570382 632898 570466 633134
rect 570702 632898 580386 633134
rect 580622 632898 580706 633134
rect 580942 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 545466 626614
rect 545702 626378 545786 626614
rect 546022 626378 555706 626614
rect 555942 626378 556026 626614
rect 556262 626378 565946 626614
rect 566182 626378 566266 626614
rect 566502 626378 576186 626614
rect 576422 626378 576506 626614
rect 576742 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 545466 626294
rect 545702 626058 545786 626294
rect 546022 626058 555706 626294
rect 555942 626058 556026 626294
rect 556262 626058 565946 626294
rect 566182 626058 566266 626294
rect 566502 626058 576186 626294
rect 576422 626058 576506 626294
rect 576742 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 541746 622894
rect 541982 622658 542066 622894
rect 542302 622658 551986 622894
rect 552222 622658 552306 622894
rect 552542 622658 562226 622894
rect 562462 622658 562546 622894
rect 562782 622658 572466 622894
rect 572702 622658 572786 622894
rect 573022 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 541746 622574
rect 541982 622338 542066 622574
rect 542302 622338 551986 622574
rect 552222 622338 552306 622574
rect 552542 622338 562226 622574
rect 562462 622338 562546 622574
rect 562782 622338 572466 622574
rect 572702 622338 572786 622574
rect 573022 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 15786 619174
rect 16022 618938 16106 619174
rect 16342 618938 548266 619174
rect 548502 618938 548586 619174
rect 548822 618938 558506 619174
rect 558742 618938 558826 619174
rect 559062 618938 568746 619174
rect 568982 618938 569066 619174
rect 569302 618938 578986 619174
rect 579222 618938 579306 619174
rect 579542 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 15786 618854
rect 16022 618618 16106 618854
rect 16342 618618 548266 618854
rect 548502 618618 548586 618854
rect 548822 618618 558506 618854
rect 558742 618618 558826 618854
rect 559062 618618 568746 618854
rect 568982 618618 569066 618854
rect 569302 618618 578986 618854
rect 579222 618618 579306 618854
rect 579542 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 12066 615454
rect 12302 615218 12386 615454
rect 12622 615218 23330 615454
rect 23566 615218 33570 615454
rect 33806 615218 43810 615454
rect 44046 615218 54050 615454
rect 54286 615218 64290 615454
rect 64526 615218 74530 615454
rect 74766 615218 84770 615454
rect 85006 615218 95010 615454
rect 95246 615218 105250 615454
rect 105486 615218 115490 615454
rect 115726 615218 125730 615454
rect 125966 615218 135970 615454
rect 136206 615218 146210 615454
rect 146446 615218 156450 615454
rect 156686 615218 166690 615454
rect 166926 615218 176930 615454
rect 177166 615218 187170 615454
rect 187406 615218 197410 615454
rect 197646 615218 207650 615454
rect 207886 615218 217890 615454
rect 218126 615218 228130 615454
rect 228366 615218 238370 615454
rect 238606 615218 248610 615454
rect 248846 615218 258850 615454
rect 259086 615218 269090 615454
rect 269326 615218 279330 615454
rect 279566 615218 289570 615454
rect 289806 615218 299810 615454
rect 300046 615218 310050 615454
rect 310286 615218 320290 615454
rect 320526 615218 330530 615454
rect 330766 615218 340770 615454
rect 341006 615218 351010 615454
rect 351246 615218 361250 615454
rect 361486 615218 371490 615454
rect 371726 615218 381730 615454
rect 381966 615218 391970 615454
rect 392206 615218 402210 615454
rect 402446 615218 412450 615454
rect 412686 615218 422690 615454
rect 422926 615218 432930 615454
rect 433166 615218 443170 615454
rect 443406 615218 453410 615454
rect 453646 615218 463650 615454
rect 463886 615218 473890 615454
rect 474126 615218 484130 615454
rect 484366 615218 494370 615454
rect 494606 615218 504610 615454
rect 504846 615218 514850 615454
rect 515086 615218 525090 615454
rect 525326 615218 535330 615454
rect 535566 615218 544546 615454
rect 544782 615218 544866 615454
rect 545102 615218 554786 615454
rect 555022 615218 555106 615454
rect 555342 615218 565026 615454
rect 565262 615218 565346 615454
rect 565582 615218 575266 615454
rect 575502 615218 575586 615454
rect 575822 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 12066 615134
rect 12302 614898 12386 615134
rect 12622 614898 23330 615134
rect 23566 614898 33570 615134
rect 33806 614898 43810 615134
rect 44046 614898 54050 615134
rect 54286 614898 64290 615134
rect 64526 614898 74530 615134
rect 74766 614898 84770 615134
rect 85006 614898 95010 615134
rect 95246 614898 105250 615134
rect 105486 614898 115490 615134
rect 115726 614898 125730 615134
rect 125966 614898 135970 615134
rect 136206 614898 146210 615134
rect 146446 614898 156450 615134
rect 156686 614898 166690 615134
rect 166926 614898 176930 615134
rect 177166 614898 187170 615134
rect 187406 614898 197410 615134
rect 197646 614898 207650 615134
rect 207886 614898 217890 615134
rect 218126 614898 228130 615134
rect 228366 614898 238370 615134
rect 238606 614898 248610 615134
rect 248846 614898 258850 615134
rect 259086 614898 269090 615134
rect 269326 614898 279330 615134
rect 279566 614898 289570 615134
rect 289806 614898 299810 615134
rect 300046 614898 310050 615134
rect 310286 614898 320290 615134
rect 320526 614898 330530 615134
rect 330766 614898 340770 615134
rect 341006 614898 351010 615134
rect 351246 614898 361250 615134
rect 361486 614898 371490 615134
rect 371726 614898 381730 615134
rect 381966 614898 391970 615134
rect 392206 614898 402210 615134
rect 402446 614898 412450 615134
rect 412686 614898 422690 615134
rect 422926 614898 432930 615134
rect 433166 614898 443170 615134
rect 443406 614898 453410 615134
rect 453646 614898 463650 615134
rect 463886 614898 473890 615134
rect 474126 614898 484130 615134
rect 484366 614898 494370 615134
rect 494606 614898 504610 615134
rect 504846 614898 514850 615134
rect 515086 614898 525090 615134
rect 525326 614898 535330 615134
rect 535566 614898 544546 615134
rect 544782 614898 544866 615134
rect 545102 614898 554786 615134
rect 555022 614898 555106 615134
rect 555342 614898 565026 615134
rect 565262 614898 565346 615134
rect 565582 614898 575266 615134
rect 575502 614898 575586 615134
rect 575822 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 550586 608614
rect 550822 608378 550906 608614
rect 551142 608378 560826 608614
rect 561062 608378 561146 608614
rect 561382 608378 571066 608614
rect 571302 608378 571386 608614
rect 571622 608378 581306 608614
rect 581542 608378 581626 608614
rect 581862 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 550586 608294
rect 550822 608058 550906 608294
rect 551142 608058 560826 608294
rect 561062 608058 561146 608294
rect 561382 608058 571066 608294
rect 571302 608058 571386 608294
rect 571622 608058 581306 608294
rect 581542 608058 581626 608294
rect 581862 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 14386 604894
rect 14622 604658 14706 604894
rect 14942 604658 546866 604894
rect 547102 604658 547186 604894
rect 547422 604658 557106 604894
rect 557342 604658 557426 604894
rect 557662 604658 567346 604894
rect 567582 604658 567666 604894
rect 567902 604658 577586 604894
rect 577822 604658 577906 604894
rect 578142 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 14386 604574
rect 14622 604338 14706 604574
rect 14942 604338 546866 604574
rect 547102 604338 547186 604574
rect 547422 604338 557106 604574
rect 557342 604338 557426 604574
rect 557662 604338 567346 604574
rect 567582 604338 567666 604574
rect 567902 604338 577586 604574
rect 577822 604338 577906 604574
rect 578142 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 10666 601174
rect 10902 600938 10986 601174
rect 11222 600938 543146 601174
rect 543382 600938 543466 601174
rect 543702 600938 553386 601174
rect 553622 600938 553706 601174
rect 553942 600938 563626 601174
rect 563862 600938 563946 601174
rect 564182 600938 573866 601174
rect 574102 600938 574186 601174
rect 574422 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 10666 600854
rect 10902 600618 10986 600854
rect 11222 600618 543146 600854
rect 543382 600618 543466 600854
rect 543702 600618 553386 600854
rect 553622 600618 553706 600854
rect 553942 600618 563626 600854
rect 563862 600618 563946 600854
rect 564182 600618 573866 600854
rect 574102 600618 574186 600854
rect 574422 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 6946 597454
rect 7182 597218 7266 597454
rect 7502 597218 28450 597454
rect 28686 597218 38690 597454
rect 38926 597218 48930 597454
rect 49166 597218 59170 597454
rect 59406 597218 69410 597454
rect 69646 597218 79650 597454
rect 79886 597218 89890 597454
rect 90126 597218 100130 597454
rect 100366 597218 110370 597454
rect 110606 597218 120610 597454
rect 120846 597218 130850 597454
rect 131086 597218 141090 597454
rect 141326 597218 151330 597454
rect 151566 597218 161570 597454
rect 161806 597218 171810 597454
rect 172046 597218 182050 597454
rect 182286 597218 192290 597454
rect 192526 597218 202530 597454
rect 202766 597218 212770 597454
rect 213006 597218 223010 597454
rect 223246 597218 233250 597454
rect 233486 597218 243490 597454
rect 243726 597218 253730 597454
rect 253966 597218 263970 597454
rect 264206 597218 274210 597454
rect 274446 597218 284450 597454
rect 284686 597218 294690 597454
rect 294926 597218 304930 597454
rect 305166 597218 315170 597454
rect 315406 597218 325410 597454
rect 325646 597218 335650 597454
rect 335886 597218 345890 597454
rect 346126 597218 356130 597454
rect 356366 597218 366370 597454
rect 366606 597218 376610 597454
rect 376846 597218 386850 597454
rect 387086 597218 397090 597454
rect 397326 597218 407330 597454
rect 407566 597218 417570 597454
rect 417806 597218 427810 597454
rect 428046 597218 438050 597454
rect 438286 597218 448290 597454
rect 448526 597218 458530 597454
rect 458766 597218 468770 597454
rect 469006 597218 479010 597454
rect 479246 597218 489250 597454
rect 489486 597218 499490 597454
rect 499726 597218 509730 597454
rect 509966 597218 519970 597454
rect 520206 597218 530210 597454
rect 530446 597218 549666 597454
rect 549902 597218 549986 597454
rect 550222 597218 559906 597454
rect 560142 597218 560226 597454
rect 560462 597218 570146 597454
rect 570382 597218 570466 597454
rect 570702 597218 580386 597454
rect 580622 597218 580706 597454
rect 580942 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 6946 597134
rect 7182 596898 7266 597134
rect 7502 596898 28450 597134
rect 28686 596898 38690 597134
rect 38926 596898 48930 597134
rect 49166 596898 59170 597134
rect 59406 596898 69410 597134
rect 69646 596898 79650 597134
rect 79886 596898 89890 597134
rect 90126 596898 100130 597134
rect 100366 596898 110370 597134
rect 110606 596898 120610 597134
rect 120846 596898 130850 597134
rect 131086 596898 141090 597134
rect 141326 596898 151330 597134
rect 151566 596898 161570 597134
rect 161806 596898 171810 597134
rect 172046 596898 182050 597134
rect 182286 596898 192290 597134
rect 192526 596898 202530 597134
rect 202766 596898 212770 597134
rect 213006 596898 223010 597134
rect 223246 596898 233250 597134
rect 233486 596898 243490 597134
rect 243726 596898 253730 597134
rect 253966 596898 263970 597134
rect 264206 596898 274210 597134
rect 274446 596898 284450 597134
rect 284686 596898 294690 597134
rect 294926 596898 304930 597134
rect 305166 596898 315170 597134
rect 315406 596898 325410 597134
rect 325646 596898 335650 597134
rect 335886 596898 345890 597134
rect 346126 596898 356130 597134
rect 356366 596898 366370 597134
rect 366606 596898 376610 597134
rect 376846 596898 386850 597134
rect 387086 596898 397090 597134
rect 397326 596898 407330 597134
rect 407566 596898 417570 597134
rect 417806 596898 427810 597134
rect 428046 596898 438050 597134
rect 438286 596898 448290 597134
rect 448526 596898 458530 597134
rect 458766 596898 468770 597134
rect 469006 596898 479010 597134
rect 479246 596898 489250 597134
rect 489486 596898 499490 597134
rect 499726 596898 509730 597134
rect 509966 596898 519970 597134
rect 520206 596898 530210 597134
rect 530446 596898 549666 597134
rect 549902 596898 549986 597134
rect 550222 596898 559906 597134
rect 560142 596898 560226 597134
rect 560462 596898 570146 597134
rect 570382 596898 570466 597134
rect 570702 596898 580386 597134
rect 580622 596898 580706 597134
rect 580942 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 545466 590614
rect 545702 590378 545786 590614
rect 546022 590378 555706 590614
rect 555942 590378 556026 590614
rect 556262 590378 565946 590614
rect 566182 590378 566266 590614
rect 566502 590378 576186 590614
rect 576422 590378 576506 590614
rect 576742 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 545466 590294
rect 545702 590058 545786 590294
rect 546022 590058 555706 590294
rect 555942 590058 556026 590294
rect 556262 590058 565946 590294
rect 566182 590058 566266 590294
rect 566502 590058 576186 590294
rect 576422 590058 576506 590294
rect 576742 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 541746 586894
rect 541982 586658 542066 586894
rect 542302 586658 551986 586894
rect 552222 586658 552306 586894
rect 552542 586658 562226 586894
rect 562462 586658 562546 586894
rect 562782 586658 572466 586894
rect 572702 586658 572786 586894
rect 573022 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 541746 586574
rect 541982 586338 542066 586574
rect 542302 586338 551986 586574
rect 552222 586338 552306 586574
rect 552542 586338 562226 586574
rect 562462 586338 562546 586574
rect 562782 586338 572466 586574
rect 572702 586338 572786 586574
rect 573022 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 15786 583174
rect 16022 582938 16106 583174
rect 16342 582938 548266 583174
rect 548502 582938 548586 583174
rect 548822 582938 558506 583174
rect 558742 582938 558826 583174
rect 559062 582938 568746 583174
rect 568982 582938 569066 583174
rect 569302 582938 578986 583174
rect 579222 582938 579306 583174
rect 579542 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 15786 582854
rect 16022 582618 16106 582854
rect 16342 582618 548266 582854
rect 548502 582618 548586 582854
rect 548822 582618 558506 582854
rect 558742 582618 558826 582854
rect 559062 582618 568746 582854
rect 568982 582618 569066 582854
rect 569302 582618 578986 582854
rect 579222 582618 579306 582854
rect 579542 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 12066 579454
rect 12302 579218 12386 579454
rect 12622 579218 23330 579454
rect 23566 579218 33570 579454
rect 33806 579218 43810 579454
rect 44046 579218 54050 579454
rect 54286 579218 64290 579454
rect 64526 579218 74530 579454
rect 74766 579218 84770 579454
rect 85006 579218 95010 579454
rect 95246 579218 105250 579454
rect 105486 579218 115490 579454
rect 115726 579218 125730 579454
rect 125966 579218 135970 579454
rect 136206 579218 146210 579454
rect 146446 579218 156450 579454
rect 156686 579218 166690 579454
rect 166926 579218 176930 579454
rect 177166 579218 187170 579454
rect 187406 579218 197410 579454
rect 197646 579218 207650 579454
rect 207886 579218 217890 579454
rect 218126 579218 228130 579454
rect 228366 579218 238370 579454
rect 238606 579218 248610 579454
rect 248846 579218 258850 579454
rect 259086 579218 269090 579454
rect 269326 579218 279330 579454
rect 279566 579218 289570 579454
rect 289806 579218 299810 579454
rect 300046 579218 310050 579454
rect 310286 579218 320290 579454
rect 320526 579218 330530 579454
rect 330766 579218 340770 579454
rect 341006 579218 351010 579454
rect 351246 579218 361250 579454
rect 361486 579218 371490 579454
rect 371726 579218 381730 579454
rect 381966 579218 391970 579454
rect 392206 579218 402210 579454
rect 402446 579218 412450 579454
rect 412686 579218 422690 579454
rect 422926 579218 432930 579454
rect 433166 579218 443170 579454
rect 443406 579218 453410 579454
rect 453646 579218 463650 579454
rect 463886 579218 473890 579454
rect 474126 579218 484130 579454
rect 484366 579218 494370 579454
rect 494606 579218 504610 579454
rect 504846 579218 514850 579454
rect 515086 579218 525090 579454
rect 525326 579218 535330 579454
rect 535566 579218 544546 579454
rect 544782 579218 544866 579454
rect 545102 579218 554786 579454
rect 555022 579218 555106 579454
rect 555342 579218 565026 579454
rect 565262 579218 565346 579454
rect 565582 579218 575266 579454
rect 575502 579218 575586 579454
rect 575822 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 12066 579134
rect 12302 578898 12386 579134
rect 12622 578898 23330 579134
rect 23566 578898 33570 579134
rect 33806 578898 43810 579134
rect 44046 578898 54050 579134
rect 54286 578898 64290 579134
rect 64526 578898 74530 579134
rect 74766 578898 84770 579134
rect 85006 578898 95010 579134
rect 95246 578898 105250 579134
rect 105486 578898 115490 579134
rect 115726 578898 125730 579134
rect 125966 578898 135970 579134
rect 136206 578898 146210 579134
rect 146446 578898 156450 579134
rect 156686 578898 166690 579134
rect 166926 578898 176930 579134
rect 177166 578898 187170 579134
rect 187406 578898 197410 579134
rect 197646 578898 207650 579134
rect 207886 578898 217890 579134
rect 218126 578898 228130 579134
rect 228366 578898 238370 579134
rect 238606 578898 248610 579134
rect 248846 578898 258850 579134
rect 259086 578898 269090 579134
rect 269326 578898 279330 579134
rect 279566 578898 289570 579134
rect 289806 578898 299810 579134
rect 300046 578898 310050 579134
rect 310286 578898 320290 579134
rect 320526 578898 330530 579134
rect 330766 578898 340770 579134
rect 341006 578898 351010 579134
rect 351246 578898 361250 579134
rect 361486 578898 371490 579134
rect 371726 578898 381730 579134
rect 381966 578898 391970 579134
rect 392206 578898 402210 579134
rect 402446 578898 412450 579134
rect 412686 578898 422690 579134
rect 422926 578898 432930 579134
rect 433166 578898 443170 579134
rect 443406 578898 453410 579134
rect 453646 578898 463650 579134
rect 463886 578898 473890 579134
rect 474126 578898 484130 579134
rect 484366 578898 494370 579134
rect 494606 578898 504610 579134
rect 504846 578898 514850 579134
rect 515086 578898 525090 579134
rect 525326 578898 535330 579134
rect 535566 578898 544546 579134
rect 544782 578898 544866 579134
rect 545102 578898 554786 579134
rect 555022 578898 555106 579134
rect 555342 578898 565026 579134
rect 565262 578898 565346 579134
rect 565582 578898 575266 579134
rect 575502 578898 575586 579134
rect 575822 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 550586 572614
rect 550822 572378 550906 572614
rect 551142 572378 560826 572614
rect 561062 572378 561146 572614
rect 561382 572378 571066 572614
rect 571302 572378 571386 572614
rect 571622 572378 581306 572614
rect 581542 572378 581626 572614
rect 581862 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 550586 572294
rect 550822 572058 550906 572294
rect 551142 572058 560826 572294
rect 561062 572058 561146 572294
rect 561382 572058 571066 572294
rect 571302 572058 571386 572294
rect 571622 572058 581306 572294
rect 581542 572058 581626 572294
rect 581862 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 14386 568894
rect 14622 568658 14706 568894
rect 14942 568658 546866 568894
rect 547102 568658 547186 568894
rect 547422 568658 557106 568894
rect 557342 568658 557426 568894
rect 557662 568658 567346 568894
rect 567582 568658 567666 568894
rect 567902 568658 577586 568894
rect 577822 568658 577906 568894
rect 578142 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 14386 568574
rect 14622 568338 14706 568574
rect 14942 568338 546866 568574
rect 547102 568338 547186 568574
rect 547422 568338 557106 568574
rect 557342 568338 557426 568574
rect 557662 568338 567346 568574
rect 567582 568338 567666 568574
rect 567902 568338 577586 568574
rect 577822 568338 577906 568574
rect 578142 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 10666 565174
rect 10902 564938 10986 565174
rect 11222 564938 543146 565174
rect 543382 564938 543466 565174
rect 543702 564938 553386 565174
rect 553622 564938 553706 565174
rect 553942 564938 563626 565174
rect 563862 564938 563946 565174
rect 564182 564938 573866 565174
rect 574102 564938 574186 565174
rect 574422 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 10666 564854
rect 10902 564618 10986 564854
rect 11222 564618 543146 564854
rect 543382 564618 543466 564854
rect 543702 564618 553386 564854
rect 553622 564618 553706 564854
rect 553942 564618 563626 564854
rect 563862 564618 563946 564854
rect 564182 564618 573866 564854
rect 574102 564618 574186 564854
rect 574422 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 6946 561454
rect 7182 561218 7266 561454
rect 7502 561218 28450 561454
rect 28686 561218 38690 561454
rect 38926 561218 48930 561454
rect 49166 561218 59170 561454
rect 59406 561218 69410 561454
rect 69646 561218 79650 561454
rect 79886 561218 89890 561454
rect 90126 561218 100130 561454
rect 100366 561218 110370 561454
rect 110606 561218 120610 561454
rect 120846 561218 130850 561454
rect 131086 561218 141090 561454
rect 141326 561218 151330 561454
rect 151566 561218 161570 561454
rect 161806 561218 171810 561454
rect 172046 561218 182050 561454
rect 182286 561218 192290 561454
rect 192526 561218 202530 561454
rect 202766 561218 212770 561454
rect 213006 561218 223010 561454
rect 223246 561218 233250 561454
rect 233486 561218 243490 561454
rect 243726 561218 253730 561454
rect 253966 561218 263970 561454
rect 264206 561218 274210 561454
rect 274446 561218 284450 561454
rect 284686 561218 294690 561454
rect 294926 561218 304930 561454
rect 305166 561218 315170 561454
rect 315406 561218 325410 561454
rect 325646 561218 335650 561454
rect 335886 561218 345890 561454
rect 346126 561218 356130 561454
rect 356366 561218 366370 561454
rect 366606 561218 376610 561454
rect 376846 561218 386850 561454
rect 387086 561218 397090 561454
rect 397326 561218 407330 561454
rect 407566 561218 417570 561454
rect 417806 561218 427810 561454
rect 428046 561218 438050 561454
rect 438286 561218 448290 561454
rect 448526 561218 458530 561454
rect 458766 561218 468770 561454
rect 469006 561218 479010 561454
rect 479246 561218 489250 561454
rect 489486 561218 499490 561454
rect 499726 561218 509730 561454
rect 509966 561218 519970 561454
rect 520206 561218 530210 561454
rect 530446 561218 549666 561454
rect 549902 561218 549986 561454
rect 550222 561218 559906 561454
rect 560142 561218 560226 561454
rect 560462 561218 570146 561454
rect 570382 561218 570466 561454
rect 570702 561218 580386 561454
rect 580622 561218 580706 561454
rect 580942 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 6946 561134
rect 7182 560898 7266 561134
rect 7502 560898 28450 561134
rect 28686 560898 38690 561134
rect 38926 560898 48930 561134
rect 49166 560898 59170 561134
rect 59406 560898 69410 561134
rect 69646 560898 79650 561134
rect 79886 560898 89890 561134
rect 90126 560898 100130 561134
rect 100366 560898 110370 561134
rect 110606 560898 120610 561134
rect 120846 560898 130850 561134
rect 131086 560898 141090 561134
rect 141326 560898 151330 561134
rect 151566 560898 161570 561134
rect 161806 560898 171810 561134
rect 172046 560898 182050 561134
rect 182286 560898 192290 561134
rect 192526 560898 202530 561134
rect 202766 560898 212770 561134
rect 213006 560898 223010 561134
rect 223246 560898 233250 561134
rect 233486 560898 243490 561134
rect 243726 560898 253730 561134
rect 253966 560898 263970 561134
rect 264206 560898 274210 561134
rect 274446 560898 284450 561134
rect 284686 560898 294690 561134
rect 294926 560898 304930 561134
rect 305166 560898 315170 561134
rect 315406 560898 325410 561134
rect 325646 560898 335650 561134
rect 335886 560898 345890 561134
rect 346126 560898 356130 561134
rect 356366 560898 366370 561134
rect 366606 560898 376610 561134
rect 376846 560898 386850 561134
rect 387086 560898 397090 561134
rect 397326 560898 407330 561134
rect 407566 560898 417570 561134
rect 417806 560898 427810 561134
rect 428046 560898 438050 561134
rect 438286 560898 448290 561134
rect 448526 560898 458530 561134
rect 458766 560898 468770 561134
rect 469006 560898 479010 561134
rect 479246 560898 489250 561134
rect 489486 560898 499490 561134
rect 499726 560898 509730 561134
rect 509966 560898 519970 561134
rect 520206 560898 530210 561134
rect 530446 560898 549666 561134
rect 549902 560898 549986 561134
rect 550222 560898 559906 561134
rect 560142 560898 560226 561134
rect 560462 560898 570146 561134
rect 570382 560898 570466 561134
rect 570702 560898 580386 561134
rect 580622 560898 580706 561134
rect 580942 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 545466 554614
rect 545702 554378 545786 554614
rect 546022 554378 555706 554614
rect 555942 554378 556026 554614
rect 556262 554378 565946 554614
rect 566182 554378 566266 554614
rect 566502 554378 576186 554614
rect 576422 554378 576506 554614
rect 576742 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 545466 554294
rect 545702 554058 545786 554294
rect 546022 554058 555706 554294
rect 555942 554058 556026 554294
rect 556262 554058 565946 554294
rect 566182 554058 566266 554294
rect 566502 554058 576186 554294
rect 576422 554058 576506 554294
rect 576742 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 541746 550894
rect 541982 550658 542066 550894
rect 542302 550658 551986 550894
rect 552222 550658 552306 550894
rect 552542 550658 562226 550894
rect 562462 550658 562546 550894
rect 562782 550658 572466 550894
rect 572702 550658 572786 550894
rect 573022 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 541746 550574
rect 541982 550338 542066 550574
rect 542302 550338 551986 550574
rect 552222 550338 552306 550574
rect 552542 550338 562226 550574
rect 562462 550338 562546 550574
rect 562782 550338 572466 550574
rect 572702 550338 572786 550574
rect 573022 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 15786 547174
rect 16022 546938 16106 547174
rect 16342 546938 548266 547174
rect 548502 546938 548586 547174
rect 548822 546938 558506 547174
rect 558742 546938 558826 547174
rect 559062 546938 568746 547174
rect 568982 546938 569066 547174
rect 569302 546938 578986 547174
rect 579222 546938 579306 547174
rect 579542 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 15786 546854
rect 16022 546618 16106 546854
rect 16342 546618 548266 546854
rect 548502 546618 548586 546854
rect 548822 546618 558506 546854
rect 558742 546618 558826 546854
rect 559062 546618 568746 546854
rect 568982 546618 569066 546854
rect 569302 546618 578986 546854
rect 579222 546618 579306 546854
rect 579542 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 12066 543454
rect 12302 543218 12386 543454
rect 12622 543218 23330 543454
rect 23566 543218 33570 543454
rect 33806 543218 43810 543454
rect 44046 543218 54050 543454
rect 54286 543218 64290 543454
rect 64526 543218 74530 543454
rect 74766 543218 84770 543454
rect 85006 543218 95010 543454
rect 95246 543218 105250 543454
rect 105486 543218 115490 543454
rect 115726 543218 125730 543454
rect 125966 543218 135970 543454
rect 136206 543218 146210 543454
rect 146446 543218 156450 543454
rect 156686 543218 166690 543454
rect 166926 543218 176930 543454
rect 177166 543218 187170 543454
rect 187406 543218 197410 543454
rect 197646 543218 207650 543454
rect 207886 543218 217890 543454
rect 218126 543218 228130 543454
rect 228366 543218 238370 543454
rect 238606 543218 248610 543454
rect 248846 543218 258850 543454
rect 259086 543218 269090 543454
rect 269326 543218 279330 543454
rect 279566 543218 289570 543454
rect 289806 543218 299810 543454
rect 300046 543218 310050 543454
rect 310286 543218 320290 543454
rect 320526 543218 330530 543454
rect 330766 543218 340770 543454
rect 341006 543218 351010 543454
rect 351246 543218 361250 543454
rect 361486 543218 371490 543454
rect 371726 543218 381730 543454
rect 381966 543218 391970 543454
rect 392206 543218 402210 543454
rect 402446 543218 412450 543454
rect 412686 543218 422690 543454
rect 422926 543218 432930 543454
rect 433166 543218 443170 543454
rect 443406 543218 453410 543454
rect 453646 543218 463650 543454
rect 463886 543218 473890 543454
rect 474126 543218 484130 543454
rect 484366 543218 494370 543454
rect 494606 543218 504610 543454
rect 504846 543218 514850 543454
rect 515086 543218 525090 543454
rect 525326 543218 535330 543454
rect 535566 543218 544546 543454
rect 544782 543218 544866 543454
rect 545102 543218 554786 543454
rect 555022 543218 555106 543454
rect 555342 543218 565026 543454
rect 565262 543218 565346 543454
rect 565582 543218 575266 543454
rect 575502 543218 575586 543454
rect 575822 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 12066 543134
rect 12302 542898 12386 543134
rect 12622 542898 23330 543134
rect 23566 542898 33570 543134
rect 33806 542898 43810 543134
rect 44046 542898 54050 543134
rect 54286 542898 64290 543134
rect 64526 542898 74530 543134
rect 74766 542898 84770 543134
rect 85006 542898 95010 543134
rect 95246 542898 105250 543134
rect 105486 542898 115490 543134
rect 115726 542898 125730 543134
rect 125966 542898 135970 543134
rect 136206 542898 146210 543134
rect 146446 542898 156450 543134
rect 156686 542898 166690 543134
rect 166926 542898 176930 543134
rect 177166 542898 187170 543134
rect 187406 542898 197410 543134
rect 197646 542898 207650 543134
rect 207886 542898 217890 543134
rect 218126 542898 228130 543134
rect 228366 542898 238370 543134
rect 238606 542898 248610 543134
rect 248846 542898 258850 543134
rect 259086 542898 269090 543134
rect 269326 542898 279330 543134
rect 279566 542898 289570 543134
rect 289806 542898 299810 543134
rect 300046 542898 310050 543134
rect 310286 542898 320290 543134
rect 320526 542898 330530 543134
rect 330766 542898 340770 543134
rect 341006 542898 351010 543134
rect 351246 542898 361250 543134
rect 361486 542898 371490 543134
rect 371726 542898 381730 543134
rect 381966 542898 391970 543134
rect 392206 542898 402210 543134
rect 402446 542898 412450 543134
rect 412686 542898 422690 543134
rect 422926 542898 432930 543134
rect 433166 542898 443170 543134
rect 443406 542898 453410 543134
rect 453646 542898 463650 543134
rect 463886 542898 473890 543134
rect 474126 542898 484130 543134
rect 484366 542898 494370 543134
rect 494606 542898 504610 543134
rect 504846 542898 514850 543134
rect 515086 542898 525090 543134
rect 525326 542898 535330 543134
rect 535566 542898 544546 543134
rect 544782 542898 544866 543134
rect 545102 542898 554786 543134
rect 555022 542898 555106 543134
rect 555342 542898 565026 543134
rect 565262 542898 565346 543134
rect 565582 542898 575266 543134
rect 575502 542898 575586 543134
rect 575822 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 550586 536614
rect 550822 536378 550906 536614
rect 551142 536378 560826 536614
rect 561062 536378 561146 536614
rect 561382 536378 571066 536614
rect 571302 536378 571386 536614
rect 571622 536378 581306 536614
rect 581542 536378 581626 536614
rect 581862 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 550586 536294
rect 550822 536058 550906 536294
rect 551142 536058 560826 536294
rect 561062 536058 561146 536294
rect 561382 536058 571066 536294
rect 571302 536058 571386 536294
rect 571622 536058 581306 536294
rect 581542 536058 581626 536294
rect 581862 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 14386 532894
rect 14622 532658 14706 532894
rect 14942 532658 546866 532894
rect 547102 532658 547186 532894
rect 547422 532658 557106 532894
rect 557342 532658 557426 532894
rect 557662 532658 567346 532894
rect 567582 532658 567666 532894
rect 567902 532658 577586 532894
rect 577822 532658 577906 532894
rect 578142 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 14386 532574
rect 14622 532338 14706 532574
rect 14942 532338 546866 532574
rect 547102 532338 547186 532574
rect 547422 532338 557106 532574
rect 557342 532338 557426 532574
rect 557662 532338 567346 532574
rect 567582 532338 567666 532574
rect 567902 532338 577586 532574
rect 577822 532338 577906 532574
rect 578142 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 10666 529174
rect 10902 528938 10986 529174
rect 11222 528938 543146 529174
rect 543382 528938 543466 529174
rect 543702 528938 553386 529174
rect 553622 528938 553706 529174
rect 553942 528938 563626 529174
rect 563862 528938 563946 529174
rect 564182 528938 573866 529174
rect 574102 528938 574186 529174
rect 574422 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 10666 528854
rect 10902 528618 10986 528854
rect 11222 528618 543146 528854
rect 543382 528618 543466 528854
rect 543702 528618 553386 528854
rect 553622 528618 553706 528854
rect 553942 528618 563626 528854
rect 563862 528618 563946 528854
rect 564182 528618 573866 528854
rect 574102 528618 574186 528854
rect 574422 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 6946 525454
rect 7182 525218 7266 525454
rect 7502 525218 28450 525454
rect 28686 525218 38690 525454
rect 38926 525218 48930 525454
rect 49166 525218 59170 525454
rect 59406 525218 69410 525454
rect 69646 525218 79650 525454
rect 79886 525218 89890 525454
rect 90126 525218 100130 525454
rect 100366 525218 110370 525454
rect 110606 525218 120610 525454
rect 120846 525218 130850 525454
rect 131086 525218 141090 525454
rect 141326 525218 151330 525454
rect 151566 525218 161570 525454
rect 161806 525218 171810 525454
rect 172046 525218 182050 525454
rect 182286 525218 192290 525454
rect 192526 525218 202530 525454
rect 202766 525218 212770 525454
rect 213006 525218 223010 525454
rect 223246 525218 233250 525454
rect 233486 525218 243490 525454
rect 243726 525218 253730 525454
rect 253966 525218 263970 525454
rect 264206 525218 274210 525454
rect 274446 525218 284450 525454
rect 284686 525218 294690 525454
rect 294926 525218 304930 525454
rect 305166 525218 315170 525454
rect 315406 525218 325410 525454
rect 325646 525218 335650 525454
rect 335886 525218 345890 525454
rect 346126 525218 356130 525454
rect 356366 525218 366370 525454
rect 366606 525218 376610 525454
rect 376846 525218 386850 525454
rect 387086 525218 397090 525454
rect 397326 525218 407330 525454
rect 407566 525218 417570 525454
rect 417806 525218 427810 525454
rect 428046 525218 438050 525454
rect 438286 525218 448290 525454
rect 448526 525218 458530 525454
rect 458766 525218 468770 525454
rect 469006 525218 479010 525454
rect 479246 525218 489250 525454
rect 489486 525218 499490 525454
rect 499726 525218 509730 525454
rect 509966 525218 519970 525454
rect 520206 525218 530210 525454
rect 530446 525218 549666 525454
rect 549902 525218 549986 525454
rect 550222 525218 559906 525454
rect 560142 525218 560226 525454
rect 560462 525218 570146 525454
rect 570382 525218 570466 525454
rect 570702 525218 580386 525454
rect 580622 525218 580706 525454
rect 580942 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 6946 525134
rect 7182 524898 7266 525134
rect 7502 524898 28450 525134
rect 28686 524898 38690 525134
rect 38926 524898 48930 525134
rect 49166 524898 59170 525134
rect 59406 524898 69410 525134
rect 69646 524898 79650 525134
rect 79886 524898 89890 525134
rect 90126 524898 100130 525134
rect 100366 524898 110370 525134
rect 110606 524898 120610 525134
rect 120846 524898 130850 525134
rect 131086 524898 141090 525134
rect 141326 524898 151330 525134
rect 151566 524898 161570 525134
rect 161806 524898 171810 525134
rect 172046 524898 182050 525134
rect 182286 524898 192290 525134
rect 192526 524898 202530 525134
rect 202766 524898 212770 525134
rect 213006 524898 223010 525134
rect 223246 524898 233250 525134
rect 233486 524898 243490 525134
rect 243726 524898 253730 525134
rect 253966 524898 263970 525134
rect 264206 524898 274210 525134
rect 274446 524898 284450 525134
rect 284686 524898 294690 525134
rect 294926 524898 304930 525134
rect 305166 524898 315170 525134
rect 315406 524898 325410 525134
rect 325646 524898 335650 525134
rect 335886 524898 345890 525134
rect 346126 524898 356130 525134
rect 356366 524898 366370 525134
rect 366606 524898 376610 525134
rect 376846 524898 386850 525134
rect 387086 524898 397090 525134
rect 397326 524898 407330 525134
rect 407566 524898 417570 525134
rect 417806 524898 427810 525134
rect 428046 524898 438050 525134
rect 438286 524898 448290 525134
rect 448526 524898 458530 525134
rect 458766 524898 468770 525134
rect 469006 524898 479010 525134
rect 479246 524898 489250 525134
rect 489486 524898 499490 525134
rect 499726 524898 509730 525134
rect 509966 524898 519970 525134
rect 520206 524898 530210 525134
rect 530446 524898 549666 525134
rect 549902 524898 549986 525134
rect 550222 524898 559906 525134
rect 560142 524898 560226 525134
rect 560462 524898 570146 525134
rect 570382 524898 570466 525134
rect 570702 524898 580386 525134
rect 580622 524898 580706 525134
rect 580942 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 545466 518614
rect 545702 518378 545786 518614
rect 546022 518378 555706 518614
rect 555942 518378 556026 518614
rect 556262 518378 565946 518614
rect 566182 518378 566266 518614
rect 566502 518378 576186 518614
rect 576422 518378 576506 518614
rect 576742 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 545466 518294
rect 545702 518058 545786 518294
rect 546022 518058 555706 518294
rect 555942 518058 556026 518294
rect 556262 518058 565946 518294
rect 566182 518058 566266 518294
rect 566502 518058 576186 518294
rect 576422 518058 576506 518294
rect 576742 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 541746 514894
rect 541982 514658 542066 514894
rect 542302 514658 551986 514894
rect 552222 514658 552306 514894
rect 552542 514658 562226 514894
rect 562462 514658 562546 514894
rect 562782 514658 572466 514894
rect 572702 514658 572786 514894
rect 573022 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 541746 514574
rect 541982 514338 542066 514574
rect 542302 514338 551986 514574
rect 552222 514338 552306 514574
rect 552542 514338 562226 514574
rect 562462 514338 562546 514574
rect 562782 514338 572466 514574
rect 572702 514338 572786 514574
rect 573022 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 15786 511174
rect 16022 510938 16106 511174
rect 16342 510938 548266 511174
rect 548502 510938 548586 511174
rect 548822 510938 558506 511174
rect 558742 510938 558826 511174
rect 559062 510938 568746 511174
rect 568982 510938 569066 511174
rect 569302 510938 578986 511174
rect 579222 510938 579306 511174
rect 579542 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 15786 510854
rect 16022 510618 16106 510854
rect 16342 510618 548266 510854
rect 548502 510618 548586 510854
rect 548822 510618 558506 510854
rect 558742 510618 558826 510854
rect 559062 510618 568746 510854
rect 568982 510618 569066 510854
rect 569302 510618 578986 510854
rect 579222 510618 579306 510854
rect 579542 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 12066 507454
rect 12302 507218 12386 507454
rect 12622 507218 23330 507454
rect 23566 507218 33570 507454
rect 33806 507218 43810 507454
rect 44046 507218 54050 507454
rect 54286 507218 64290 507454
rect 64526 507218 74530 507454
rect 74766 507218 84770 507454
rect 85006 507218 95010 507454
rect 95246 507218 105250 507454
rect 105486 507218 115490 507454
rect 115726 507218 125730 507454
rect 125966 507218 135970 507454
rect 136206 507218 146210 507454
rect 146446 507218 156450 507454
rect 156686 507218 166690 507454
rect 166926 507218 176930 507454
rect 177166 507218 187170 507454
rect 187406 507218 197410 507454
rect 197646 507218 207650 507454
rect 207886 507218 217890 507454
rect 218126 507218 228130 507454
rect 228366 507218 238370 507454
rect 238606 507218 248610 507454
rect 248846 507218 258850 507454
rect 259086 507218 269090 507454
rect 269326 507218 279330 507454
rect 279566 507218 289570 507454
rect 289806 507218 299810 507454
rect 300046 507218 310050 507454
rect 310286 507218 320290 507454
rect 320526 507218 330530 507454
rect 330766 507218 340770 507454
rect 341006 507218 351010 507454
rect 351246 507218 361250 507454
rect 361486 507218 371490 507454
rect 371726 507218 381730 507454
rect 381966 507218 391970 507454
rect 392206 507218 402210 507454
rect 402446 507218 412450 507454
rect 412686 507218 422690 507454
rect 422926 507218 432930 507454
rect 433166 507218 443170 507454
rect 443406 507218 453410 507454
rect 453646 507218 463650 507454
rect 463886 507218 473890 507454
rect 474126 507218 484130 507454
rect 484366 507218 494370 507454
rect 494606 507218 504610 507454
rect 504846 507218 514850 507454
rect 515086 507218 525090 507454
rect 525326 507218 535330 507454
rect 535566 507218 544546 507454
rect 544782 507218 544866 507454
rect 545102 507218 554786 507454
rect 555022 507218 555106 507454
rect 555342 507218 565026 507454
rect 565262 507218 565346 507454
rect 565582 507218 575266 507454
rect 575502 507218 575586 507454
rect 575822 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 12066 507134
rect 12302 506898 12386 507134
rect 12622 506898 23330 507134
rect 23566 506898 33570 507134
rect 33806 506898 43810 507134
rect 44046 506898 54050 507134
rect 54286 506898 64290 507134
rect 64526 506898 74530 507134
rect 74766 506898 84770 507134
rect 85006 506898 95010 507134
rect 95246 506898 105250 507134
rect 105486 506898 115490 507134
rect 115726 506898 125730 507134
rect 125966 506898 135970 507134
rect 136206 506898 146210 507134
rect 146446 506898 156450 507134
rect 156686 506898 166690 507134
rect 166926 506898 176930 507134
rect 177166 506898 187170 507134
rect 187406 506898 197410 507134
rect 197646 506898 207650 507134
rect 207886 506898 217890 507134
rect 218126 506898 228130 507134
rect 228366 506898 238370 507134
rect 238606 506898 248610 507134
rect 248846 506898 258850 507134
rect 259086 506898 269090 507134
rect 269326 506898 279330 507134
rect 279566 506898 289570 507134
rect 289806 506898 299810 507134
rect 300046 506898 310050 507134
rect 310286 506898 320290 507134
rect 320526 506898 330530 507134
rect 330766 506898 340770 507134
rect 341006 506898 351010 507134
rect 351246 506898 361250 507134
rect 361486 506898 371490 507134
rect 371726 506898 381730 507134
rect 381966 506898 391970 507134
rect 392206 506898 402210 507134
rect 402446 506898 412450 507134
rect 412686 506898 422690 507134
rect 422926 506898 432930 507134
rect 433166 506898 443170 507134
rect 443406 506898 453410 507134
rect 453646 506898 463650 507134
rect 463886 506898 473890 507134
rect 474126 506898 484130 507134
rect 484366 506898 494370 507134
rect 494606 506898 504610 507134
rect 504846 506898 514850 507134
rect 515086 506898 525090 507134
rect 525326 506898 535330 507134
rect 535566 506898 544546 507134
rect 544782 506898 544866 507134
rect 545102 506898 554786 507134
rect 555022 506898 555106 507134
rect 555342 506898 565026 507134
rect 565262 506898 565346 507134
rect 565582 506898 575266 507134
rect 575502 506898 575586 507134
rect 575822 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 550586 500614
rect 550822 500378 550906 500614
rect 551142 500378 560826 500614
rect 561062 500378 561146 500614
rect 561382 500378 571066 500614
rect 571302 500378 571386 500614
rect 571622 500378 581306 500614
rect 581542 500378 581626 500614
rect 581862 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 550586 500294
rect 550822 500058 550906 500294
rect 551142 500058 560826 500294
rect 561062 500058 561146 500294
rect 561382 500058 571066 500294
rect 571302 500058 571386 500294
rect 571622 500058 581306 500294
rect 581542 500058 581626 500294
rect 581862 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 14386 496894
rect 14622 496658 14706 496894
rect 14942 496658 546866 496894
rect 547102 496658 547186 496894
rect 547422 496658 557106 496894
rect 557342 496658 557426 496894
rect 557662 496658 567346 496894
rect 567582 496658 567666 496894
rect 567902 496658 577586 496894
rect 577822 496658 577906 496894
rect 578142 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 14386 496574
rect 14622 496338 14706 496574
rect 14942 496338 546866 496574
rect 547102 496338 547186 496574
rect 547422 496338 557106 496574
rect 557342 496338 557426 496574
rect 557662 496338 567346 496574
rect 567582 496338 567666 496574
rect 567902 496338 577586 496574
rect 577822 496338 577906 496574
rect 578142 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 10666 493174
rect 10902 492938 10986 493174
rect 11222 492938 543146 493174
rect 543382 492938 543466 493174
rect 543702 492938 553386 493174
rect 553622 492938 553706 493174
rect 553942 492938 563626 493174
rect 563862 492938 563946 493174
rect 564182 492938 573866 493174
rect 574102 492938 574186 493174
rect 574422 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 10666 492854
rect 10902 492618 10986 492854
rect 11222 492618 543146 492854
rect 543382 492618 543466 492854
rect 543702 492618 553386 492854
rect 553622 492618 553706 492854
rect 553942 492618 563626 492854
rect 563862 492618 563946 492854
rect 564182 492618 573866 492854
rect 574102 492618 574186 492854
rect 574422 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 6946 489454
rect 7182 489218 7266 489454
rect 7502 489218 28450 489454
rect 28686 489218 38690 489454
rect 38926 489218 48930 489454
rect 49166 489218 59170 489454
rect 59406 489218 69410 489454
rect 69646 489218 79650 489454
rect 79886 489218 89890 489454
rect 90126 489218 100130 489454
rect 100366 489218 110370 489454
rect 110606 489218 120610 489454
rect 120846 489218 130850 489454
rect 131086 489218 141090 489454
rect 141326 489218 151330 489454
rect 151566 489218 161570 489454
rect 161806 489218 171810 489454
rect 172046 489218 182050 489454
rect 182286 489218 192290 489454
rect 192526 489218 202530 489454
rect 202766 489218 212770 489454
rect 213006 489218 223010 489454
rect 223246 489218 233250 489454
rect 233486 489218 243490 489454
rect 243726 489218 253730 489454
rect 253966 489218 263970 489454
rect 264206 489218 274210 489454
rect 274446 489218 284450 489454
rect 284686 489218 294690 489454
rect 294926 489218 304930 489454
rect 305166 489218 315170 489454
rect 315406 489218 325410 489454
rect 325646 489218 335650 489454
rect 335886 489218 345890 489454
rect 346126 489218 356130 489454
rect 356366 489218 366370 489454
rect 366606 489218 376610 489454
rect 376846 489218 386850 489454
rect 387086 489218 397090 489454
rect 397326 489218 407330 489454
rect 407566 489218 417570 489454
rect 417806 489218 427810 489454
rect 428046 489218 438050 489454
rect 438286 489218 448290 489454
rect 448526 489218 458530 489454
rect 458766 489218 468770 489454
rect 469006 489218 479010 489454
rect 479246 489218 489250 489454
rect 489486 489218 499490 489454
rect 499726 489218 509730 489454
rect 509966 489218 519970 489454
rect 520206 489218 530210 489454
rect 530446 489218 549666 489454
rect 549902 489218 549986 489454
rect 550222 489218 559906 489454
rect 560142 489218 560226 489454
rect 560462 489218 570146 489454
rect 570382 489218 570466 489454
rect 570702 489218 580386 489454
rect 580622 489218 580706 489454
rect 580942 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 6946 489134
rect 7182 488898 7266 489134
rect 7502 488898 28450 489134
rect 28686 488898 38690 489134
rect 38926 488898 48930 489134
rect 49166 488898 59170 489134
rect 59406 488898 69410 489134
rect 69646 488898 79650 489134
rect 79886 488898 89890 489134
rect 90126 488898 100130 489134
rect 100366 488898 110370 489134
rect 110606 488898 120610 489134
rect 120846 488898 130850 489134
rect 131086 488898 141090 489134
rect 141326 488898 151330 489134
rect 151566 488898 161570 489134
rect 161806 488898 171810 489134
rect 172046 488898 182050 489134
rect 182286 488898 192290 489134
rect 192526 488898 202530 489134
rect 202766 488898 212770 489134
rect 213006 488898 223010 489134
rect 223246 488898 233250 489134
rect 233486 488898 243490 489134
rect 243726 488898 253730 489134
rect 253966 488898 263970 489134
rect 264206 488898 274210 489134
rect 274446 488898 284450 489134
rect 284686 488898 294690 489134
rect 294926 488898 304930 489134
rect 305166 488898 315170 489134
rect 315406 488898 325410 489134
rect 325646 488898 335650 489134
rect 335886 488898 345890 489134
rect 346126 488898 356130 489134
rect 356366 488898 366370 489134
rect 366606 488898 376610 489134
rect 376846 488898 386850 489134
rect 387086 488898 397090 489134
rect 397326 488898 407330 489134
rect 407566 488898 417570 489134
rect 417806 488898 427810 489134
rect 428046 488898 438050 489134
rect 438286 488898 448290 489134
rect 448526 488898 458530 489134
rect 458766 488898 468770 489134
rect 469006 488898 479010 489134
rect 479246 488898 489250 489134
rect 489486 488898 499490 489134
rect 499726 488898 509730 489134
rect 509966 488898 519970 489134
rect 520206 488898 530210 489134
rect 530446 488898 549666 489134
rect 549902 488898 549986 489134
rect 550222 488898 559906 489134
rect 560142 488898 560226 489134
rect 560462 488898 570146 489134
rect 570382 488898 570466 489134
rect 570702 488898 580386 489134
rect 580622 488898 580706 489134
rect 580942 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 545466 482614
rect 545702 482378 545786 482614
rect 546022 482378 555706 482614
rect 555942 482378 556026 482614
rect 556262 482378 565946 482614
rect 566182 482378 566266 482614
rect 566502 482378 576186 482614
rect 576422 482378 576506 482614
rect 576742 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 545466 482294
rect 545702 482058 545786 482294
rect 546022 482058 555706 482294
rect 555942 482058 556026 482294
rect 556262 482058 565946 482294
rect 566182 482058 566266 482294
rect 566502 482058 576186 482294
rect 576422 482058 576506 482294
rect 576742 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 541746 478894
rect 541982 478658 542066 478894
rect 542302 478658 551986 478894
rect 552222 478658 552306 478894
rect 552542 478658 562226 478894
rect 562462 478658 562546 478894
rect 562782 478658 572466 478894
rect 572702 478658 572786 478894
rect 573022 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 541746 478574
rect 541982 478338 542066 478574
rect 542302 478338 551986 478574
rect 552222 478338 552306 478574
rect 552542 478338 562226 478574
rect 562462 478338 562546 478574
rect 562782 478338 572466 478574
rect 572702 478338 572786 478574
rect 573022 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 15786 475174
rect 16022 474938 16106 475174
rect 16342 474938 548266 475174
rect 548502 474938 548586 475174
rect 548822 474938 558506 475174
rect 558742 474938 558826 475174
rect 559062 474938 568746 475174
rect 568982 474938 569066 475174
rect 569302 474938 578986 475174
rect 579222 474938 579306 475174
rect 579542 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 15786 474854
rect 16022 474618 16106 474854
rect 16342 474618 548266 474854
rect 548502 474618 548586 474854
rect 548822 474618 558506 474854
rect 558742 474618 558826 474854
rect 559062 474618 568746 474854
rect 568982 474618 569066 474854
rect 569302 474618 578986 474854
rect 579222 474618 579306 474854
rect 579542 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 12066 471454
rect 12302 471218 12386 471454
rect 12622 471218 23330 471454
rect 23566 471218 33570 471454
rect 33806 471218 43810 471454
rect 44046 471218 54050 471454
rect 54286 471218 64290 471454
rect 64526 471218 74530 471454
rect 74766 471218 84770 471454
rect 85006 471218 95010 471454
rect 95246 471218 105250 471454
rect 105486 471218 115490 471454
rect 115726 471218 125730 471454
rect 125966 471218 135970 471454
rect 136206 471218 146210 471454
rect 146446 471218 156450 471454
rect 156686 471218 166690 471454
rect 166926 471218 176930 471454
rect 177166 471218 187170 471454
rect 187406 471218 197410 471454
rect 197646 471218 207650 471454
rect 207886 471218 217890 471454
rect 218126 471218 228130 471454
rect 228366 471218 238370 471454
rect 238606 471218 248610 471454
rect 248846 471218 258850 471454
rect 259086 471218 269090 471454
rect 269326 471218 279330 471454
rect 279566 471218 289570 471454
rect 289806 471218 299810 471454
rect 300046 471218 310050 471454
rect 310286 471218 320290 471454
rect 320526 471218 330530 471454
rect 330766 471218 340770 471454
rect 341006 471218 351010 471454
rect 351246 471218 361250 471454
rect 361486 471218 371490 471454
rect 371726 471218 381730 471454
rect 381966 471218 391970 471454
rect 392206 471218 402210 471454
rect 402446 471218 412450 471454
rect 412686 471218 422690 471454
rect 422926 471218 432930 471454
rect 433166 471218 443170 471454
rect 443406 471218 453410 471454
rect 453646 471218 463650 471454
rect 463886 471218 473890 471454
rect 474126 471218 484130 471454
rect 484366 471218 494370 471454
rect 494606 471218 504610 471454
rect 504846 471218 514850 471454
rect 515086 471218 525090 471454
rect 525326 471218 535330 471454
rect 535566 471218 544546 471454
rect 544782 471218 544866 471454
rect 545102 471218 554786 471454
rect 555022 471218 555106 471454
rect 555342 471218 565026 471454
rect 565262 471218 565346 471454
rect 565582 471218 575266 471454
rect 575502 471218 575586 471454
rect 575822 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 12066 471134
rect 12302 470898 12386 471134
rect 12622 470898 23330 471134
rect 23566 470898 33570 471134
rect 33806 470898 43810 471134
rect 44046 470898 54050 471134
rect 54286 470898 64290 471134
rect 64526 470898 74530 471134
rect 74766 470898 84770 471134
rect 85006 470898 95010 471134
rect 95246 470898 105250 471134
rect 105486 470898 115490 471134
rect 115726 470898 125730 471134
rect 125966 470898 135970 471134
rect 136206 470898 146210 471134
rect 146446 470898 156450 471134
rect 156686 470898 166690 471134
rect 166926 470898 176930 471134
rect 177166 470898 187170 471134
rect 187406 470898 197410 471134
rect 197646 470898 207650 471134
rect 207886 470898 217890 471134
rect 218126 470898 228130 471134
rect 228366 470898 238370 471134
rect 238606 470898 248610 471134
rect 248846 470898 258850 471134
rect 259086 470898 269090 471134
rect 269326 470898 279330 471134
rect 279566 470898 289570 471134
rect 289806 470898 299810 471134
rect 300046 470898 310050 471134
rect 310286 470898 320290 471134
rect 320526 470898 330530 471134
rect 330766 470898 340770 471134
rect 341006 470898 351010 471134
rect 351246 470898 361250 471134
rect 361486 470898 371490 471134
rect 371726 470898 381730 471134
rect 381966 470898 391970 471134
rect 392206 470898 402210 471134
rect 402446 470898 412450 471134
rect 412686 470898 422690 471134
rect 422926 470898 432930 471134
rect 433166 470898 443170 471134
rect 443406 470898 453410 471134
rect 453646 470898 463650 471134
rect 463886 470898 473890 471134
rect 474126 470898 484130 471134
rect 484366 470898 494370 471134
rect 494606 470898 504610 471134
rect 504846 470898 514850 471134
rect 515086 470898 525090 471134
rect 525326 470898 535330 471134
rect 535566 470898 544546 471134
rect 544782 470898 544866 471134
rect 545102 470898 554786 471134
rect 555022 470898 555106 471134
rect 555342 470898 565026 471134
rect 565262 470898 565346 471134
rect 565582 470898 575266 471134
rect 575502 470898 575586 471134
rect 575822 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 550586 464614
rect 550822 464378 550906 464614
rect 551142 464378 560826 464614
rect 561062 464378 561146 464614
rect 561382 464378 571066 464614
rect 571302 464378 571386 464614
rect 571622 464378 581306 464614
rect 581542 464378 581626 464614
rect 581862 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 550586 464294
rect 550822 464058 550906 464294
rect 551142 464058 560826 464294
rect 561062 464058 561146 464294
rect 561382 464058 571066 464294
rect 571302 464058 571386 464294
rect 571622 464058 581306 464294
rect 581542 464058 581626 464294
rect 581862 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 14386 460894
rect 14622 460658 14706 460894
rect 14942 460658 546866 460894
rect 547102 460658 547186 460894
rect 547422 460658 557106 460894
rect 557342 460658 557426 460894
rect 557662 460658 567346 460894
rect 567582 460658 567666 460894
rect 567902 460658 577586 460894
rect 577822 460658 577906 460894
rect 578142 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 14386 460574
rect 14622 460338 14706 460574
rect 14942 460338 546866 460574
rect 547102 460338 547186 460574
rect 547422 460338 557106 460574
rect 557342 460338 557426 460574
rect 557662 460338 567346 460574
rect 567582 460338 567666 460574
rect 567902 460338 577586 460574
rect 577822 460338 577906 460574
rect 578142 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 10666 457174
rect 10902 456938 10986 457174
rect 11222 456938 543146 457174
rect 543382 456938 543466 457174
rect 543702 456938 553386 457174
rect 553622 456938 553706 457174
rect 553942 456938 563626 457174
rect 563862 456938 563946 457174
rect 564182 456938 573866 457174
rect 574102 456938 574186 457174
rect 574422 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 10666 456854
rect 10902 456618 10986 456854
rect 11222 456618 543146 456854
rect 543382 456618 543466 456854
rect 543702 456618 553386 456854
rect 553622 456618 553706 456854
rect 553942 456618 563626 456854
rect 563862 456618 563946 456854
rect 564182 456618 573866 456854
rect 574102 456618 574186 456854
rect 574422 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 6946 453454
rect 7182 453218 7266 453454
rect 7502 453218 28450 453454
rect 28686 453218 38690 453454
rect 38926 453218 48930 453454
rect 49166 453218 59170 453454
rect 59406 453218 69410 453454
rect 69646 453218 79650 453454
rect 79886 453218 89890 453454
rect 90126 453218 100130 453454
rect 100366 453218 110370 453454
rect 110606 453218 120610 453454
rect 120846 453218 130850 453454
rect 131086 453218 141090 453454
rect 141326 453218 151330 453454
rect 151566 453218 161570 453454
rect 161806 453218 171810 453454
rect 172046 453218 182050 453454
rect 182286 453218 192290 453454
rect 192526 453218 202530 453454
rect 202766 453218 212770 453454
rect 213006 453218 223010 453454
rect 223246 453218 233250 453454
rect 233486 453218 243490 453454
rect 243726 453218 253730 453454
rect 253966 453218 263970 453454
rect 264206 453218 274210 453454
rect 274446 453218 284450 453454
rect 284686 453218 294690 453454
rect 294926 453218 304930 453454
rect 305166 453218 315170 453454
rect 315406 453218 325410 453454
rect 325646 453218 335650 453454
rect 335886 453218 345890 453454
rect 346126 453218 356130 453454
rect 356366 453218 366370 453454
rect 366606 453218 376610 453454
rect 376846 453218 386850 453454
rect 387086 453218 397090 453454
rect 397326 453218 407330 453454
rect 407566 453218 417570 453454
rect 417806 453218 427810 453454
rect 428046 453218 438050 453454
rect 438286 453218 448290 453454
rect 448526 453218 458530 453454
rect 458766 453218 468770 453454
rect 469006 453218 479010 453454
rect 479246 453218 489250 453454
rect 489486 453218 499490 453454
rect 499726 453218 509730 453454
rect 509966 453218 519970 453454
rect 520206 453218 530210 453454
rect 530446 453218 549666 453454
rect 549902 453218 549986 453454
rect 550222 453218 559906 453454
rect 560142 453218 560226 453454
rect 560462 453218 570146 453454
rect 570382 453218 570466 453454
rect 570702 453218 580386 453454
rect 580622 453218 580706 453454
rect 580942 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 6946 453134
rect 7182 452898 7266 453134
rect 7502 452898 28450 453134
rect 28686 452898 38690 453134
rect 38926 452898 48930 453134
rect 49166 452898 59170 453134
rect 59406 452898 69410 453134
rect 69646 452898 79650 453134
rect 79886 452898 89890 453134
rect 90126 452898 100130 453134
rect 100366 452898 110370 453134
rect 110606 452898 120610 453134
rect 120846 452898 130850 453134
rect 131086 452898 141090 453134
rect 141326 452898 151330 453134
rect 151566 452898 161570 453134
rect 161806 452898 171810 453134
rect 172046 452898 182050 453134
rect 182286 452898 192290 453134
rect 192526 452898 202530 453134
rect 202766 452898 212770 453134
rect 213006 452898 223010 453134
rect 223246 452898 233250 453134
rect 233486 452898 243490 453134
rect 243726 452898 253730 453134
rect 253966 452898 263970 453134
rect 264206 452898 274210 453134
rect 274446 452898 284450 453134
rect 284686 452898 294690 453134
rect 294926 452898 304930 453134
rect 305166 452898 315170 453134
rect 315406 452898 325410 453134
rect 325646 452898 335650 453134
rect 335886 452898 345890 453134
rect 346126 452898 356130 453134
rect 356366 452898 366370 453134
rect 366606 452898 376610 453134
rect 376846 452898 386850 453134
rect 387086 452898 397090 453134
rect 397326 452898 407330 453134
rect 407566 452898 417570 453134
rect 417806 452898 427810 453134
rect 428046 452898 438050 453134
rect 438286 452898 448290 453134
rect 448526 452898 458530 453134
rect 458766 452898 468770 453134
rect 469006 452898 479010 453134
rect 479246 452898 489250 453134
rect 489486 452898 499490 453134
rect 499726 452898 509730 453134
rect 509966 452898 519970 453134
rect 520206 452898 530210 453134
rect 530446 452898 549666 453134
rect 549902 452898 549986 453134
rect 550222 452898 559906 453134
rect 560142 452898 560226 453134
rect 560462 452898 570146 453134
rect 570382 452898 570466 453134
rect 570702 452898 580386 453134
rect 580622 452898 580706 453134
rect 580942 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 545466 446614
rect 545702 446378 545786 446614
rect 546022 446378 555706 446614
rect 555942 446378 556026 446614
rect 556262 446378 565946 446614
rect 566182 446378 566266 446614
rect 566502 446378 576186 446614
rect 576422 446378 576506 446614
rect 576742 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 545466 446294
rect 545702 446058 545786 446294
rect 546022 446058 555706 446294
rect 555942 446058 556026 446294
rect 556262 446058 565946 446294
rect 566182 446058 566266 446294
rect 566502 446058 576186 446294
rect 576422 446058 576506 446294
rect 576742 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 541746 442894
rect 541982 442658 542066 442894
rect 542302 442658 551986 442894
rect 552222 442658 552306 442894
rect 552542 442658 562226 442894
rect 562462 442658 562546 442894
rect 562782 442658 572466 442894
rect 572702 442658 572786 442894
rect 573022 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 541746 442574
rect 541982 442338 542066 442574
rect 542302 442338 551986 442574
rect 552222 442338 552306 442574
rect 552542 442338 562226 442574
rect 562462 442338 562546 442574
rect 562782 442338 572466 442574
rect 572702 442338 572786 442574
rect 573022 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 15786 439174
rect 16022 438938 16106 439174
rect 16342 438938 548266 439174
rect 548502 438938 548586 439174
rect 548822 438938 558506 439174
rect 558742 438938 558826 439174
rect 559062 438938 568746 439174
rect 568982 438938 569066 439174
rect 569302 438938 578986 439174
rect 579222 438938 579306 439174
rect 579542 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 15786 438854
rect 16022 438618 16106 438854
rect 16342 438618 548266 438854
rect 548502 438618 548586 438854
rect 548822 438618 558506 438854
rect 558742 438618 558826 438854
rect 559062 438618 568746 438854
rect 568982 438618 569066 438854
rect 569302 438618 578986 438854
rect 579222 438618 579306 438854
rect 579542 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 12066 435454
rect 12302 435218 12386 435454
rect 12622 435218 23330 435454
rect 23566 435218 33570 435454
rect 33806 435218 43810 435454
rect 44046 435218 54050 435454
rect 54286 435218 64290 435454
rect 64526 435218 74530 435454
rect 74766 435218 84770 435454
rect 85006 435218 95010 435454
rect 95246 435218 105250 435454
rect 105486 435218 115490 435454
rect 115726 435218 125730 435454
rect 125966 435218 135970 435454
rect 136206 435218 146210 435454
rect 146446 435218 156450 435454
rect 156686 435218 166690 435454
rect 166926 435218 176930 435454
rect 177166 435218 187170 435454
rect 187406 435218 197410 435454
rect 197646 435218 207650 435454
rect 207886 435218 217890 435454
rect 218126 435218 228130 435454
rect 228366 435218 238370 435454
rect 238606 435218 248610 435454
rect 248846 435218 258850 435454
rect 259086 435218 269090 435454
rect 269326 435218 279330 435454
rect 279566 435218 289570 435454
rect 289806 435218 299810 435454
rect 300046 435218 310050 435454
rect 310286 435218 320290 435454
rect 320526 435218 330530 435454
rect 330766 435218 340770 435454
rect 341006 435218 351010 435454
rect 351246 435218 361250 435454
rect 361486 435218 371490 435454
rect 371726 435218 381730 435454
rect 381966 435218 391970 435454
rect 392206 435218 402210 435454
rect 402446 435218 412450 435454
rect 412686 435218 422690 435454
rect 422926 435218 432930 435454
rect 433166 435218 443170 435454
rect 443406 435218 453410 435454
rect 453646 435218 463650 435454
rect 463886 435218 473890 435454
rect 474126 435218 484130 435454
rect 484366 435218 494370 435454
rect 494606 435218 504610 435454
rect 504846 435218 514850 435454
rect 515086 435218 525090 435454
rect 525326 435218 535330 435454
rect 535566 435218 544546 435454
rect 544782 435218 544866 435454
rect 545102 435218 554786 435454
rect 555022 435218 555106 435454
rect 555342 435218 565026 435454
rect 565262 435218 565346 435454
rect 565582 435218 575266 435454
rect 575502 435218 575586 435454
rect 575822 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 12066 435134
rect 12302 434898 12386 435134
rect 12622 434898 23330 435134
rect 23566 434898 33570 435134
rect 33806 434898 43810 435134
rect 44046 434898 54050 435134
rect 54286 434898 64290 435134
rect 64526 434898 74530 435134
rect 74766 434898 84770 435134
rect 85006 434898 95010 435134
rect 95246 434898 105250 435134
rect 105486 434898 115490 435134
rect 115726 434898 125730 435134
rect 125966 434898 135970 435134
rect 136206 434898 146210 435134
rect 146446 434898 156450 435134
rect 156686 434898 166690 435134
rect 166926 434898 176930 435134
rect 177166 434898 187170 435134
rect 187406 434898 197410 435134
rect 197646 434898 207650 435134
rect 207886 434898 217890 435134
rect 218126 434898 228130 435134
rect 228366 434898 238370 435134
rect 238606 434898 248610 435134
rect 248846 434898 258850 435134
rect 259086 434898 269090 435134
rect 269326 434898 279330 435134
rect 279566 434898 289570 435134
rect 289806 434898 299810 435134
rect 300046 434898 310050 435134
rect 310286 434898 320290 435134
rect 320526 434898 330530 435134
rect 330766 434898 340770 435134
rect 341006 434898 351010 435134
rect 351246 434898 361250 435134
rect 361486 434898 371490 435134
rect 371726 434898 381730 435134
rect 381966 434898 391970 435134
rect 392206 434898 402210 435134
rect 402446 434898 412450 435134
rect 412686 434898 422690 435134
rect 422926 434898 432930 435134
rect 433166 434898 443170 435134
rect 443406 434898 453410 435134
rect 453646 434898 463650 435134
rect 463886 434898 473890 435134
rect 474126 434898 484130 435134
rect 484366 434898 494370 435134
rect 494606 434898 504610 435134
rect 504846 434898 514850 435134
rect 515086 434898 525090 435134
rect 525326 434898 535330 435134
rect 535566 434898 544546 435134
rect 544782 434898 544866 435134
rect 545102 434898 554786 435134
rect 555022 434898 555106 435134
rect 555342 434898 565026 435134
rect 565262 434898 565346 435134
rect 565582 434898 575266 435134
rect 575502 434898 575586 435134
rect 575822 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 550586 428614
rect 550822 428378 550906 428614
rect 551142 428378 560826 428614
rect 561062 428378 561146 428614
rect 561382 428378 571066 428614
rect 571302 428378 571386 428614
rect 571622 428378 581306 428614
rect 581542 428378 581626 428614
rect 581862 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 550586 428294
rect 550822 428058 550906 428294
rect 551142 428058 560826 428294
rect 561062 428058 561146 428294
rect 561382 428058 571066 428294
rect 571302 428058 571386 428294
rect 571622 428058 581306 428294
rect 581542 428058 581626 428294
rect 581862 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 14386 424894
rect 14622 424658 14706 424894
rect 14942 424658 546866 424894
rect 547102 424658 547186 424894
rect 547422 424658 557106 424894
rect 557342 424658 557426 424894
rect 557662 424658 567346 424894
rect 567582 424658 567666 424894
rect 567902 424658 577586 424894
rect 577822 424658 577906 424894
rect 578142 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 14386 424574
rect 14622 424338 14706 424574
rect 14942 424338 546866 424574
rect 547102 424338 547186 424574
rect 547422 424338 557106 424574
rect 557342 424338 557426 424574
rect 557662 424338 567346 424574
rect 567582 424338 567666 424574
rect 567902 424338 577586 424574
rect 577822 424338 577906 424574
rect 578142 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 10666 421174
rect 10902 420938 10986 421174
rect 11222 420938 543146 421174
rect 543382 420938 543466 421174
rect 543702 420938 553386 421174
rect 553622 420938 553706 421174
rect 553942 420938 563626 421174
rect 563862 420938 563946 421174
rect 564182 420938 573866 421174
rect 574102 420938 574186 421174
rect 574422 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 10666 420854
rect 10902 420618 10986 420854
rect 11222 420618 543146 420854
rect 543382 420618 543466 420854
rect 543702 420618 553386 420854
rect 553622 420618 553706 420854
rect 553942 420618 563626 420854
rect 563862 420618 563946 420854
rect 564182 420618 573866 420854
rect 574102 420618 574186 420854
rect 574422 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 6946 417454
rect 7182 417218 7266 417454
rect 7502 417218 28450 417454
rect 28686 417218 38690 417454
rect 38926 417218 48930 417454
rect 49166 417218 59170 417454
rect 59406 417218 69410 417454
rect 69646 417218 79650 417454
rect 79886 417218 89890 417454
rect 90126 417218 100130 417454
rect 100366 417218 110370 417454
rect 110606 417218 120610 417454
rect 120846 417218 130850 417454
rect 131086 417218 141090 417454
rect 141326 417218 151330 417454
rect 151566 417218 161570 417454
rect 161806 417218 171810 417454
rect 172046 417218 182050 417454
rect 182286 417218 192290 417454
rect 192526 417218 202530 417454
rect 202766 417218 212770 417454
rect 213006 417218 223010 417454
rect 223246 417218 233250 417454
rect 233486 417218 243490 417454
rect 243726 417218 253730 417454
rect 253966 417218 263970 417454
rect 264206 417218 274210 417454
rect 274446 417218 284450 417454
rect 284686 417218 294690 417454
rect 294926 417218 304930 417454
rect 305166 417218 315170 417454
rect 315406 417218 325410 417454
rect 325646 417218 335650 417454
rect 335886 417218 345890 417454
rect 346126 417218 356130 417454
rect 356366 417218 366370 417454
rect 366606 417218 376610 417454
rect 376846 417218 386850 417454
rect 387086 417218 397090 417454
rect 397326 417218 407330 417454
rect 407566 417218 417570 417454
rect 417806 417218 427810 417454
rect 428046 417218 438050 417454
rect 438286 417218 448290 417454
rect 448526 417218 458530 417454
rect 458766 417218 468770 417454
rect 469006 417218 479010 417454
rect 479246 417218 489250 417454
rect 489486 417218 499490 417454
rect 499726 417218 509730 417454
rect 509966 417218 519970 417454
rect 520206 417218 530210 417454
rect 530446 417218 549666 417454
rect 549902 417218 549986 417454
rect 550222 417218 559906 417454
rect 560142 417218 560226 417454
rect 560462 417218 570146 417454
rect 570382 417218 570466 417454
rect 570702 417218 580386 417454
rect 580622 417218 580706 417454
rect 580942 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 6946 417134
rect 7182 416898 7266 417134
rect 7502 416898 28450 417134
rect 28686 416898 38690 417134
rect 38926 416898 48930 417134
rect 49166 416898 59170 417134
rect 59406 416898 69410 417134
rect 69646 416898 79650 417134
rect 79886 416898 89890 417134
rect 90126 416898 100130 417134
rect 100366 416898 110370 417134
rect 110606 416898 120610 417134
rect 120846 416898 130850 417134
rect 131086 416898 141090 417134
rect 141326 416898 151330 417134
rect 151566 416898 161570 417134
rect 161806 416898 171810 417134
rect 172046 416898 182050 417134
rect 182286 416898 192290 417134
rect 192526 416898 202530 417134
rect 202766 416898 212770 417134
rect 213006 416898 223010 417134
rect 223246 416898 233250 417134
rect 233486 416898 243490 417134
rect 243726 416898 253730 417134
rect 253966 416898 263970 417134
rect 264206 416898 274210 417134
rect 274446 416898 284450 417134
rect 284686 416898 294690 417134
rect 294926 416898 304930 417134
rect 305166 416898 315170 417134
rect 315406 416898 325410 417134
rect 325646 416898 335650 417134
rect 335886 416898 345890 417134
rect 346126 416898 356130 417134
rect 356366 416898 366370 417134
rect 366606 416898 376610 417134
rect 376846 416898 386850 417134
rect 387086 416898 397090 417134
rect 397326 416898 407330 417134
rect 407566 416898 417570 417134
rect 417806 416898 427810 417134
rect 428046 416898 438050 417134
rect 438286 416898 448290 417134
rect 448526 416898 458530 417134
rect 458766 416898 468770 417134
rect 469006 416898 479010 417134
rect 479246 416898 489250 417134
rect 489486 416898 499490 417134
rect 499726 416898 509730 417134
rect 509966 416898 519970 417134
rect 520206 416898 530210 417134
rect 530446 416898 549666 417134
rect 549902 416898 549986 417134
rect 550222 416898 559906 417134
rect 560142 416898 560226 417134
rect 560462 416898 570146 417134
rect 570382 416898 570466 417134
rect 570702 416898 580386 417134
rect 580622 416898 580706 417134
rect 580942 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 545466 410614
rect 545702 410378 545786 410614
rect 546022 410378 555706 410614
rect 555942 410378 556026 410614
rect 556262 410378 565946 410614
rect 566182 410378 566266 410614
rect 566502 410378 576186 410614
rect 576422 410378 576506 410614
rect 576742 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 545466 410294
rect 545702 410058 545786 410294
rect 546022 410058 555706 410294
rect 555942 410058 556026 410294
rect 556262 410058 565946 410294
rect 566182 410058 566266 410294
rect 566502 410058 576186 410294
rect 576422 410058 576506 410294
rect 576742 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 541746 406894
rect 541982 406658 542066 406894
rect 542302 406658 551986 406894
rect 552222 406658 552306 406894
rect 552542 406658 562226 406894
rect 562462 406658 562546 406894
rect 562782 406658 572466 406894
rect 572702 406658 572786 406894
rect 573022 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 541746 406574
rect 541982 406338 542066 406574
rect 542302 406338 551986 406574
rect 552222 406338 552306 406574
rect 552542 406338 562226 406574
rect 562462 406338 562546 406574
rect 562782 406338 572466 406574
rect 572702 406338 572786 406574
rect 573022 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 15786 403174
rect 16022 402938 16106 403174
rect 16342 402938 548266 403174
rect 548502 402938 548586 403174
rect 548822 402938 558506 403174
rect 558742 402938 558826 403174
rect 559062 402938 568746 403174
rect 568982 402938 569066 403174
rect 569302 402938 578986 403174
rect 579222 402938 579306 403174
rect 579542 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 15786 402854
rect 16022 402618 16106 402854
rect 16342 402618 548266 402854
rect 548502 402618 548586 402854
rect 548822 402618 558506 402854
rect 558742 402618 558826 402854
rect 559062 402618 568746 402854
rect 568982 402618 569066 402854
rect 569302 402618 578986 402854
rect 579222 402618 579306 402854
rect 579542 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 12066 399454
rect 12302 399218 12386 399454
rect 12622 399218 23330 399454
rect 23566 399218 33570 399454
rect 33806 399218 43810 399454
rect 44046 399218 54050 399454
rect 54286 399218 64290 399454
rect 64526 399218 74530 399454
rect 74766 399218 84770 399454
rect 85006 399218 95010 399454
rect 95246 399218 105250 399454
rect 105486 399218 115490 399454
rect 115726 399218 125730 399454
rect 125966 399218 135970 399454
rect 136206 399218 146210 399454
rect 146446 399218 156450 399454
rect 156686 399218 166690 399454
rect 166926 399218 176930 399454
rect 177166 399218 187170 399454
rect 187406 399218 197410 399454
rect 197646 399218 207650 399454
rect 207886 399218 217890 399454
rect 218126 399218 228130 399454
rect 228366 399218 238370 399454
rect 238606 399218 248610 399454
rect 248846 399218 258850 399454
rect 259086 399218 269090 399454
rect 269326 399218 279330 399454
rect 279566 399218 289570 399454
rect 289806 399218 299810 399454
rect 300046 399218 310050 399454
rect 310286 399218 320290 399454
rect 320526 399218 330530 399454
rect 330766 399218 340770 399454
rect 341006 399218 351010 399454
rect 351246 399218 361250 399454
rect 361486 399218 371490 399454
rect 371726 399218 381730 399454
rect 381966 399218 391970 399454
rect 392206 399218 402210 399454
rect 402446 399218 412450 399454
rect 412686 399218 422690 399454
rect 422926 399218 432930 399454
rect 433166 399218 443170 399454
rect 443406 399218 453410 399454
rect 453646 399218 463650 399454
rect 463886 399218 473890 399454
rect 474126 399218 484130 399454
rect 484366 399218 494370 399454
rect 494606 399218 504610 399454
rect 504846 399218 514850 399454
rect 515086 399218 525090 399454
rect 525326 399218 535330 399454
rect 535566 399218 544546 399454
rect 544782 399218 544866 399454
rect 545102 399218 554786 399454
rect 555022 399218 555106 399454
rect 555342 399218 565026 399454
rect 565262 399218 565346 399454
rect 565582 399218 575266 399454
rect 575502 399218 575586 399454
rect 575822 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 12066 399134
rect 12302 398898 12386 399134
rect 12622 398898 23330 399134
rect 23566 398898 33570 399134
rect 33806 398898 43810 399134
rect 44046 398898 54050 399134
rect 54286 398898 64290 399134
rect 64526 398898 74530 399134
rect 74766 398898 84770 399134
rect 85006 398898 95010 399134
rect 95246 398898 105250 399134
rect 105486 398898 115490 399134
rect 115726 398898 125730 399134
rect 125966 398898 135970 399134
rect 136206 398898 146210 399134
rect 146446 398898 156450 399134
rect 156686 398898 166690 399134
rect 166926 398898 176930 399134
rect 177166 398898 187170 399134
rect 187406 398898 197410 399134
rect 197646 398898 207650 399134
rect 207886 398898 217890 399134
rect 218126 398898 228130 399134
rect 228366 398898 238370 399134
rect 238606 398898 248610 399134
rect 248846 398898 258850 399134
rect 259086 398898 269090 399134
rect 269326 398898 279330 399134
rect 279566 398898 289570 399134
rect 289806 398898 299810 399134
rect 300046 398898 310050 399134
rect 310286 398898 320290 399134
rect 320526 398898 330530 399134
rect 330766 398898 340770 399134
rect 341006 398898 351010 399134
rect 351246 398898 361250 399134
rect 361486 398898 371490 399134
rect 371726 398898 381730 399134
rect 381966 398898 391970 399134
rect 392206 398898 402210 399134
rect 402446 398898 412450 399134
rect 412686 398898 422690 399134
rect 422926 398898 432930 399134
rect 433166 398898 443170 399134
rect 443406 398898 453410 399134
rect 453646 398898 463650 399134
rect 463886 398898 473890 399134
rect 474126 398898 484130 399134
rect 484366 398898 494370 399134
rect 494606 398898 504610 399134
rect 504846 398898 514850 399134
rect 515086 398898 525090 399134
rect 525326 398898 535330 399134
rect 535566 398898 544546 399134
rect 544782 398898 544866 399134
rect 545102 398898 554786 399134
rect 555022 398898 555106 399134
rect 555342 398898 565026 399134
rect 565262 398898 565346 399134
rect 565582 398898 575266 399134
rect 575502 398898 575586 399134
rect 575822 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 550586 392614
rect 550822 392378 550906 392614
rect 551142 392378 560826 392614
rect 561062 392378 561146 392614
rect 561382 392378 571066 392614
rect 571302 392378 571386 392614
rect 571622 392378 581306 392614
rect 581542 392378 581626 392614
rect 581862 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 550586 392294
rect 550822 392058 550906 392294
rect 551142 392058 560826 392294
rect 561062 392058 561146 392294
rect 561382 392058 571066 392294
rect 571302 392058 571386 392294
rect 571622 392058 581306 392294
rect 581542 392058 581626 392294
rect 581862 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 14386 388894
rect 14622 388658 14706 388894
rect 14942 388658 546866 388894
rect 547102 388658 547186 388894
rect 547422 388658 557106 388894
rect 557342 388658 557426 388894
rect 557662 388658 567346 388894
rect 567582 388658 567666 388894
rect 567902 388658 577586 388894
rect 577822 388658 577906 388894
rect 578142 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 14386 388574
rect 14622 388338 14706 388574
rect 14942 388338 546866 388574
rect 547102 388338 547186 388574
rect 547422 388338 557106 388574
rect 557342 388338 557426 388574
rect 557662 388338 567346 388574
rect 567582 388338 567666 388574
rect 567902 388338 577586 388574
rect 577822 388338 577906 388574
rect 578142 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 10666 385174
rect 10902 384938 10986 385174
rect 11222 384938 543146 385174
rect 543382 384938 543466 385174
rect 543702 384938 553386 385174
rect 553622 384938 553706 385174
rect 553942 384938 563626 385174
rect 563862 384938 563946 385174
rect 564182 384938 573866 385174
rect 574102 384938 574186 385174
rect 574422 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 10666 384854
rect 10902 384618 10986 384854
rect 11222 384618 543146 384854
rect 543382 384618 543466 384854
rect 543702 384618 553386 384854
rect 553622 384618 553706 384854
rect 553942 384618 563626 384854
rect 563862 384618 563946 384854
rect 564182 384618 573866 384854
rect 574102 384618 574186 384854
rect 574422 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 6946 381454
rect 7182 381218 7266 381454
rect 7502 381218 28450 381454
rect 28686 381218 38690 381454
rect 38926 381218 48930 381454
rect 49166 381218 59170 381454
rect 59406 381218 69410 381454
rect 69646 381218 79650 381454
rect 79886 381218 89890 381454
rect 90126 381218 100130 381454
rect 100366 381218 110370 381454
rect 110606 381218 120610 381454
rect 120846 381218 130850 381454
rect 131086 381218 141090 381454
rect 141326 381218 151330 381454
rect 151566 381218 161570 381454
rect 161806 381218 171810 381454
rect 172046 381218 182050 381454
rect 182286 381218 192290 381454
rect 192526 381218 202530 381454
rect 202766 381218 212770 381454
rect 213006 381218 223010 381454
rect 223246 381218 233250 381454
rect 233486 381218 243490 381454
rect 243726 381218 253730 381454
rect 253966 381218 263970 381454
rect 264206 381218 274210 381454
rect 274446 381218 284450 381454
rect 284686 381218 294690 381454
rect 294926 381218 304930 381454
rect 305166 381218 315170 381454
rect 315406 381218 325410 381454
rect 325646 381218 335650 381454
rect 335886 381218 345890 381454
rect 346126 381218 356130 381454
rect 356366 381218 366370 381454
rect 366606 381218 376610 381454
rect 376846 381218 386850 381454
rect 387086 381218 397090 381454
rect 397326 381218 407330 381454
rect 407566 381218 417570 381454
rect 417806 381218 427810 381454
rect 428046 381218 438050 381454
rect 438286 381218 448290 381454
rect 448526 381218 458530 381454
rect 458766 381218 468770 381454
rect 469006 381218 479010 381454
rect 479246 381218 489250 381454
rect 489486 381218 499490 381454
rect 499726 381218 509730 381454
rect 509966 381218 519970 381454
rect 520206 381218 530210 381454
rect 530446 381218 549666 381454
rect 549902 381218 549986 381454
rect 550222 381218 559906 381454
rect 560142 381218 560226 381454
rect 560462 381218 570146 381454
rect 570382 381218 570466 381454
rect 570702 381218 580386 381454
rect 580622 381218 580706 381454
rect 580942 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 6946 381134
rect 7182 380898 7266 381134
rect 7502 380898 28450 381134
rect 28686 380898 38690 381134
rect 38926 380898 48930 381134
rect 49166 380898 59170 381134
rect 59406 380898 69410 381134
rect 69646 380898 79650 381134
rect 79886 380898 89890 381134
rect 90126 380898 100130 381134
rect 100366 380898 110370 381134
rect 110606 380898 120610 381134
rect 120846 380898 130850 381134
rect 131086 380898 141090 381134
rect 141326 380898 151330 381134
rect 151566 380898 161570 381134
rect 161806 380898 171810 381134
rect 172046 380898 182050 381134
rect 182286 380898 192290 381134
rect 192526 380898 202530 381134
rect 202766 380898 212770 381134
rect 213006 380898 223010 381134
rect 223246 380898 233250 381134
rect 233486 380898 243490 381134
rect 243726 380898 253730 381134
rect 253966 380898 263970 381134
rect 264206 380898 274210 381134
rect 274446 380898 284450 381134
rect 284686 380898 294690 381134
rect 294926 380898 304930 381134
rect 305166 380898 315170 381134
rect 315406 380898 325410 381134
rect 325646 380898 335650 381134
rect 335886 380898 345890 381134
rect 346126 380898 356130 381134
rect 356366 380898 366370 381134
rect 366606 380898 376610 381134
rect 376846 380898 386850 381134
rect 387086 380898 397090 381134
rect 397326 380898 407330 381134
rect 407566 380898 417570 381134
rect 417806 380898 427810 381134
rect 428046 380898 438050 381134
rect 438286 380898 448290 381134
rect 448526 380898 458530 381134
rect 458766 380898 468770 381134
rect 469006 380898 479010 381134
rect 479246 380898 489250 381134
rect 489486 380898 499490 381134
rect 499726 380898 509730 381134
rect 509966 380898 519970 381134
rect 520206 380898 530210 381134
rect 530446 380898 549666 381134
rect 549902 380898 549986 381134
rect 550222 380898 559906 381134
rect 560142 380898 560226 381134
rect 560462 380898 570146 381134
rect 570382 380898 570466 381134
rect 570702 380898 580386 381134
rect 580622 380898 580706 381134
rect 580942 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 545466 374614
rect 545702 374378 545786 374614
rect 546022 374378 555706 374614
rect 555942 374378 556026 374614
rect 556262 374378 565946 374614
rect 566182 374378 566266 374614
rect 566502 374378 576186 374614
rect 576422 374378 576506 374614
rect 576742 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 545466 374294
rect 545702 374058 545786 374294
rect 546022 374058 555706 374294
rect 555942 374058 556026 374294
rect 556262 374058 565946 374294
rect 566182 374058 566266 374294
rect 566502 374058 576186 374294
rect 576422 374058 576506 374294
rect 576742 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 541746 370894
rect 541982 370658 542066 370894
rect 542302 370658 551986 370894
rect 552222 370658 552306 370894
rect 552542 370658 562226 370894
rect 562462 370658 562546 370894
rect 562782 370658 572466 370894
rect 572702 370658 572786 370894
rect 573022 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 541746 370574
rect 541982 370338 542066 370574
rect 542302 370338 551986 370574
rect 552222 370338 552306 370574
rect 552542 370338 562226 370574
rect 562462 370338 562546 370574
rect 562782 370338 572466 370574
rect 572702 370338 572786 370574
rect 573022 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 15786 367174
rect 16022 366938 16106 367174
rect 16342 366938 548266 367174
rect 548502 366938 548586 367174
rect 548822 366938 558506 367174
rect 558742 366938 558826 367174
rect 559062 366938 568746 367174
rect 568982 366938 569066 367174
rect 569302 366938 578986 367174
rect 579222 366938 579306 367174
rect 579542 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 15786 366854
rect 16022 366618 16106 366854
rect 16342 366618 548266 366854
rect 548502 366618 548586 366854
rect 548822 366618 558506 366854
rect 558742 366618 558826 366854
rect 559062 366618 568746 366854
rect 568982 366618 569066 366854
rect 569302 366618 578986 366854
rect 579222 366618 579306 366854
rect 579542 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 12066 363454
rect 12302 363218 12386 363454
rect 12622 363218 23330 363454
rect 23566 363218 33570 363454
rect 33806 363218 43810 363454
rect 44046 363218 54050 363454
rect 54286 363218 64290 363454
rect 64526 363218 74530 363454
rect 74766 363218 84770 363454
rect 85006 363218 95010 363454
rect 95246 363218 105250 363454
rect 105486 363218 115490 363454
rect 115726 363218 125730 363454
rect 125966 363218 135970 363454
rect 136206 363218 146210 363454
rect 146446 363218 156450 363454
rect 156686 363218 166690 363454
rect 166926 363218 176930 363454
rect 177166 363218 187170 363454
rect 187406 363218 197410 363454
rect 197646 363218 207650 363454
rect 207886 363218 217890 363454
rect 218126 363218 228130 363454
rect 228366 363218 238370 363454
rect 238606 363218 248610 363454
rect 248846 363218 258850 363454
rect 259086 363218 269090 363454
rect 269326 363218 279330 363454
rect 279566 363218 289570 363454
rect 289806 363218 299810 363454
rect 300046 363218 310050 363454
rect 310286 363218 320290 363454
rect 320526 363218 330530 363454
rect 330766 363218 340770 363454
rect 341006 363218 351010 363454
rect 351246 363218 361250 363454
rect 361486 363218 371490 363454
rect 371726 363218 381730 363454
rect 381966 363218 391970 363454
rect 392206 363218 402210 363454
rect 402446 363218 412450 363454
rect 412686 363218 422690 363454
rect 422926 363218 432930 363454
rect 433166 363218 443170 363454
rect 443406 363218 453410 363454
rect 453646 363218 463650 363454
rect 463886 363218 473890 363454
rect 474126 363218 484130 363454
rect 484366 363218 494370 363454
rect 494606 363218 504610 363454
rect 504846 363218 514850 363454
rect 515086 363218 525090 363454
rect 525326 363218 535330 363454
rect 535566 363218 544546 363454
rect 544782 363218 544866 363454
rect 545102 363218 554786 363454
rect 555022 363218 555106 363454
rect 555342 363218 565026 363454
rect 565262 363218 565346 363454
rect 565582 363218 575266 363454
rect 575502 363218 575586 363454
rect 575822 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 12066 363134
rect 12302 362898 12386 363134
rect 12622 362898 23330 363134
rect 23566 362898 33570 363134
rect 33806 362898 43810 363134
rect 44046 362898 54050 363134
rect 54286 362898 64290 363134
rect 64526 362898 74530 363134
rect 74766 362898 84770 363134
rect 85006 362898 95010 363134
rect 95246 362898 105250 363134
rect 105486 362898 115490 363134
rect 115726 362898 125730 363134
rect 125966 362898 135970 363134
rect 136206 362898 146210 363134
rect 146446 362898 156450 363134
rect 156686 362898 166690 363134
rect 166926 362898 176930 363134
rect 177166 362898 187170 363134
rect 187406 362898 197410 363134
rect 197646 362898 207650 363134
rect 207886 362898 217890 363134
rect 218126 362898 228130 363134
rect 228366 362898 238370 363134
rect 238606 362898 248610 363134
rect 248846 362898 258850 363134
rect 259086 362898 269090 363134
rect 269326 362898 279330 363134
rect 279566 362898 289570 363134
rect 289806 362898 299810 363134
rect 300046 362898 310050 363134
rect 310286 362898 320290 363134
rect 320526 362898 330530 363134
rect 330766 362898 340770 363134
rect 341006 362898 351010 363134
rect 351246 362898 361250 363134
rect 361486 362898 371490 363134
rect 371726 362898 381730 363134
rect 381966 362898 391970 363134
rect 392206 362898 402210 363134
rect 402446 362898 412450 363134
rect 412686 362898 422690 363134
rect 422926 362898 432930 363134
rect 433166 362898 443170 363134
rect 443406 362898 453410 363134
rect 453646 362898 463650 363134
rect 463886 362898 473890 363134
rect 474126 362898 484130 363134
rect 484366 362898 494370 363134
rect 494606 362898 504610 363134
rect 504846 362898 514850 363134
rect 515086 362898 525090 363134
rect 525326 362898 535330 363134
rect 535566 362898 544546 363134
rect 544782 362898 544866 363134
rect 545102 362898 554786 363134
rect 555022 362898 555106 363134
rect 555342 362898 565026 363134
rect 565262 362898 565346 363134
rect 565582 362898 575266 363134
rect 575502 362898 575586 363134
rect 575822 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 550586 356614
rect 550822 356378 550906 356614
rect 551142 356378 560826 356614
rect 561062 356378 561146 356614
rect 561382 356378 571066 356614
rect 571302 356378 571386 356614
rect 571622 356378 581306 356614
rect 581542 356378 581626 356614
rect 581862 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 550586 356294
rect 550822 356058 550906 356294
rect 551142 356058 560826 356294
rect 561062 356058 561146 356294
rect 561382 356058 571066 356294
rect 571302 356058 571386 356294
rect 571622 356058 581306 356294
rect 581542 356058 581626 356294
rect 581862 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 14386 352894
rect 14622 352658 14706 352894
rect 14942 352658 546866 352894
rect 547102 352658 547186 352894
rect 547422 352658 557106 352894
rect 557342 352658 557426 352894
rect 557662 352658 567346 352894
rect 567582 352658 567666 352894
rect 567902 352658 577586 352894
rect 577822 352658 577906 352894
rect 578142 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 14386 352574
rect 14622 352338 14706 352574
rect 14942 352338 546866 352574
rect 547102 352338 547186 352574
rect 547422 352338 557106 352574
rect 557342 352338 557426 352574
rect 557662 352338 567346 352574
rect 567582 352338 567666 352574
rect 567902 352338 577586 352574
rect 577822 352338 577906 352574
rect 578142 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 10666 349174
rect 10902 348938 10986 349174
rect 11222 348938 543146 349174
rect 543382 348938 543466 349174
rect 543702 348938 553386 349174
rect 553622 348938 553706 349174
rect 553942 348938 563626 349174
rect 563862 348938 563946 349174
rect 564182 348938 573866 349174
rect 574102 348938 574186 349174
rect 574422 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 10666 348854
rect 10902 348618 10986 348854
rect 11222 348618 543146 348854
rect 543382 348618 543466 348854
rect 543702 348618 553386 348854
rect 553622 348618 553706 348854
rect 553942 348618 563626 348854
rect 563862 348618 563946 348854
rect 564182 348618 573866 348854
rect 574102 348618 574186 348854
rect 574422 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 6946 345454
rect 7182 345218 7266 345454
rect 7502 345218 28450 345454
rect 28686 345218 38690 345454
rect 38926 345218 48930 345454
rect 49166 345218 59170 345454
rect 59406 345218 69410 345454
rect 69646 345218 79650 345454
rect 79886 345218 89890 345454
rect 90126 345218 100130 345454
rect 100366 345218 110370 345454
rect 110606 345218 120610 345454
rect 120846 345218 130850 345454
rect 131086 345218 141090 345454
rect 141326 345218 151330 345454
rect 151566 345218 161570 345454
rect 161806 345218 171810 345454
rect 172046 345218 182050 345454
rect 182286 345218 192290 345454
rect 192526 345218 202530 345454
rect 202766 345218 212770 345454
rect 213006 345218 223010 345454
rect 223246 345218 233250 345454
rect 233486 345218 243490 345454
rect 243726 345218 253730 345454
rect 253966 345218 263970 345454
rect 264206 345218 274210 345454
rect 274446 345218 284450 345454
rect 284686 345218 294690 345454
rect 294926 345218 304930 345454
rect 305166 345218 315170 345454
rect 315406 345218 325410 345454
rect 325646 345218 335650 345454
rect 335886 345218 345890 345454
rect 346126 345218 356130 345454
rect 356366 345218 366370 345454
rect 366606 345218 376610 345454
rect 376846 345218 386850 345454
rect 387086 345218 397090 345454
rect 397326 345218 407330 345454
rect 407566 345218 417570 345454
rect 417806 345218 427810 345454
rect 428046 345218 438050 345454
rect 438286 345218 448290 345454
rect 448526 345218 458530 345454
rect 458766 345218 468770 345454
rect 469006 345218 479010 345454
rect 479246 345218 489250 345454
rect 489486 345218 499490 345454
rect 499726 345218 509730 345454
rect 509966 345218 519970 345454
rect 520206 345218 530210 345454
rect 530446 345218 549666 345454
rect 549902 345218 549986 345454
rect 550222 345218 559906 345454
rect 560142 345218 560226 345454
rect 560462 345218 570146 345454
rect 570382 345218 570466 345454
rect 570702 345218 580386 345454
rect 580622 345218 580706 345454
rect 580942 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 6946 345134
rect 7182 344898 7266 345134
rect 7502 344898 28450 345134
rect 28686 344898 38690 345134
rect 38926 344898 48930 345134
rect 49166 344898 59170 345134
rect 59406 344898 69410 345134
rect 69646 344898 79650 345134
rect 79886 344898 89890 345134
rect 90126 344898 100130 345134
rect 100366 344898 110370 345134
rect 110606 344898 120610 345134
rect 120846 344898 130850 345134
rect 131086 344898 141090 345134
rect 141326 344898 151330 345134
rect 151566 344898 161570 345134
rect 161806 344898 171810 345134
rect 172046 344898 182050 345134
rect 182286 344898 192290 345134
rect 192526 344898 202530 345134
rect 202766 344898 212770 345134
rect 213006 344898 223010 345134
rect 223246 344898 233250 345134
rect 233486 344898 243490 345134
rect 243726 344898 253730 345134
rect 253966 344898 263970 345134
rect 264206 344898 274210 345134
rect 274446 344898 284450 345134
rect 284686 344898 294690 345134
rect 294926 344898 304930 345134
rect 305166 344898 315170 345134
rect 315406 344898 325410 345134
rect 325646 344898 335650 345134
rect 335886 344898 345890 345134
rect 346126 344898 356130 345134
rect 356366 344898 366370 345134
rect 366606 344898 376610 345134
rect 376846 344898 386850 345134
rect 387086 344898 397090 345134
rect 397326 344898 407330 345134
rect 407566 344898 417570 345134
rect 417806 344898 427810 345134
rect 428046 344898 438050 345134
rect 438286 344898 448290 345134
rect 448526 344898 458530 345134
rect 458766 344898 468770 345134
rect 469006 344898 479010 345134
rect 479246 344898 489250 345134
rect 489486 344898 499490 345134
rect 499726 344898 509730 345134
rect 509966 344898 519970 345134
rect 520206 344898 530210 345134
rect 530446 344898 549666 345134
rect 549902 344898 549986 345134
rect 550222 344898 559906 345134
rect 560142 344898 560226 345134
rect 560462 344898 570146 345134
rect 570382 344898 570466 345134
rect 570702 344898 580386 345134
rect 580622 344898 580706 345134
rect 580942 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 545466 338614
rect 545702 338378 545786 338614
rect 546022 338378 555706 338614
rect 555942 338378 556026 338614
rect 556262 338378 565946 338614
rect 566182 338378 566266 338614
rect 566502 338378 576186 338614
rect 576422 338378 576506 338614
rect 576742 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 545466 338294
rect 545702 338058 545786 338294
rect 546022 338058 555706 338294
rect 555942 338058 556026 338294
rect 556262 338058 565946 338294
rect 566182 338058 566266 338294
rect 566502 338058 576186 338294
rect 576422 338058 576506 338294
rect 576742 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 541746 334894
rect 541982 334658 542066 334894
rect 542302 334658 551986 334894
rect 552222 334658 552306 334894
rect 552542 334658 562226 334894
rect 562462 334658 562546 334894
rect 562782 334658 572466 334894
rect 572702 334658 572786 334894
rect 573022 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 541746 334574
rect 541982 334338 542066 334574
rect 542302 334338 551986 334574
rect 552222 334338 552306 334574
rect 552542 334338 562226 334574
rect 562462 334338 562546 334574
rect 562782 334338 572466 334574
rect 572702 334338 572786 334574
rect 573022 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 15786 331174
rect 16022 330938 16106 331174
rect 16342 330938 548266 331174
rect 548502 330938 548586 331174
rect 548822 330938 558506 331174
rect 558742 330938 558826 331174
rect 559062 330938 568746 331174
rect 568982 330938 569066 331174
rect 569302 330938 578986 331174
rect 579222 330938 579306 331174
rect 579542 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 15786 330854
rect 16022 330618 16106 330854
rect 16342 330618 548266 330854
rect 548502 330618 548586 330854
rect 548822 330618 558506 330854
rect 558742 330618 558826 330854
rect 559062 330618 568746 330854
rect 568982 330618 569066 330854
rect 569302 330618 578986 330854
rect 579222 330618 579306 330854
rect 579542 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 12066 327454
rect 12302 327218 12386 327454
rect 12622 327218 23330 327454
rect 23566 327218 33570 327454
rect 33806 327218 43810 327454
rect 44046 327218 54050 327454
rect 54286 327218 64290 327454
rect 64526 327218 74530 327454
rect 74766 327218 84770 327454
rect 85006 327218 95010 327454
rect 95246 327218 105250 327454
rect 105486 327218 115490 327454
rect 115726 327218 125730 327454
rect 125966 327218 135970 327454
rect 136206 327218 146210 327454
rect 146446 327218 156450 327454
rect 156686 327218 166690 327454
rect 166926 327218 176930 327454
rect 177166 327218 187170 327454
rect 187406 327218 197410 327454
rect 197646 327218 207650 327454
rect 207886 327218 217890 327454
rect 218126 327218 228130 327454
rect 228366 327218 238370 327454
rect 238606 327218 248610 327454
rect 248846 327218 258850 327454
rect 259086 327218 269090 327454
rect 269326 327218 279330 327454
rect 279566 327218 289570 327454
rect 289806 327218 299810 327454
rect 300046 327218 310050 327454
rect 310286 327218 320290 327454
rect 320526 327218 330530 327454
rect 330766 327218 340770 327454
rect 341006 327218 351010 327454
rect 351246 327218 361250 327454
rect 361486 327218 371490 327454
rect 371726 327218 381730 327454
rect 381966 327218 391970 327454
rect 392206 327218 402210 327454
rect 402446 327218 412450 327454
rect 412686 327218 422690 327454
rect 422926 327218 432930 327454
rect 433166 327218 443170 327454
rect 443406 327218 453410 327454
rect 453646 327218 463650 327454
rect 463886 327218 473890 327454
rect 474126 327218 484130 327454
rect 484366 327218 494370 327454
rect 494606 327218 504610 327454
rect 504846 327218 514850 327454
rect 515086 327218 525090 327454
rect 525326 327218 535330 327454
rect 535566 327218 544546 327454
rect 544782 327218 544866 327454
rect 545102 327218 554786 327454
rect 555022 327218 555106 327454
rect 555342 327218 565026 327454
rect 565262 327218 565346 327454
rect 565582 327218 575266 327454
rect 575502 327218 575586 327454
rect 575822 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 12066 327134
rect 12302 326898 12386 327134
rect 12622 326898 23330 327134
rect 23566 326898 33570 327134
rect 33806 326898 43810 327134
rect 44046 326898 54050 327134
rect 54286 326898 64290 327134
rect 64526 326898 74530 327134
rect 74766 326898 84770 327134
rect 85006 326898 95010 327134
rect 95246 326898 105250 327134
rect 105486 326898 115490 327134
rect 115726 326898 125730 327134
rect 125966 326898 135970 327134
rect 136206 326898 146210 327134
rect 146446 326898 156450 327134
rect 156686 326898 166690 327134
rect 166926 326898 176930 327134
rect 177166 326898 187170 327134
rect 187406 326898 197410 327134
rect 197646 326898 207650 327134
rect 207886 326898 217890 327134
rect 218126 326898 228130 327134
rect 228366 326898 238370 327134
rect 238606 326898 248610 327134
rect 248846 326898 258850 327134
rect 259086 326898 269090 327134
rect 269326 326898 279330 327134
rect 279566 326898 289570 327134
rect 289806 326898 299810 327134
rect 300046 326898 310050 327134
rect 310286 326898 320290 327134
rect 320526 326898 330530 327134
rect 330766 326898 340770 327134
rect 341006 326898 351010 327134
rect 351246 326898 361250 327134
rect 361486 326898 371490 327134
rect 371726 326898 381730 327134
rect 381966 326898 391970 327134
rect 392206 326898 402210 327134
rect 402446 326898 412450 327134
rect 412686 326898 422690 327134
rect 422926 326898 432930 327134
rect 433166 326898 443170 327134
rect 443406 326898 453410 327134
rect 453646 326898 463650 327134
rect 463886 326898 473890 327134
rect 474126 326898 484130 327134
rect 484366 326898 494370 327134
rect 494606 326898 504610 327134
rect 504846 326898 514850 327134
rect 515086 326898 525090 327134
rect 525326 326898 535330 327134
rect 535566 326898 544546 327134
rect 544782 326898 544866 327134
rect 545102 326898 554786 327134
rect 555022 326898 555106 327134
rect 555342 326898 565026 327134
rect 565262 326898 565346 327134
rect 565582 326898 575266 327134
rect 575502 326898 575586 327134
rect 575822 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 550586 320614
rect 550822 320378 550906 320614
rect 551142 320378 560826 320614
rect 561062 320378 561146 320614
rect 561382 320378 571066 320614
rect 571302 320378 571386 320614
rect 571622 320378 581306 320614
rect 581542 320378 581626 320614
rect 581862 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 550586 320294
rect 550822 320058 550906 320294
rect 551142 320058 560826 320294
rect 561062 320058 561146 320294
rect 561382 320058 571066 320294
rect 571302 320058 571386 320294
rect 571622 320058 581306 320294
rect 581542 320058 581626 320294
rect 581862 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 14386 316894
rect 14622 316658 14706 316894
rect 14942 316658 546866 316894
rect 547102 316658 547186 316894
rect 547422 316658 557106 316894
rect 557342 316658 557426 316894
rect 557662 316658 567346 316894
rect 567582 316658 567666 316894
rect 567902 316658 577586 316894
rect 577822 316658 577906 316894
rect 578142 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 14386 316574
rect 14622 316338 14706 316574
rect 14942 316338 546866 316574
rect 547102 316338 547186 316574
rect 547422 316338 557106 316574
rect 557342 316338 557426 316574
rect 557662 316338 567346 316574
rect 567582 316338 567666 316574
rect 567902 316338 577586 316574
rect 577822 316338 577906 316574
rect 578142 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 10666 313174
rect 10902 312938 10986 313174
rect 11222 312938 543146 313174
rect 543382 312938 543466 313174
rect 543702 312938 553386 313174
rect 553622 312938 553706 313174
rect 553942 312938 563626 313174
rect 563862 312938 563946 313174
rect 564182 312938 573866 313174
rect 574102 312938 574186 313174
rect 574422 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 10666 312854
rect 10902 312618 10986 312854
rect 11222 312618 543146 312854
rect 543382 312618 543466 312854
rect 543702 312618 553386 312854
rect 553622 312618 553706 312854
rect 553942 312618 563626 312854
rect 563862 312618 563946 312854
rect 564182 312618 573866 312854
rect 574102 312618 574186 312854
rect 574422 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 6946 309454
rect 7182 309218 7266 309454
rect 7502 309218 28450 309454
rect 28686 309218 38690 309454
rect 38926 309218 48930 309454
rect 49166 309218 59170 309454
rect 59406 309218 69410 309454
rect 69646 309218 79650 309454
rect 79886 309218 89890 309454
rect 90126 309218 100130 309454
rect 100366 309218 110370 309454
rect 110606 309218 120610 309454
rect 120846 309218 130850 309454
rect 131086 309218 141090 309454
rect 141326 309218 151330 309454
rect 151566 309218 161570 309454
rect 161806 309218 171810 309454
rect 172046 309218 182050 309454
rect 182286 309218 192290 309454
rect 192526 309218 202530 309454
rect 202766 309218 212770 309454
rect 213006 309218 223010 309454
rect 223246 309218 233250 309454
rect 233486 309218 243490 309454
rect 243726 309218 253730 309454
rect 253966 309218 263970 309454
rect 264206 309218 274210 309454
rect 274446 309218 284450 309454
rect 284686 309218 294690 309454
rect 294926 309218 304930 309454
rect 305166 309218 315170 309454
rect 315406 309218 325410 309454
rect 325646 309218 335650 309454
rect 335886 309218 345890 309454
rect 346126 309218 356130 309454
rect 356366 309218 366370 309454
rect 366606 309218 376610 309454
rect 376846 309218 386850 309454
rect 387086 309218 397090 309454
rect 397326 309218 407330 309454
rect 407566 309218 417570 309454
rect 417806 309218 427810 309454
rect 428046 309218 438050 309454
rect 438286 309218 448290 309454
rect 448526 309218 458530 309454
rect 458766 309218 468770 309454
rect 469006 309218 479010 309454
rect 479246 309218 489250 309454
rect 489486 309218 499490 309454
rect 499726 309218 509730 309454
rect 509966 309218 519970 309454
rect 520206 309218 530210 309454
rect 530446 309218 549666 309454
rect 549902 309218 549986 309454
rect 550222 309218 559906 309454
rect 560142 309218 560226 309454
rect 560462 309218 570146 309454
rect 570382 309218 570466 309454
rect 570702 309218 580386 309454
rect 580622 309218 580706 309454
rect 580942 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 6946 309134
rect 7182 308898 7266 309134
rect 7502 308898 28450 309134
rect 28686 308898 38690 309134
rect 38926 308898 48930 309134
rect 49166 308898 59170 309134
rect 59406 308898 69410 309134
rect 69646 308898 79650 309134
rect 79886 308898 89890 309134
rect 90126 308898 100130 309134
rect 100366 308898 110370 309134
rect 110606 308898 120610 309134
rect 120846 308898 130850 309134
rect 131086 308898 141090 309134
rect 141326 308898 151330 309134
rect 151566 308898 161570 309134
rect 161806 308898 171810 309134
rect 172046 308898 182050 309134
rect 182286 308898 192290 309134
rect 192526 308898 202530 309134
rect 202766 308898 212770 309134
rect 213006 308898 223010 309134
rect 223246 308898 233250 309134
rect 233486 308898 243490 309134
rect 243726 308898 253730 309134
rect 253966 308898 263970 309134
rect 264206 308898 274210 309134
rect 274446 308898 284450 309134
rect 284686 308898 294690 309134
rect 294926 308898 304930 309134
rect 305166 308898 315170 309134
rect 315406 308898 325410 309134
rect 325646 308898 335650 309134
rect 335886 308898 345890 309134
rect 346126 308898 356130 309134
rect 356366 308898 366370 309134
rect 366606 308898 376610 309134
rect 376846 308898 386850 309134
rect 387086 308898 397090 309134
rect 397326 308898 407330 309134
rect 407566 308898 417570 309134
rect 417806 308898 427810 309134
rect 428046 308898 438050 309134
rect 438286 308898 448290 309134
rect 448526 308898 458530 309134
rect 458766 308898 468770 309134
rect 469006 308898 479010 309134
rect 479246 308898 489250 309134
rect 489486 308898 499490 309134
rect 499726 308898 509730 309134
rect 509966 308898 519970 309134
rect 520206 308898 530210 309134
rect 530446 308898 549666 309134
rect 549902 308898 549986 309134
rect 550222 308898 559906 309134
rect 560142 308898 560226 309134
rect 560462 308898 570146 309134
rect 570382 308898 570466 309134
rect 570702 308898 580386 309134
rect 580622 308898 580706 309134
rect 580942 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 545466 302614
rect 545702 302378 545786 302614
rect 546022 302378 555706 302614
rect 555942 302378 556026 302614
rect 556262 302378 565946 302614
rect 566182 302378 566266 302614
rect 566502 302378 576186 302614
rect 576422 302378 576506 302614
rect 576742 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 545466 302294
rect 545702 302058 545786 302294
rect 546022 302058 555706 302294
rect 555942 302058 556026 302294
rect 556262 302058 565946 302294
rect 566182 302058 566266 302294
rect 566502 302058 576186 302294
rect 576422 302058 576506 302294
rect 576742 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 541746 298894
rect 541982 298658 542066 298894
rect 542302 298658 551986 298894
rect 552222 298658 552306 298894
rect 552542 298658 562226 298894
rect 562462 298658 562546 298894
rect 562782 298658 572466 298894
rect 572702 298658 572786 298894
rect 573022 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 541746 298574
rect 541982 298338 542066 298574
rect 542302 298338 551986 298574
rect 552222 298338 552306 298574
rect 552542 298338 562226 298574
rect 562462 298338 562546 298574
rect 562782 298338 572466 298574
rect 572702 298338 572786 298574
rect 573022 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 15786 295174
rect 16022 294938 16106 295174
rect 16342 294938 548266 295174
rect 548502 294938 548586 295174
rect 548822 294938 558506 295174
rect 558742 294938 558826 295174
rect 559062 294938 568746 295174
rect 568982 294938 569066 295174
rect 569302 294938 578986 295174
rect 579222 294938 579306 295174
rect 579542 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 15786 294854
rect 16022 294618 16106 294854
rect 16342 294618 548266 294854
rect 548502 294618 548586 294854
rect 548822 294618 558506 294854
rect 558742 294618 558826 294854
rect 559062 294618 568746 294854
rect 568982 294618 569066 294854
rect 569302 294618 578986 294854
rect 579222 294618 579306 294854
rect 579542 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 12066 291454
rect 12302 291218 12386 291454
rect 12622 291218 23330 291454
rect 23566 291218 33570 291454
rect 33806 291218 43810 291454
rect 44046 291218 54050 291454
rect 54286 291218 64290 291454
rect 64526 291218 74530 291454
rect 74766 291218 84770 291454
rect 85006 291218 95010 291454
rect 95246 291218 105250 291454
rect 105486 291218 115490 291454
rect 115726 291218 125730 291454
rect 125966 291218 135970 291454
rect 136206 291218 146210 291454
rect 146446 291218 156450 291454
rect 156686 291218 166690 291454
rect 166926 291218 176930 291454
rect 177166 291218 187170 291454
rect 187406 291218 197410 291454
rect 197646 291218 207650 291454
rect 207886 291218 217890 291454
rect 218126 291218 228130 291454
rect 228366 291218 238370 291454
rect 238606 291218 248610 291454
rect 248846 291218 258850 291454
rect 259086 291218 269090 291454
rect 269326 291218 279330 291454
rect 279566 291218 289570 291454
rect 289806 291218 299810 291454
rect 300046 291218 310050 291454
rect 310286 291218 320290 291454
rect 320526 291218 330530 291454
rect 330766 291218 340770 291454
rect 341006 291218 351010 291454
rect 351246 291218 361250 291454
rect 361486 291218 371490 291454
rect 371726 291218 381730 291454
rect 381966 291218 391970 291454
rect 392206 291218 402210 291454
rect 402446 291218 412450 291454
rect 412686 291218 422690 291454
rect 422926 291218 432930 291454
rect 433166 291218 443170 291454
rect 443406 291218 453410 291454
rect 453646 291218 463650 291454
rect 463886 291218 473890 291454
rect 474126 291218 484130 291454
rect 484366 291218 494370 291454
rect 494606 291218 504610 291454
rect 504846 291218 514850 291454
rect 515086 291218 525090 291454
rect 525326 291218 535330 291454
rect 535566 291218 544546 291454
rect 544782 291218 544866 291454
rect 545102 291218 554786 291454
rect 555022 291218 555106 291454
rect 555342 291218 565026 291454
rect 565262 291218 565346 291454
rect 565582 291218 575266 291454
rect 575502 291218 575586 291454
rect 575822 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 12066 291134
rect 12302 290898 12386 291134
rect 12622 290898 23330 291134
rect 23566 290898 33570 291134
rect 33806 290898 43810 291134
rect 44046 290898 54050 291134
rect 54286 290898 64290 291134
rect 64526 290898 74530 291134
rect 74766 290898 84770 291134
rect 85006 290898 95010 291134
rect 95246 290898 105250 291134
rect 105486 290898 115490 291134
rect 115726 290898 125730 291134
rect 125966 290898 135970 291134
rect 136206 290898 146210 291134
rect 146446 290898 156450 291134
rect 156686 290898 166690 291134
rect 166926 290898 176930 291134
rect 177166 290898 187170 291134
rect 187406 290898 197410 291134
rect 197646 290898 207650 291134
rect 207886 290898 217890 291134
rect 218126 290898 228130 291134
rect 228366 290898 238370 291134
rect 238606 290898 248610 291134
rect 248846 290898 258850 291134
rect 259086 290898 269090 291134
rect 269326 290898 279330 291134
rect 279566 290898 289570 291134
rect 289806 290898 299810 291134
rect 300046 290898 310050 291134
rect 310286 290898 320290 291134
rect 320526 290898 330530 291134
rect 330766 290898 340770 291134
rect 341006 290898 351010 291134
rect 351246 290898 361250 291134
rect 361486 290898 371490 291134
rect 371726 290898 381730 291134
rect 381966 290898 391970 291134
rect 392206 290898 402210 291134
rect 402446 290898 412450 291134
rect 412686 290898 422690 291134
rect 422926 290898 432930 291134
rect 433166 290898 443170 291134
rect 443406 290898 453410 291134
rect 453646 290898 463650 291134
rect 463886 290898 473890 291134
rect 474126 290898 484130 291134
rect 484366 290898 494370 291134
rect 494606 290898 504610 291134
rect 504846 290898 514850 291134
rect 515086 290898 525090 291134
rect 525326 290898 535330 291134
rect 535566 290898 544546 291134
rect 544782 290898 544866 291134
rect 545102 290898 554786 291134
rect 555022 290898 555106 291134
rect 555342 290898 565026 291134
rect 565262 290898 565346 291134
rect 565582 290898 575266 291134
rect 575502 290898 575586 291134
rect 575822 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 550586 284614
rect 550822 284378 550906 284614
rect 551142 284378 560826 284614
rect 561062 284378 561146 284614
rect 561382 284378 571066 284614
rect 571302 284378 571386 284614
rect 571622 284378 581306 284614
rect 581542 284378 581626 284614
rect 581862 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 550586 284294
rect 550822 284058 550906 284294
rect 551142 284058 560826 284294
rect 561062 284058 561146 284294
rect 561382 284058 571066 284294
rect 571302 284058 571386 284294
rect 571622 284058 581306 284294
rect 581542 284058 581626 284294
rect 581862 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 14386 280894
rect 14622 280658 14706 280894
rect 14942 280658 546866 280894
rect 547102 280658 547186 280894
rect 547422 280658 557106 280894
rect 557342 280658 557426 280894
rect 557662 280658 567346 280894
rect 567582 280658 567666 280894
rect 567902 280658 577586 280894
rect 577822 280658 577906 280894
rect 578142 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 14386 280574
rect 14622 280338 14706 280574
rect 14942 280338 546866 280574
rect 547102 280338 547186 280574
rect 547422 280338 557106 280574
rect 557342 280338 557426 280574
rect 557662 280338 567346 280574
rect 567582 280338 567666 280574
rect 567902 280338 577586 280574
rect 577822 280338 577906 280574
rect 578142 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 10666 277174
rect 10902 276938 10986 277174
rect 11222 276938 543146 277174
rect 543382 276938 543466 277174
rect 543702 276938 553386 277174
rect 553622 276938 553706 277174
rect 553942 276938 563626 277174
rect 563862 276938 563946 277174
rect 564182 276938 573866 277174
rect 574102 276938 574186 277174
rect 574422 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 10666 276854
rect 10902 276618 10986 276854
rect 11222 276618 543146 276854
rect 543382 276618 543466 276854
rect 543702 276618 553386 276854
rect 553622 276618 553706 276854
rect 553942 276618 563626 276854
rect 563862 276618 563946 276854
rect 564182 276618 573866 276854
rect 574102 276618 574186 276854
rect 574422 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 6946 273454
rect 7182 273218 7266 273454
rect 7502 273218 28450 273454
rect 28686 273218 38690 273454
rect 38926 273218 48930 273454
rect 49166 273218 59170 273454
rect 59406 273218 69410 273454
rect 69646 273218 79650 273454
rect 79886 273218 89890 273454
rect 90126 273218 100130 273454
rect 100366 273218 110370 273454
rect 110606 273218 120610 273454
rect 120846 273218 130850 273454
rect 131086 273218 141090 273454
rect 141326 273218 151330 273454
rect 151566 273218 161570 273454
rect 161806 273218 171810 273454
rect 172046 273218 182050 273454
rect 182286 273218 192290 273454
rect 192526 273218 202530 273454
rect 202766 273218 212770 273454
rect 213006 273218 223010 273454
rect 223246 273218 233250 273454
rect 233486 273218 243490 273454
rect 243726 273218 253730 273454
rect 253966 273218 263970 273454
rect 264206 273218 274210 273454
rect 274446 273218 284450 273454
rect 284686 273218 294690 273454
rect 294926 273218 304930 273454
rect 305166 273218 315170 273454
rect 315406 273218 325410 273454
rect 325646 273218 335650 273454
rect 335886 273218 345890 273454
rect 346126 273218 356130 273454
rect 356366 273218 366370 273454
rect 366606 273218 376610 273454
rect 376846 273218 386850 273454
rect 387086 273218 397090 273454
rect 397326 273218 407330 273454
rect 407566 273218 417570 273454
rect 417806 273218 427810 273454
rect 428046 273218 438050 273454
rect 438286 273218 448290 273454
rect 448526 273218 458530 273454
rect 458766 273218 468770 273454
rect 469006 273218 479010 273454
rect 479246 273218 489250 273454
rect 489486 273218 499490 273454
rect 499726 273218 509730 273454
rect 509966 273218 519970 273454
rect 520206 273218 530210 273454
rect 530446 273218 549666 273454
rect 549902 273218 549986 273454
rect 550222 273218 559906 273454
rect 560142 273218 560226 273454
rect 560462 273218 570146 273454
rect 570382 273218 570466 273454
rect 570702 273218 580386 273454
rect 580622 273218 580706 273454
rect 580942 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 6946 273134
rect 7182 272898 7266 273134
rect 7502 272898 28450 273134
rect 28686 272898 38690 273134
rect 38926 272898 48930 273134
rect 49166 272898 59170 273134
rect 59406 272898 69410 273134
rect 69646 272898 79650 273134
rect 79886 272898 89890 273134
rect 90126 272898 100130 273134
rect 100366 272898 110370 273134
rect 110606 272898 120610 273134
rect 120846 272898 130850 273134
rect 131086 272898 141090 273134
rect 141326 272898 151330 273134
rect 151566 272898 161570 273134
rect 161806 272898 171810 273134
rect 172046 272898 182050 273134
rect 182286 272898 192290 273134
rect 192526 272898 202530 273134
rect 202766 272898 212770 273134
rect 213006 272898 223010 273134
rect 223246 272898 233250 273134
rect 233486 272898 243490 273134
rect 243726 272898 253730 273134
rect 253966 272898 263970 273134
rect 264206 272898 274210 273134
rect 274446 272898 284450 273134
rect 284686 272898 294690 273134
rect 294926 272898 304930 273134
rect 305166 272898 315170 273134
rect 315406 272898 325410 273134
rect 325646 272898 335650 273134
rect 335886 272898 345890 273134
rect 346126 272898 356130 273134
rect 356366 272898 366370 273134
rect 366606 272898 376610 273134
rect 376846 272898 386850 273134
rect 387086 272898 397090 273134
rect 397326 272898 407330 273134
rect 407566 272898 417570 273134
rect 417806 272898 427810 273134
rect 428046 272898 438050 273134
rect 438286 272898 448290 273134
rect 448526 272898 458530 273134
rect 458766 272898 468770 273134
rect 469006 272898 479010 273134
rect 479246 272898 489250 273134
rect 489486 272898 499490 273134
rect 499726 272898 509730 273134
rect 509966 272898 519970 273134
rect 520206 272898 530210 273134
rect 530446 272898 549666 273134
rect 549902 272898 549986 273134
rect 550222 272898 559906 273134
rect 560142 272898 560226 273134
rect 560462 272898 570146 273134
rect 570382 272898 570466 273134
rect 570702 272898 580386 273134
rect 580622 272898 580706 273134
rect 580942 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 545466 266614
rect 545702 266378 545786 266614
rect 546022 266378 555706 266614
rect 555942 266378 556026 266614
rect 556262 266378 565946 266614
rect 566182 266378 566266 266614
rect 566502 266378 576186 266614
rect 576422 266378 576506 266614
rect 576742 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 545466 266294
rect 545702 266058 545786 266294
rect 546022 266058 555706 266294
rect 555942 266058 556026 266294
rect 556262 266058 565946 266294
rect 566182 266058 566266 266294
rect 566502 266058 576186 266294
rect 576422 266058 576506 266294
rect 576742 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 541746 262894
rect 541982 262658 542066 262894
rect 542302 262658 551986 262894
rect 552222 262658 552306 262894
rect 552542 262658 562226 262894
rect 562462 262658 562546 262894
rect 562782 262658 572466 262894
rect 572702 262658 572786 262894
rect 573022 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 541746 262574
rect 541982 262338 542066 262574
rect 542302 262338 551986 262574
rect 552222 262338 552306 262574
rect 552542 262338 562226 262574
rect 562462 262338 562546 262574
rect 562782 262338 572466 262574
rect 572702 262338 572786 262574
rect 573022 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 15786 259174
rect 16022 258938 16106 259174
rect 16342 258938 548266 259174
rect 548502 258938 548586 259174
rect 548822 258938 558506 259174
rect 558742 258938 558826 259174
rect 559062 258938 568746 259174
rect 568982 258938 569066 259174
rect 569302 258938 578986 259174
rect 579222 258938 579306 259174
rect 579542 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 15786 258854
rect 16022 258618 16106 258854
rect 16342 258618 548266 258854
rect 548502 258618 548586 258854
rect 548822 258618 558506 258854
rect 558742 258618 558826 258854
rect 559062 258618 568746 258854
rect 568982 258618 569066 258854
rect 569302 258618 578986 258854
rect 579222 258618 579306 258854
rect 579542 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 12066 255454
rect 12302 255218 12386 255454
rect 12622 255218 23330 255454
rect 23566 255218 33570 255454
rect 33806 255218 43810 255454
rect 44046 255218 54050 255454
rect 54286 255218 64290 255454
rect 64526 255218 74530 255454
rect 74766 255218 84770 255454
rect 85006 255218 95010 255454
rect 95246 255218 105250 255454
rect 105486 255218 115490 255454
rect 115726 255218 125730 255454
rect 125966 255218 135970 255454
rect 136206 255218 146210 255454
rect 146446 255218 156450 255454
rect 156686 255218 166690 255454
rect 166926 255218 176930 255454
rect 177166 255218 187170 255454
rect 187406 255218 197410 255454
rect 197646 255218 207650 255454
rect 207886 255218 217890 255454
rect 218126 255218 228130 255454
rect 228366 255218 238370 255454
rect 238606 255218 248610 255454
rect 248846 255218 258850 255454
rect 259086 255218 269090 255454
rect 269326 255218 279330 255454
rect 279566 255218 289570 255454
rect 289806 255218 299810 255454
rect 300046 255218 310050 255454
rect 310286 255218 320290 255454
rect 320526 255218 330530 255454
rect 330766 255218 340770 255454
rect 341006 255218 351010 255454
rect 351246 255218 361250 255454
rect 361486 255218 371490 255454
rect 371726 255218 381730 255454
rect 381966 255218 391970 255454
rect 392206 255218 402210 255454
rect 402446 255218 412450 255454
rect 412686 255218 422690 255454
rect 422926 255218 432930 255454
rect 433166 255218 443170 255454
rect 443406 255218 453410 255454
rect 453646 255218 463650 255454
rect 463886 255218 473890 255454
rect 474126 255218 484130 255454
rect 484366 255218 494370 255454
rect 494606 255218 504610 255454
rect 504846 255218 514850 255454
rect 515086 255218 525090 255454
rect 525326 255218 535330 255454
rect 535566 255218 544546 255454
rect 544782 255218 544866 255454
rect 545102 255218 554786 255454
rect 555022 255218 555106 255454
rect 555342 255218 565026 255454
rect 565262 255218 565346 255454
rect 565582 255218 575266 255454
rect 575502 255218 575586 255454
rect 575822 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 12066 255134
rect 12302 254898 12386 255134
rect 12622 254898 23330 255134
rect 23566 254898 33570 255134
rect 33806 254898 43810 255134
rect 44046 254898 54050 255134
rect 54286 254898 64290 255134
rect 64526 254898 74530 255134
rect 74766 254898 84770 255134
rect 85006 254898 95010 255134
rect 95246 254898 105250 255134
rect 105486 254898 115490 255134
rect 115726 254898 125730 255134
rect 125966 254898 135970 255134
rect 136206 254898 146210 255134
rect 146446 254898 156450 255134
rect 156686 254898 166690 255134
rect 166926 254898 176930 255134
rect 177166 254898 187170 255134
rect 187406 254898 197410 255134
rect 197646 254898 207650 255134
rect 207886 254898 217890 255134
rect 218126 254898 228130 255134
rect 228366 254898 238370 255134
rect 238606 254898 248610 255134
rect 248846 254898 258850 255134
rect 259086 254898 269090 255134
rect 269326 254898 279330 255134
rect 279566 254898 289570 255134
rect 289806 254898 299810 255134
rect 300046 254898 310050 255134
rect 310286 254898 320290 255134
rect 320526 254898 330530 255134
rect 330766 254898 340770 255134
rect 341006 254898 351010 255134
rect 351246 254898 361250 255134
rect 361486 254898 371490 255134
rect 371726 254898 381730 255134
rect 381966 254898 391970 255134
rect 392206 254898 402210 255134
rect 402446 254898 412450 255134
rect 412686 254898 422690 255134
rect 422926 254898 432930 255134
rect 433166 254898 443170 255134
rect 443406 254898 453410 255134
rect 453646 254898 463650 255134
rect 463886 254898 473890 255134
rect 474126 254898 484130 255134
rect 484366 254898 494370 255134
rect 494606 254898 504610 255134
rect 504846 254898 514850 255134
rect 515086 254898 525090 255134
rect 525326 254898 535330 255134
rect 535566 254898 544546 255134
rect 544782 254898 544866 255134
rect 545102 254898 554786 255134
rect 555022 254898 555106 255134
rect 555342 254898 565026 255134
rect 565262 254898 565346 255134
rect 565582 254898 575266 255134
rect 575502 254898 575586 255134
rect 575822 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 550586 248614
rect 550822 248378 550906 248614
rect 551142 248378 560826 248614
rect 561062 248378 561146 248614
rect 561382 248378 571066 248614
rect 571302 248378 571386 248614
rect 571622 248378 581306 248614
rect 581542 248378 581626 248614
rect 581862 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 550586 248294
rect 550822 248058 550906 248294
rect 551142 248058 560826 248294
rect 561062 248058 561146 248294
rect 561382 248058 571066 248294
rect 571302 248058 571386 248294
rect 571622 248058 581306 248294
rect 581542 248058 581626 248294
rect 581862 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 14386 244894
rect 14622 244658 14706 244894
rect 14942 244658 546866 244894
rect 547102 244658 547186 244894
rect 547422 244658 557106 244894
rect 557342 244658 557426 244894
rect 557662 244658 567346 244894
rect 567582 244658 567666 244894
rect 567902 244658 577586 244894
rect 577822 244658 577906 244894
rect 578142 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 14386 244574
rect 14622 244338 14706 244574
rect 14942 244338 546866 244574
rect 547102 244338 547186 244574
rect 547422 244338 557106 244574
rect 557342 244338 557426 244574
rect 557662 244338 567346 244574
rect 567582 244338 567666 244574
rect 567902 244338 577586 244574
rect 577822 244338 577906 244574
rect 578142 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 10666 241174
rect 10902 240938 10986 241174
rect 11222 240938 543146 241174
rect 543382 240938 543466 241174
rect 543702 240938 553386 241174
rect 553622 240938 553706 241174
rect 553942 240938 563626 241174
rect 563862 240938 563946 241174
rect 564182 240938 573866 241174
rect 574102 240938 574186 241174
rect 574422 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 10666 240854
rect 10902 240618 10986 240854
rect 11222 240618 543146 240854
rect 543382 240618 543466 240854
rect 543702 240618 553386 240854
rect 553622 240618 553706 240854
rect 553942 240618 563626 240854
rect 563862 240618 563946 240854
rect 564182 240618 573866 240854
rect 574102 240618 574186 240854
rect 574422 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 6946 237454
rect 7182 237218 7266 237454
rect 7502 237218 28450 237454
rect 28686 237218 38690 237454
rect 38926 237218 48930 237454
rect 49166 237218 59170 237454
rect 59406 237218 69410 237454
rect 69646 237218 79650 237454
rect 79886 237218 89890 237454
rect 90126 237218 100130 237454
rect 100366 237218 110370 237454
rect 110606 237218 120610 237454
rect 120846 237218 130850 237454
rect 131086 237218 141090 237454
rect 141326 237218 151330 237454
rect 151566 237218 161570 237454
rect 161806 237218 171810 237454
rect 172046 237218 182050 237454
rect 182286 237218 192290 237454
rect 192526 237218 202530 237454
rect 202766 237218 212770 237454
rect 213006 237218 223010 237454
rect 223246 237218 233250 237454
rect 233486 237218 243490 237454
rect 243726 237218 253730 237454
rect 253966 237218 263970 237454
rect 264206 237218 274210 237454
rect 274446 237218 284450 237454
rect 284686 237218 294690 237454
rect 294926 237218 304930 237454
rect 305166 237218 315170 237454
rect 315406 237218 325410 237454
rect 325646 237218 335650 237454
rect 335886 237218 345890 237454
rect 346126 237218 356130 237454
rect 356366 237218 366370 237454
rect 366606 237218 376610 237454
rect 376846 237218 386850 237454
rect 387086 237218 397090 237454
rect 397326 237218 407330 237454
rect 407566 237218 417570 237454
rect 417806 237218 427810 237454
rect 428046 237218 438050 237454
rect 438286 237218 448290 237454
rect 448526 237218 458530 237454
rect 458766 237218 468770 237454
rect 469006 237218 479010 237454
rect 479246 237218 489250 237454
rect 489486 237218 499490 237454
rect 499726 237218 509730 237454
rect 509966 237218 519970 237454
rect 520206 237218 530210 237454
rect 530446 237218 549666 237454
rect 549902 237218 549986 237454
rect 550222 237218 559906 237454
rect 560142 237218 560226 237454
rect 560462 237218 570146 237454
rect 570382 237218 570466 237454
rect 570702 237218 580386 237454
rect 580622 237218 580706 237454
rect 580942 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 6946 237134
rect 7182 236898 7266 237134
rect 7502 236898 28450 237134
rect 28686 236898 38690 237134
rect 38926 236898 48930 237134
rect 49166 236898 59170 237134
rect 59406 236898 69410 237134
rect 69646 236898 79650 237134
rect 79886 236898 89890 237134
rect 90126 236898 100130 237134
rect 100366 236898 110370 237134
rect 110606 236898 120610 237134
rect 120846 236898 130850 237134
rect 131086 236898 141090 237134
rect 141326 236898 151330 237134
rect 151566 236898 161570 237134
rect 161806 236898 171810 237134
rect 172046 236898 182050 237134
rect 182286 236898 192290 237134
rect 192526 236898 202530 237134
rect 202766 236898 212770 237134
rect 213006 236898 223010 237134
rect 223246 236898 233250 237134
rect 233486 236898 243490 237134
rect 243726 236898 253730 237134
rect 253966 236898 263970 237134
rect 264206 236898 274210 237134
rect 274446 236898 284450 237134
rect 284686 236898 294690 237134
rect 294926 236898 304930 237134
rect 305166 236898 315170 237134
rect 315406 236898 325410 237134
rect 325646 236898 335650 237134
rect 335886 236898 345890 237134
rect 346126 236898 356130 237134
rect 356366 236898 366370 237134
rect 366606 236898 376610 237134
rect 376846 236898 386850 237134
rect 387086 236898 397090 237134
rect 397326 236898 407330 237134
rect 407566 236898 417570 237134
rect 417806 236898 427810 237134
rect 428046 236898 438050 237134
rect 438286 236898 448290 237134
rect 448526 236898 458530 237134
rect 458766 236898 468770 237134
rect 469006 236898 479010 237134
rect 479246 236898 489250 237134
rect 489486 236898 499490 237134
rect 499726 236898 509730 237134
rect 509966 236898 519970 237134
rect 520206 236898 530210 237134
rect 530446 236898 549666 237134
rect 549902 236898 549986 237134
rect 550222 236898 559906 237134
rect 560142 236898 560226 237134
rect 560462 236898 570146 237134
rect 570382 236898 570466 237134
rect 570702 236898 580386 237134
rect 580622 236898 580706 237134
rect 580942 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 545466 230614
rect 545702 230378 545786 230614
rect 546022 230378 555706 230614
rect 555942 230378 556026 230614
rect 556262 230378 565946 230614
rect 566182 230378 566266 230614
rect 566502 230378 576186 230614
rect 576422 230378 576506 230614
rect 576742 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 545466 230294
rect 545702 230058 545786 230294
rect 546022 230058 555706 230294
rect 555942 230058 556026 230294
rect 556262 230058 565946 230294
rect 566182 230058 566266 230294
rect 566502 230058 576186 230294
rect 576422 230058 576506 230294
rect 576742 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 541746 226894
rect 541982 226658 542066 226894
rect 542302 226658 551986 226894
rect 552222 226658 552306 226894
rect 552542 226658 562226 226894
rect 562462 226658 562546 226894
rect 562782 226658 572466 226894
rect 572702 226658 572786 226894
rect 573022 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 541746 226574
rect 541982 226338 542066 226574
rect 542302 226338 551986 226574
rect 552222 226338 552306 226574
rect 552542 226338 562226 226574
rect 562462 226338 562546 226574
rect 562782 226338 572466 226574
rect 572702 226338 572786 226574
rect 573022 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 15786 223174
rect 16022 222938 16106 223174
rect 16342 222938 548266 223174
rect 548502 222938 548586 223174
rect 548822 222938 558506 223174
rect 558742 222938 558826 223174
rect 559062 222938 568746 223174
rect 568982 222938 569066 223174
rect 569302 222938 578986 223174
rect 579222 222938 579306 223174
rect 579542 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 15786 222854
rect 16022 222618 16106 222854
rect 16342 222618 548266 222854
rect 548502 222618 548586 222854
rect 548822 222618 558506 222854
rect 558742 222618 558826 222854
rect 559062 222618 568746 222854
rect 568982 222618 569066 222854
rect 569302 222618 578986 222854
rect 579222 222618 579306 222854
rect 579542 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 12066 219454
rect 12302 219218 12386 219454
rect 12622 219218 23330 219454
rect 23566 219218 33570 219454
rect 33806 219218 43810 219454
rect 44046 219218 54050 219454
rect 54286 219218 64290 219454
rect 64526 219218 74530 219454
rect 74766 219218 84770 219454
rect 85006 219218 95010 219454
rect 95246 219218 105250 219454
rect 105486 219218 115490 219454
rect 115726 219218 125730 219454
rect 125966 219218 135970 219454
rect 136206 219218 146210 219454
rect 146446 219218 156450 219454
rect 156686 219218 166690 219454
rect 166926 219218 176930 219454
rect 177166 219218 187170 219454
rect 187406 219218 197410 219454
rect 197646 219218 207650 219454
rect 207886 219218 217890 219454
rect 218126 219218 228130 219454
rect 228366 219218 238370 219454
rect 238606 219218 248610 219454
rect 248846 219218 258850 219454
rect 259086 219218 269090 219454
rect 269326 219218 279330 219454
rect 279566 219218 289570 219454
rect 289806 219218 299810 219454
rect 300046 219218 310050 219454
rect 310286 219218 320290 219454
rect 320526 219218 330530 219454
rect 330766 219218 340770 219454
rect 341006 219218 351010 219454
rect 351246 219218 361250 219454
rect 361486 219218 371490 219454
rect 371726 219218 381730 219454
rect 381966 219218 391970 219454
rect 392206 219218 402210 219454
rect 402446 219218 412450 219454
rect 412686 219218 422690 219454
rect 422926 219218 432930 219454
rect 433166 219218 443170 219454
rect 443406 219218 453410 219454
rect 453646 219218 463650 219454
rect 463886 219218 473890 219454
rect 474126 219218 484130 219454
rect 484366 219218 494370 219454
rect 494606 219218 504610 219454
rect 504846 219218 514850 219454
rect 515086 219218 525090 219454
rect 525326 219218 535330 219454
rect 535566 219218 544546 219454
rect 544782 219218 544866 219454
rect 545102 219218 554786 219454
rect 555022 219218 555106 219454
rect 555342 219218 565026 219454
rect 565262 219218 565346 219454
rect 565582 219218 575266 219454
rect 575502 219218 575586 219454
rect 575822 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 12066 219134
rect 12302 218898 12386 219134
rect 12622 218898 23330 219134
rect 23566 218898 33570 219134
rect 33806 218898 43810 219134
rect 44046 218898 54050 219134
rect 54286 218898 64290 219134
rect 64526 218898 74530 219134
rect 74766 218898 84770 219134
rect 85006 218898 95010 219134
rect 95246 218898 105250 219134
rect 105486 218898 115490 219134
rect 115726 218898 125730 219134
rect 125966 218898 135970 219134
rect 136206 218898 146210 219134
rect 146446 218898 156450 219134
rect 156686 218898 166690 219134
rect 166926 218898 176930 219134
rect 177166 218898 187170 219134
rect 187406 218898 197410 219134
rect 197646 218898 207650 219134
rect 207886 218898 217890 219134
rect 218126 218898 228130 219134
rect 228366 218898 238370 219134
rect 238606 218898 248610 219134
rect 248846 218898 258850 219134
rect 259086 218898 269090 219134
rect 269326 218898 279330 219134
rect 279566 218898 289570 219134
rect 289806 218898 299810 219134
rect 300046 218898 310050 219134
rect 310286 218898 320290 219134
rect 320526 218898 330530 219134
rect 330766 218898 340770 219134
rect 341006 218898 351010 219134
rect 351246 218898 361250 219134
rect 361486 218898 371490 219134
rect 371726 218898 381730 219134
rect 381966 218898 391970 219134
rect 392206 218898 402210 219134
rect 402446 218898 412450 219134
rect 412686 218898 422690 219134
rect 422926 218898 432930 219134
rect 433166 218898 443170 219134
rect 443406 218898 453410 219134
rect 453646 218898 463650 219134
rect 463886 218898 473890 219134
rect 474126 218898 484130 219134
rect 484366 218898 494370 219134
rect 494606 218898 504610 219134
rect 504846 218898 514850 219134
rect 515086 218898 525090 219134
rect 525326 218898 535330 219134
rect 535566 218898 544546 219134
rect 544782 218898 544866 219134
rect 545102 218898 554786 219134
rect 555022 218898 555106 219134
rect 555342 218898 565026 219134
rect 565262 218898 565346 219134
rect 565582 218898 575266 219134
rect 575502 218898 575586 219134
rect 575822 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 550586 212614
rect 550822 212378 550906 212614
rect 551142 212378 560826 212614
rect 561062 212378 561146 212614
rect 561382 212378 571066 212614
rect 571302 212378 571386 212614
rect 571622 212378 581306 212614
rect 581542 212378 581626 212614
rect 581862 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 550586 212294
rect 550822 212058 550906 212294
rect 551142 212058 560826 212294
rect 561062 212058 561146 212294
rect 561382 212058 571066 212294
rect 571302 212058 571386 212294
rect 571622 212058 581306 212294
rect 581542 212058 581626 212294
rect 581862 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 14386 208894
rect 14622 208658 14706 208894
rect 14942 208658 546866 208894
rect 547102 208658 547186 208894
rect 547422 208658 557106 208894
rect 557342 208658 557426 208894
rect 557662 208658 567346 208894
rect 567582 208658 567666 208894
rect 567902 208658 577586 208894
rect 577822 208658 577906 208894
rect 578142 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 14386 208574
rect 14622 208338 14706 208574
rect 14942 208338 546866 208574
rect 547102 208338 547186 208574
rect 547422 208338 557106 208574
rect 557342 208338 557426 208574
rect 557662 208338 567346 208574
rect 567582 208338 567666 208574
rect 567902 208338 577586 208574
rect 577822 208338 577906 208574
rect 578142 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 10666 205174
rect 10902 204938 10986 205174
rect 11222 204938 543146 205174
rect 543382 204938 543466 205174
rect 543702 204938 553386 205174
rect 553622 204938 553706 205174
rect 553942 204938 563626 205174
rect 563862 204938 563946 205174
rect 564182 204938 573866 205174
rect 574102 204938 574186 205174
rect 574422 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 10666 204854
rect 10902 204618 10986 204854
rect 11222 204618 543146 204854
rect 543382 204618 543466 204854
rect 543702 204618 553386 204854
rect 553622 204618 553706 204854
rect 553942 204618 563626 204854
rect 563862 204618 563946 204854
rect 564182 204618 573866 204854
rect 574102 204618 574186 204854
rect 574422 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 6946 201454
rect 7182 201218 7266 201454
rect 7502 201218 28450 201454
rect 28686 201218 38690 201454
rect 38926 201218 48930 201454
rect 49166 201218 59170 201454
rect 59406 201218 69410 201454
rect 69646 201218 79650 201454
rect 79886 201218 89890 201454
rect 90126 201218 100130 201454
rect 100366 201218 110370 201454
rect 110606 201218 120610 201454
rect 120846 201218 130850 201454
rect 131086 201218 141090 201454
rect 141326 201218 151330 201454
rect 151566 201218 161570 201454
rect 161806 201218 171810 201454
rect 172046 201218 182050 201454
rect 182286 201218 192290 201454
rect 192526 201218 202530 201454
rect 202766 201218 212770 201454
rect 213006 201218 223010 201454
rect 223246 201218 233250 201454
rect 233486 201218 243490 201454
rect 243726 201218 253730 201454
rect 253966 201218 263970 201454
rect 264206 201218 274210 201454
rect 274446 201218 284450 201454
rect 284686 201218 294690 201454
rect 294926 201218 304930 201454
rect 305166 201218 315170 201454
rect 315406 201218 325410 201454
rect 325646 201218 335650 201454
rect 335886 201218 345890 201454
rect 346126 201218 356130 201454
rect 356366 201218 366370 201454
rect 366606 201218 376610 201454
rect 376846 201218 386850 201454
rect 387086 201218 397090 201454
rect 397326 201218 407330 201454
rect 407566 201218 417570 201454
rect 417806 201218 427810 201454
rect 428046 201218 438050 201454
rect 438286 201218 448290 201454
rect 448526 201218 458530 201454
rect 458766 201218 468770 201454
rect 469006 201218 479010 201454
rect 479246 201218 489250 201454
rect 489486 201218 499490 201454
rect 499726 201218 509730 201454
rect 509966 201218 519970 201454
rect 520206 201218 530210 201454
rect 530446 201218 549666 201454
rect 549902 201218 549986 201454
rect 550222 201218 559906 201454
rect 560142 201218 560226 201454
rect 560462 201218 570146 201454
rect 570382 201218 570466 201454
rect 570702 201218 580386 201454
rect 580622 201218 580706 201454
rect 580942 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 6946 201134
rect 7182 200898 7266 201134
rect 7502 200898 28450 201134
rect 28686 200898 38690 201134
rect 38926 200898 48930 201134
rect 49166 200898 59170 201134
rect 59406 200898 69410 201134
rect 69646 200898 79650 201134
rect 79886 200898 89890 201134
rect 90126 200898 100130 201134
rect 100366 200898 110370 201134
rect 110606 200898 120610 201134
rect 120846 200898 130850 201134
rect 131086 200898 141090 201134
rect 141326 200898 151330 201134
rect 151566 200898 161570 201134
rect 161806 200898 171810 201134
rect 172046 200898 182050 201134
rect 182286 200898 192290 201134
rect 192526 200898 202530 201134
rect 202766 200898 212770 201134
rect 213006 200898 223010 201134
rect 223246 200898 233250 201134
rect 233486 200898 243490 201134
rect 243726 200898 253730 201134
rect 253966 200898 263970 201134
rect 264206 200898 274210 201134
rect 274446 200898 284450 201134
rect 284686 200898 294690 201134
rect 294926 200898 304930 201134
rect 305166 200898 315170 201134
rect 315406 200898 325410 201134
rect 325646 200898 335650 201134
rect 335886 200898 345890 201134
rect 346126 200898 356130 201134
rect 356366 200898 366370 201134
rect 366606 200898 376610 201134
rect 376846 200898 386850 201134
rect 387086 200898 397090 201134
rect 397326 200898 407330 201134
rect 407566 200898 417570 201134
rect 417806 200898 427810 201134
rect 428046 200898 438050 201134
rect 438286 200898 448290 201134
rect 448526 200898 458530 201134
rect 458766 200898 468770 201134
rect 469006 200898 479010 201134
rect 479246 200898 489250 201134
rect 489486 200898 499490 201134
rect 499726 200898 509730 201134
rect 509966 200898 519970 201134
rect 520206 200898 530210 201134
rect 530446 200898 549666 201134
rect 549902 200898 549986 201134
rect 550222 200898 559906 201134
rect 560142 200898 560226 201134
rect 560462 200898 570146 201134
rect 570382 200898 570466 201134
rect 570702 200898 580386 201134
rect 580622 200898 580706 201134
rect 580942 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 545466 194614
rect 545702 194378 545786 194614
rect 546022 194378 555706 194614
rect 555942 194378 556026 194614
rect 556262 194378 565946 194614
rect 566182 194378 566266 194614
rect 566502 194378 576186 194614
rect 576422 194378 576506 194614
rect 576742 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 545466 194294
rect 545702 194058 545786 194294
rect 546022 194058 555706 194294
rect 555942 194058 556026 194294
rect 556262 194058 565946 194294
rect 566182 194058 566266 194294
rect 566502 194058 576186 194294
rect 576422 194058 576506 194294
rect 576742 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 541746 190894
rect 541982 190658 542066 190894
rect 542302 190658 551986 190894
rect 552222 190658 552306 190894
rect 552542 190658 562226 190894
rect 562462 190658 562546 190894
rect 562782 190658 572466 190894
rect 572702 190658 572786 190894
rect 573022 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 541746 190574
rect 541982 190338 542066 190574
rect 542302 190338 551986 190574
rect 552222 190338 552306 190574
rect 552542 190338 562226 190574
rect 562462 190338 562546 190574
rect 562782 190338 572466 190574
rect 572702 190338 572786 190574
rect 573022 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 15786 187174
rect 16022 186938 16106 187174
rect 16342 186938 548266 187174
rect 548502 186938 548586 187174
rect 548822 186938 558506 187174
rect 558742 186938 558826 187174
rect 559062 186938 568746 187174
rect 568982 186938 569066 187174
rect 569302 186938 578986 187174
rect 579222 186938 579306 187174
rect 579542 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 15786 186854
rect 16022 186618 16106 186854
rect 16342 186618 548266 186854
rect 548502 186618 548586 186854
rect 548822 186618 558506 186854
rect 558742 186618 558826 186854
rect 559062 186618 568746 186854
rect 568982 186618 569066 186854
rect 569302 186618 578986 186854
rect 579222 186618 579306 186854
rect 579542 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 12066 183454
rect 12302 183218 12386 183454
rect 12622 183218 23330 183454
rect 23566 183218 33570 183454
rect 33806 183218 43810 183454
rect 44046 183218 54050 183454
rect 54286 183218 64290 183454
rect 64526 183218 74530 183454
rect 74766 183218 84770 183454
rect 85006 183218 95010 183454
rect 95246 183218 105250 183454
rect 105486 183218 115490 183454
rect 115726 183218 125730 183454
rect 125966 183218 135970 183454
rect 136206 183218 146210 183454
rect 146446 183218 156450 183454
rect 156686 183218 166690 183454
rect 166926 183218 176930 183454
rect 177166 183218 187170 183454
rect 187406 183218 197410 183454
rect 197646 183218 207650 183454
rect 207886 183218 217890 183454
rect 218126 183218 228130 183454
rect 228366 183218 238370 183454
rect 238606 183218 248610 183454
rect 248846 183218 258850 183454
rect 259086 183218 269090 183454
rect 269326 183218 279330 183454
rect 279566 183218 289570 183454
rect 289806 183218 299810 183454
rect 300046 183218 310050 183454
rect 310286 183218 320290 183454
rect 320526 183218 330530 183454
rect 330766 183218 340770 183454
rect 341006 183218 351010 183454
rect 351246 183218 361250 183454
rect 361486 183218 371490 183454
rect 371726 183218 381730 183454
rect 381966 183218 391970 183454
rect 392206 183218 402210 183454
rect 402446 183218 412450 183454
rect 412686 183218 422690 183454
rect 422926 183218 432930 183454
rect 433166 183218 443170 183454
rect 443406 183218 453410 183454
rect 453646 183218 463650 183454
rect 463886 183218 473890 183454
rect 474126 183218 484130 183454
rect 484366 183218 494370 183454
rect 494606 183218 504610 183454
rect 504846 183218 514850 183454
rect 515086 183218 525090 183454
rect 525326 183218 535330 183454
rect 535566 183218 544546 183454
rect 544782 183218 544866 183454
rect 545102 183218 554786 183454
rect 555022 183218 555106 183454
rect 555342 183218 565026 183454
rect 565262 183218 565346 183454
rect 565582 183218 575266 183454
rect 575502 183218 575586 183454
rect 575822 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 12066 183134
rect 12302 182898 12386 183134
rect 12622 182898 23330 183134
rect 23566 182898 33570 183134
rect 33806 182898 43810 183134
rect 44046 182898 54050 183134
rect 54286 182898 64290 183134
rect 64526 182898 74530 183134
rect 74766 182898 84770 183134
rect 85006 182898 95010 183134
rect 95246 182898 105250 183134
rect 105486 182898 115490 183134
rect 115726 182898 125730 183134
rect 125966 182898 135970 183134
rect 136206 182898 146210 183134
rect 146446 182898 156450 183134
rect 156686 182898 166690 183134
rect 166926 182898 176930 183134
rect 177166 182898 187170 183134
rect 187406 182898 197410 183134
rect 197646 182898 207650 183134
rect 207886 182898 217890 183134
rect 218126 182898 228130 183134
rect 228366 182898 238370 183134
rect 238606 182898 248610 183134
rect 248846 182898 258850 183134
rect 259086 182898 269090 183134
rect 269326 182898 279330 183134
rect 279566 182898 289570 183134
rect 289806 182898 299810 183134
rect 300046 182898 310050 183134
rect 310286 182898 320290 183134
rect 320526 182898 330530 183134
rect 330766 182898 340770 183134
rect 341006 182898 351010 183134
rect 351246 182898 361250 183134
rect 361486 182898 371490 183134
rect 371726 182898 381730 183134
rect 381966 182898 391970 183134
rect 392206 182898 402210 183134
rect 402446 182898 412450 183134
rect 412686 182898 422690 183134
rect 422926 182898 432930 183134
rect 433166 182898 443170 183134
rect 443406 182898 453410 183134
rect 453646 182898 463650 183134
rect 463886 182898 473890 183134
rect 474126 182898 484130 183134
rect 484366 182898 494370 183134
rect 494606 182898 504610 183134
rect 504846 182898 514850 183134
rect 515086 182898 525090 183134
rect 525326 182898 535330 183134
rect 535566 182898 544546 183134
rect 544782 182898 544866 183134
rect 545102 182898 554786 183134
rect 555022 182898 555106 183134
rect 555342 182898 565026 183134
rect 565262 182898 565346 183134
rect 565582 182898 575266 183134
rect 575502 182898 575586 183134
rect 575822 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 550586 176614
rect 550822 176378 550906 176614
rect 551142 176378 560826 176614
rect 561062 176378 561146 176614
rect 561382 176378 571066 176614
rect 571302 176378 571386 176614
rect 571622 176378 581306 176614
rect 581542 176378 581626 176614
rect 581862 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 550586 176294
rect 550822 176058 550906 176294
rect 551142 176058 560826 176294
rect 561062 176058 561146 176294
rect 561382 176058 571066 176294
rect 571302 176058 571386 176294
rect 571622 176058 581306 176294
rect 581542 176058 581626 176294
rect 581862 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 14386 172894
rect 14622 172658 14706 172894
rect 14942 172658 546866 172894
rect 547102 172658 547186 172894
rect 547422 172658 557106 172894
rect 557342 172658 557426 172894
rect 557662 172658 567346 172894
rect 567582 172658 567666 172894
rect 567902 172658 577586 172894
rect 577822 172658 577906 172894
rect 578142 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 14386 172574
rect 14622 172338 14706 172574
rect 14942 172338 546866 172574
rect 547102 172338 547186 172574
rect 547422 172338 557106 172574
rect 557342 172338 557426 172574
rect 557662 172338 567346 172574
rect 567582 172338 567666 172574
rect 567902 172338 577586 172574
rect 577822 172338 577906 172574
rect 578142 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 10666 169174
rect 10902 168938 10986 169174
rect 11222 168938 543146 169174
rect 543382 168938 543466 169174
rect 543702 168938 553386 169174
rect 553622 168938 553706 169174
rect 553942 168938 563626 169174
rect 563862 168938 563946 169174
rect 564182 168938 573866 169174
rect 574102 168938 574186 169174
rect 574422 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 10666 168854
rect 10902 168618 10986 168854
rect 11222 168618 543146 168854
rect 543382 168618 543466 168854
rect 543702 168618 553386 168854
rect 553622 168618 553706 168854
rect 553942 168618 563626 168854
rect 563862 168618 563946 168854
rect 564182 168618 573866 168854
rect 574102 168618 574186 168854
rect 574422 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 6946 165454
rect 7182 165218 7266 165454
rect 7502 165218 28450 165454
rect 28686 165218 38690 165454
rect 38926 165218 48930 165454
rect 49166 165218 59170 165454
rect 59406 165218 69410 165454
rect 69646 165218 79650 165454
rect 79886 165218 89890 165454
rect 90126 165218 100130 165454
rect 100366 165218 110370 165454
rect 110606 165218 120610 165454
rect 120846 165218 130850 165454
rect 131086 165218 141090 165454
rect 141326 165218 151330 165454
rect 151566 165218 161570 165454
rect 161806 165218 171810 165454
rect 172046 165218 182050 165454
rect 182286 165218 192290 165454
rect 192526 165218 202530 165454
rect 202766 165218 212770 165454
rect 213006 165218 223010 165454
rect 223246 165218 233250 165454
rect 233486 165218 243490 165454
rect 243726 165218 253730 165454
rect 253966 165218 263970 165454
rect 264206 165218 274210 165454
rect 274446 165218 284450 165454
rect 284686 165218 294690 165454
rect 294926 165218 304930 165454
rect 305166 165218 315170 165454
rect 315406 165218 325410 165454
rect 325646 165218 335650 165454
rect 335886 165218 345890 165454
rect 346126 165218 356130 165454
rect 356366 165218 366370 165454
rect 366606 165218 376610 165454
rect 376846 165218 386850 165454
rect 387086 165218 397090 165454
rect 397326 165218 407330 165454
rect 407566 165218 417570 165454
rect 417806 165218 427810 165454
rect 428046 165218 438050 165454
rect 438286 165218 448290 165454
rect 448526 165218 458530 165454
rect 458766 165218 468770 165454
rect 469006 165218 479010 165454
rect 479246 165218 489250 165454
rect 489486 165218 499490 165454
rect 499726 165218 509730 165454
rect 509966 165218 519970 165454
rect 520206 165218 530210 165454
rect 530446 165218 549666 165454
rect 549902 165218 549986 165454
rect 550222 165218 559906 165454
rect 560142 165218 560226 165454
rect 560462 165218 570146 165454
rect 570382 165218 570466 165454
rect 570702 165218 580386 165454
rect 580622 165218 580706 165454
rect 580942 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 6946 165134
rect 7182 164898 7266 165134
rect 7502 164898 28450 165134
rect 28686 164898 38690 165134
rect 38926 164898 48930 165134
rect 49166 164898 59170 165134
rect 59406 164898 69410 165134
rect 69646 164898 79650 165134
rect 79886 164898 89890 165134
rect 90126 164898 100130 165134
rect 100366 164898 110370 165134
rect 110606 164898 120610 165134
rect 120846 164898 130850 165134
rect 131086 164898 141090 165134
rect 141326 164898 151330 165134
rect 151566 164898 161570 165134
rect 161806 164898 171810 165134
rect 172046 164898 182050 165134
rect 182286 164898 192290 165134
rect 192526 164898 202530 165134
rect 202766 164898 212770 165134
rect 213006 164898 223010 165134
rect 223246 164898 233250 165134
rect 233486 164898 243490 165134
rect 243726 164898 253730 165134
rect 253966 164898 263970 165134
rect 264206 164898 274210 165134
rect 274446 164898 284450 165134
rect 284686 164898 294690 165134
rect 294926 164898 304930 165134
rect 305166 164898 315170 165134
rect 315406 164898 325410 165134
rect 325646 164898 335650 165134
rect 335886 164898 345890 165134
rect 346126 164898 356130 165134
rect 356366 164898 366370 165134
rect 366606 164898 376610 165134
rect 376846 164898 386850 165134
rect 387086 164898 397090 165134
rect 397326 164898 407330 165134
rect 407566 164898 417570 165134
rect 417806 164898 427810 165134
rect 428046 164898 438050 165134
rect 438286 164898 448290 165134
rect 448526 164898 458530 165134
rect 458766 164898 468770 165134
rect 469006 164898 479010 165134
rect 479246 164898 489250 165134
rect 489486 164898 499490 165134
rect 499726 164898 509730 165134
rect 509966 164898 519970 165134
rect 520206 164898 530210 165134
rect 530446 164898 549666 165134
rect 549902 164898 549986 165134
rect 550222 164898 559906 165134
rect 560142 164898 560226 165134
rect 560462 164898 570146 165134
rect 570382 164898 570466 165134
rect 570702 164898 580386 165134
rect 580622 164898 580706 165134
rect 580942 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 545466 158614
rect 545702 158378 545786 158614
rect 546022 158378 555706 158614
rect 555942 158378 556026 158614
rect 556262 158378 565946 158614
rect 566182 158378 566266 158614
rect 566502 158378 576186 158614
rect 576422 158378 576506 158614
rect 576742 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 545466 158294
rect 545702 158058 545786 158294
rect 546022 158058 555706 158294
rect 555942 158058 556026 158294
rect 556262 158058 565946 158294
rect 566182 158058 566266 158294
rect 566502 158058 576186 158294
rect 576422 158058 576506 158294
rect 576742 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 541746 154894
rect 541982 154658 542066 154894
rect 542302 154658 551986 154894
rect 552222 154658 552306 154894
rect 552542 154658 562226 154894
rect 562462 154658 562546 154894
rect 562782 154658 572466 154894
rect 572702 154658 572786 154894
rect 573022 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 541746 154574
rect 541982 154338 542066 154574
rect 542302 154338 551986 154574
rect 552222 154338 552306 154574
rect 552542 154338 562226 154574
rect 562462 154338 562546 154574
rect 562782 154338 572466 154574
rect 572702 154338 572786 154574
rect 573022 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 15786 151174
rect 16022 150938 16106 151174
rect 16342 150938 548266 151174
rect 548502 150938 548586 151174
rect 548822 150938 558506 151174
rect 558742 150938 558826 151174
rect 559062 150938 568746 151174
rect 568982 150938 569066 151174
rect 569302 150938 578986 151174
rect 579222 150938 579306 151174
rect 579542 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 15786 150854
rect 16022 150618 16106 150854
rect 16342 150618 548266 150854
rect 548502 150618 548586 150854
rect 548822 150618 558506 150854
rect 558742 150618 558826 150854
rect 559062 150618 568746 150854
rect 568982 150618 569066 150854
rect 569302 150618 578986 150854
rect 579222 150618 579306 150854
rect 579542 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 12066 147454
rect 12302 147218 12386 147454
rect 12622 147218 23330 147454
rect 23566 147218 33570 147454
rect 33806 147218 43810 147454
rect 44046 147218 54050 147454
rect 54286 147218 64290 147454
rect 64526 147218 74530 147454
rect 74766 147218 84770 147454
rect 85006 147218 95010 147454
rect 95246 147218 105250 147454
rect 105486 147218 115490 147454
rect 115726 147218 125730 147454
rect 125966 147218 135970 147454
rect 136206 147218 146210 147454
rect 146446 147218 156450 147454
rect 156686 147218 166690 147454
rect 166926 147218 176930 147454
rect 177166 147218 187170 147454
rect 187406 147218 197410 147454
rect 197646 147218 207650 147454
rect 207886 147218 217890 147454
rect 218126 147218 228130 147454
rect 228366 147218 238370 147454
rect 238606 147218 248610 147454
rect 248846 147218 258850 147454
rect 259086 147218 269090 147454
rect 269326 147218 279330 147454
rect 279566 147218 289570 147454
rect 289806 147218 299810 147454
rect 300046 147218 310050 147454
rect 310286 147218 320290 147454
rect 320526 147218 330530 147454
rect 330766 147218 340770 147454
rect 341006 147218 351010 147454
rect 351246 147218 361250 147454
rect 361486 147218 371490 147454
rect 371726 147218 381730 147454
rect 381966 147218 391970 147454
rect 392206 147218 402210 147454
rect 402446 147218 412450 147454
rect 412686 147218 422690 147454
rect 422926 147218 432930 147454
rect 433166 147218 443170 147454
rect 443406 147218 453410 147454
rect 453646 147218 463650 147454
rect 463886 147218 473890 147454
rect 474126 147218 484130 147454
rect 484366 147218 494370 147454
rect 494606 147218 504610 147454
rect 504846 147218 514850 147454
rect 515086 147218 525090 147454
rect 525326 147218 535330 147454
rect 535566 147218 544546 147454
rect 544782 147218 544866 147454
rect 545102 147218 554786 147454
rect 555022 147218 555106 147454
rect 555342 147218 565026 147454
rect 565262 147218 565346 147454
rect 565582 147218 575266 147454
rect 575502 147218 575586 147454
rect 575822 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 12066 147134
rect 12302 146898 12386 147134
rect 12622 146898 23330 147134
rect 23566 146898 33570 147134
rect 33806 146898 43810 147134
rect 44046 146898 54050 147134
rect 54286 146898 64290 147134
rect 64526 146898 74530 147134
rect 74766 146898 84770 147134
rect 85006 146898 95010 147134
rect 95246 146898 105250 147134
rect 105486 146898 115490 147134
rect 115726 146898 125730 147134
rect 125966 146898 135970 147134
rect 136206 146898 146210 147134
rect 146446 146898 156450 147134
rect 156686 146898 166690 147134
rect 166926 146898 176930 147134
rect 177166 146898 187170 147134
rect 187406 146898 197410 147134
rect 197646 146898 207650 147134
rect 207886 146898 217890 147134
rect 218126 146898 228130 147134
rect 228366 146898 238370 147134
rect 238606 146898 248610 147134
rect 248846 146898 258850 147134
rect 259086 146898 269090 147134
rect 269326 146898 279330 147134
rect 279566 146898 289570 147134
rect 289806 146898 299810 147134
rect 300046 146898 310050 147134
rect 310286 146898 320290 147134
rect 320526 146898 330530 147134
rect 330766 146898 340770 147134
rect 341006 146898 351010 147134
rect 351246 146898 361250 147134
rect 361486 146898 371490 147134
rect 371726 146898 381730 147134
rect 381966 146898 391970 147134
rect 392206 146898 402210 147134
rect 402446 146898 412450 147134
rect 412686 146898 422690 147134
rect 422926 146898 432930 147134
rect 433166 146898 443170 147134
rect 443406 146898 453410 147134
rect 453646 146898 463650 147134
rect 463886 146898 473890 147134
rect 474126 146898 484130 147134
rect 484366 146898 494370 147134
rect 494606 146898 504610 147134
rect 504846 146898 514850 147134
rect 515086 146898 525090 147134
rect 525326 146898 535330 147134
rect 535566 146898 544546 147134
rect 544782 146898 544866 147134
rect 545102 146898 554786 147134
rect 555022 146898 555106 147134
rect 555342 146898 565026 147134
rect 565262 146898 565346 147134
rect 565582 146898 575266 147134
rect 575502 146898 575586 147134
rect 575822 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 550586 140614
rect 550822 140378 550906 140614
rect 551142 140378 560826 140614
rect 561062 140378 561146 140614
rect 561382 140378 571066 140614
rect 571302 140378 571386 140614
rect 571622 140378 581306 140614
rect 581542 140378 581626 140614
rect 581862 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 550586 140294
rect 550822 140058 550906 140294
rect 551142 140058 560826 140294
rect 561062 140058 561146 140294
rect 561382 140058 571066 140294
rect 571302 140058 571386 140294
rect 571622 140058 581306 140294
rect 581542 140058 581626 140294
rect 581862 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 14386 136894
rect 14622 136658 14706 136894
rect 14942 136658 546866 136894
rect 547102 136658 547186 136894
rect 547422 136658 557106 136894
rect 557342 136658 557426 136894
rect 557662 136658 567346 136894
rect 567582 136658 567666 136894
rect 567902 136658 577586 136894
rect 577822 136658 577906 136894
rect 578142 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 14386 136574
rect 14622 136338 14706 136574
rect 14942 136338 546866 136574
rect 547102 136338 547186 136574
rect 547422 136338 557106 136574
rect 557342 136338 557426 136574
rect 557662 136338 567346 136574
rect 567582 136338 567666 136574
rect 567902 136338 577586 136574
rect 577822 136338 577906 136574
rect 578142 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 10666 133174
rect 10902 132938 10986 133174
rect 11222 132938 543146 133174
rect 543382 132938 543466 133174
rect 543702 132938 553386 133174
rect 553622 132938 553706 133174
rect 553942 132938 563626 133174
rect 563862 132938 563946 133174
rect 564182 132938 573866 133174
rect 574102 132938 574186 133174
rect 574422 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 10666 132854
rect 10902 132618 10986 132854
rect 11222 132618 543146 132854
rect 543382 132618 543466 132854
rect 543702 132618 553386 132854
rect 553622 132618 553706 132854
rect 553942 132618 563626 132854
rect 563862 132618 563946 132854
rect 564182 132618 573866 132854
rect 574102 132618 574186 132854
rect 574422 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 6946 129454
rect 7182 129218 7266 129454
rect 7502 129218 28450 129454
rect 28686 129218 38690 129454
rect 38926 129218 48930 129454
rect 49166 129218 59170 129454
rect 59406 129218 69410 129454
rect 69646 129218 79650 129454
rect 79886 129218 89890 129454
rect 90126 129218 100130 129454
rect 100366 129218 110370 129454
rect 110606 129218 120610 129454
rect 120846 129218 130850 129454
rect 131086 129218 141090 129454
rect 141326 129218 151330 129454
rect 151566 129218 161570 129454
rect 161806 129218 171810 129454
rect 172046 129218 182050 129454
rect 182286 129218 192290 129454
rect 192526 129218 202530 129454
rect 202766 129218 212770 129454
rect 213006 129218 223010 129454
rect 223246 129218 233250 129454
rect 233486 129218 243490 129454
rect 243726 129218 253730 129454
rect 253966 129218 263970 129454
rect 264206 129218 274210 129454
rect 274446 129218 284450 129454
rect 284686 129218 294690 129454
rect 294926 129218 304930 129454
rect 305166 129218 315170 129454
rect 315406 129218 325410 129454
rect 325646 129218 335650 129454
rect 335886 129218 345890 129454
rect 346126 129218 356130 129454
rect 356366 129218 366370 129454
rect 366606 129218 376610 129454
rect 376846 129218 386850 129454
rect 387086 129218 397090 129454
rect 397326 129218 407330 129454
rect 407566 129218 417570 129454
rect 417806 129218 427810 129454
rect 428046 129218 438050 129454
rect 438286 129218 448290 129454
rect 448526 129218 458530 129454
rect 458766 129218 468770 129454
rect 469006 129218 479010 129454
rect 479246 129218 489250 129454
rect 489486 129218 499490 129454
rect 499726 129218 509730 129454
rect 509966 129218 519970 129454
rect 520206 129218 530210 129454
rect 530446 129218 549666 129454
rect 549902 129218 549986 129454
rect 550222 129218 559906 129454
rect 560142 129218 560226 129454
rect 560462 129218 570146 129454
rect 570382 129218 570466 129454
rect 570702 129218 580386 129454
rect 580622 129218 580706 129454
rect 580942 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 6946 129134
rect 7182 128898 7266 129134
rect 7502 128898 28450 129134
rect 28686 128898 38690 129134
rect 38926 128898 48930 129134
rect 49166 128898 59170 129134
rect 59406 128898 69410 129134
rect 69646 128898 79650 129134
rect 79886 128898 89890 129134
rect 90126 128898 100130 129134
rect 100366 128898 110370 129134
rect 110606 128898 120610 129134
rect 120846 128898 130850 129134
rect 131086 128898 141090 129134
rect 141326 128898 151330 129134
rect 151566 128898 161570 129134
rect 161806 128898 171810 129134
rect 172046 128898 182050 129134
rect 182286 128898 192290 129134
rect 192526 128898 202530 129134
rect 202766 128898 212770 129134
rect 213006 128898 223010 129134
rect 223246 128898 233250 129134
rect 233486 128898 243490 129134
rect 243726 128898 253730 129134
rect 253966 128898 263970 129134
rect 264206 128898 274210 129134
rect 274446 128898 284450 129134
rect 284686 128898 294690 129134
rect 294926 128898 304930 129134
rect 305166 128898 315170 129134
rect 315406 128898 325410 129134
rect 325646 128898 335650 129134
rect 335886 128898 345890 129134
rect 346126 128898 356130 129134
rect 356366 128898 366370 129134
rect 366606 128898 376610 129134
rect 376846 128898 386850 129134
rect 387086 128898 397090 129134
rect 397326 128898 407330 129134
rect 407566 128898 417570 129134
rect 417806 128898 427810 129134
rect 428046 128898 438050 129134
rect 438286 128898 448290 129134
rect 448526 128898 458530 129134
rect 458766 128898 468770 129134
rect 469006 128898 479010 129134
rect 479246 128898 489250 129134
rect 489486 128898 499490 129134
rect 499726 128898 509730 129134
rect 509966 128898 519970 129134
rect 520206 128898 530210 129134
rect 530446 128898 549666 129134
rect 549902 128898 549986 129134
rect 550222 128898 559906 129134
rect 560142 128898 560226 129134
rect 560462 128898 570146 129134
rect 570382 128898 570466 129134
rect 570702 128898 580386 129134
rect 580622 128898 580706 129134
rect 580942 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 545466 122614
rect 545702 122378 545786 122614
rect 546022 122378 555706 122614
rect 555942 122378 556026 122614
rect 556262 122378 565946 122614
rect 566182 122378 566266 122614
rect 566502 122378 576186 122614
rect 576422 122378 576506 122614
rect 576742 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 545466 122294
rect 545702 122058 545786 122294
rect 546022 122058 555706 122294
rect 555942 122058 556026 122294
rect 556262 122058 565946 122294
rect 566182 122058 566266 122294
rect 566502 122058 576186 122294
rect 576422 122058 576506 122294
rect 576742 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 541746 118894
rect 541982 118658 542066 118894
rect 542302 118658 551986 118894
rect 552222 118658 552306 118894
rect 552542 118658 562226 118894
rect 562462 118658 562546 118894
rect 562782 118658 572466 118894
rect 572702 118658 572786 118894
rect 573022 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 541746 118574
rect 541982 118338 542066 118574
rect 542302 118338 551986 118574
rect 552222 118338 552306 118574
rect 552542 118338 562226 118574
rect 562462 118338 562546 118574
rect 562782 118338 572466 118574
rect 572702 118338 572786 118574
rect 573022 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 15786 115174
rect 16022 114938 16106 115174
rect 16342 114938 548266 115174
rect 548502 114938 548586 115174
rect 548822 114938 558506 115174
rect 558742 114938 558826 115174
rect 559062 114938 568746 115174
rect 568982 114938 569066 115174
rect 569302 114938 578986 115174
rect 579222 114938 579306 115174
rect 579542 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 15786 114854
rect 16022 114618 16106 114854
rect 16342 114618 548266 114854
rect 548502 114618 548586 114854
rect 548822 114618 558506 114854
rect 558742 114618 558826 114854
rect 559062 114618 568746 114854
rect 568982 114618 569066 114854
rect 569302 114618 578986 114854
rect 579222 114618 579306 114854
rect 579542 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 12066 111454
rect 12302 111218 12386 111454
rect 12622 111218 23330 111454
rect 23566 111218 33570 111454
rect 33806 111218 43810 111454
rect 44046 111218 54050 111454
rect 54286 111218 64290 111454
rect 64526 111218 74530 111454
rect 74766 111218 84770 111454
rect 85006 111218 95010 111454
rect 95246 111218 105250 111454
rect 105486 111218 115490 111454
rect 115726 111218 125730 111454
rect 125966 111218 135970 111454
rect 136206 111218 146210 111454
rect 146446 111218 156450 111454
rect 156686 111218 166690 111454
rect 166926 111218 176930 111454
rect 177166 111218 187170 111454
rect 187406 111218 197410 111454
rect 197646 111218 207650 111454
rect 207886 111218 217890 111454
rect 218126 111218 228130 111454
rect 228366 111218 238370 111454
rect 238606 111218 248610 111454
rect 248846 111218 258850 111454
rect 259086 111218 269090 111454
rect 269326 111218 279330 111454
rect 279566 111218 289570 111454
rect 289806 111218 299810 111454
rect 300046 111218 310050 111454
rect 310286 111218 320290 111454
rect 320526 111218 330530 111454
rect 330766 111218 340770 111454
rect 341006 111218 351010 111454
rect 351246 111218 361250 111454
rect 361486 111218 371490 111454
rect 371726 111218 381730 111454
rect 381966 111218 391970 111454
rect 392206 111218 402210 111454
rect 402446 111218 412450 111454
rect 412686 111218 422690 111454
rect 422926 111218 432930 111454
rect 433166 111218 443170 111454
rect 443406 111218 453410 111454
rect 453646 111218 463650 111454
rect 463886 111218 473890 111454
rect 474126 111218 484130 111454
rect 484366 111218 494370 111454
rect 494606 111218 504610 111454
rect 504846 111218 514850 111454
rect 515086 111218 525090 111454
rect 525326 111218 535330 111454
rect 535566 111218 544546 111454
rect 544782 111218 544866 111454
rect 545102 111218 554786 111454
rect 555022 111218 555106 111454
rect 555342 111218 565026 111454
rect 565262 111218 565346 111454
rect 565582 111218 575266 111454
rect 575502 111218 575586 111454
rect 575822 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 12066 111134
rect 12302 110898 12386 111134
rect 12622 110898 23330 111134
rect 23566 110898 33570 111134
rect 33806 110898 43810 111134
rect 44046 110898 54050 111134
rect 54286 110898 64290 111134
rect 64526 110898 74530 111134
rect 74766 110898 84770 111134
rect 85006 110898 95010 111134
rect 95246 110898 105250 111134
rect 105486 110898 115490 111134
rect 115726 110898 125730 111134
rect 125966 110898 135970 111134
rect 136206 110898 146210 111134
rect 146446 110898 156450 111134
rect 156686 110898 166690 111134
rect 166926 110898 176930 111134
rect 177166 110898 187170 111134
rect 187406 110898 197410 111134
rect 197646 110898 207650 111134
rect 207886 110898 217890 111134
rect 218126 110898 228130 111134
rect 228366 110898 238370 111134
rect 238606 110898 248610 111134
rect 248846 110898 258850 111134
rect 259086 110898 269090 111134
rect 269326 110898 279330 111134
rect 279566 110898 289570 111134
rect 289806 110898 299810 111134
rect 300046 110898 310050 111134
rect 310286 110898 320290 111134
rect 320526 110898 330530 111134
rect 330766 110898 340770 111134
rect 341006 110898 351010 111134
rect 351246 110898 361250 111134
rect 361486 110898 371490 111134
rect 371726 110898 381730 111134
rect 381966 110898 391970 111134
rect 392206 110898 402210 111134
rect 402446 110898 412450 111134
rect 412686 110898 422690 111134
rect 422926 110898 432930 111134
rect 433166 110898 443170 111134
rect 443406 110898 453410 111134
rect 453646 110898 463650 111134
rect 463886 110898 473890 111134
rect 474126 110898 484130 111134
rect 484366 110898 494370 111134
rect 494606 110898 504610 111134
rect 504846 110898 514850 111134
rect 515086 110898 525090 111134
rect 525326 110898 535330 111134
rect 535566 110898 544546 111134
rect 544782 110898 544866 111134
rect 545102 110898 554786 111134
rect 555022 110898 555106 111134
rect 555342 110898 565026 111134
rect 565262 110898 565346 111134
rect 565582 110898 575266 111134
rect 575502 110898 575586 111134
rect 575822 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 550586 104614
rect 550822 104378 550906 104614
rect 551142 104378 560826 104614
rect 561062 104378 561146 104614
rect 561382 104378 571066 104614
rect 571302 104378 571386 104614
rect 571622 104378 581306 104614
rect 581542 104378 581626 104614
rect 581862 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 550586 104294
rect 550822 104058 550906 104294
rect 551142 104058 560826 104294
rect 561062 104058 561146 104294
rect 561382 104058 571066 104294
rect 571302 104058 571386 104294
rect 571622 104058 581306 104294
rect 581542 104058 581626 104294
rect 581862 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 14386 100894
rect 14622 100658 14706 100894
rect 14942 100658 546866 100894
rect 547102 100658 547186 100894
rect 547422 100658 557106 100894
rect 557342 100658 557426 100894
rect 557662 100658 567346 100894
rect 567582 100658 567666 100894
rect 567902 100658 577586 100894
rect 577822 100658 577906 100894
rect 578142 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 14386 100574
rect 14622 100338 14706 100574
rect 14942 100338 546866 100574
rect 547102 100338 547186 100574
rect 547422 100338 557106 100574
rect 557342 100338 557426 100574
rect 557662 100338 567346 100574
rect 567582 100338 567666 100574
rect 567902 100338 577586 100574
rect 577822 100338 577906 100574
rect 578142 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 10666 97174
rect 10902 96938 10986 97174
rect 11222 96938 543146 97174
rect 543382 96938 543466 97174
rect 543702 96938 553386 97174
rect 553622 96938 553706 97174
rect 553942 96938 563626 97174
rect 563862 96938 563946 97174
rect 564182 96938 573866 97174
rect 574102 96938 574186 97174
rect 574422 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 10666 96854
rect 10902 96618 10986 96854
rect 11222 96618 543146 96854
rect 543382 96618 543466 96854
rect 543702 96618 553386 96854
rect 553622 96618 553706 96854
rect 553942 96618 563626 96854
rect 563862 96618 563946 96854
rect 564182 96618 573866 96854
rect 574102 96618 574186 96854
rect 574422 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 6946 93454
rect 7182 93218 7266 93454
rect 7502 93218 28450 93454
rect 28686 93218 38690 93454
rect 38926 93218 48930 93454
rect 49166 93218 59170 93454
rect 59406 93218 69410 93454
rect 69646 93218 79650 93454
rect 79886 93218 89890 93454
rect 90126 93218 100130 93454
rect 100366 93218 110370 93454
rect 110606 93218 120610 93454
rect 120846 93218 130850 93454
rect 131086 93218 141090 93454
rect 141326 93218 151330 93454
rect 151566 93218 161570 93454
rect 161806 93218 171810 93454
rect 172046 93218 182050 93454
rect 182286 93218 192290 93454
rect 192526 93218 202530 93454
rect 202766 93218 212770 93454
rect 213006 93218 223010 93454
rect 223246 93218 233250 93454
rect 233486 93218 243490 93454
rect 243726 93218 253730 93454
rect 253966 93218 263970 93454
rect 264206 93218 274210 93454
rect 274446 93218 284450 93454
rect 284686 93218 294690 93454
rect 294926 93218 304930 93454
rect 305166 93218 315170 93454
rect 315406 93218 325410 93454
rect 325646 93218 335650 93454
rect 335886 93218 345890 93454
rect 346126 93218 356130 93454
rect 356366 93218 366370 93454
rect 366606 93218 376610 93454
rect 376846 93218 386850 93454
rect 387086 93218 397090 93454
rect 397326 93218 407330 93454
rect 407566 93218 417570 93454
rect 417806 93218 427810 93454
rect 428046 93218 438050 93454
rect 438286 93218 448290 93454
rect 448526 93218 458530 93454
rect 458766 93218 468770 93454
rect 469006 93218 479010 93454
rect 479246 93218 489250 93454
rect 489486 93218 499490 93454
rect 499726 93218 509730 93454
rect 509966 93218 519970 93454
rect 520206 93218 530210 93454
rect 530446 93218 549666 93454
rect 549902 93218 549986 93454
rect 550222 93218 559906 93454
rect 560142 93218 560226 93454
rect 560462 93218 570146 93454
rect 570382 93218 570466 93454
rect 570702 93218 580386 93454
rect 580622 93218 580706 93454
rect 580942 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 6946 93134
rect 7182 92898 7266 93134
rect 7502 92898 28450 93134
rect 28686 92898 38690 93134
rect 38926 92898 48930 93134
rect 49166 92898 59170 93134
rect 59406 92898 69410 93134
rect 69646 92898 79650 93134
rect 79886 92898 89890 93134
rect 90126 92898 100130 93134
rect 100366 92898 110370 93134
rect 110606 92898 120610 93134
rect 120846 92898 130850 93134
rect 131086 92898 141090 93134
rect 141326 92898 151330 93134
rect 151566 92898 161570 93134
rect 161806 92898 171810 93134
rect 172046 92898 182050 93134
rect 182286 92898 192290 93134
rect 192526 92898 202530 93134
rect 202766 92898 212770 93134
rect 213006 92898 223010 93134
rect 223246 92898 233250 93134
rect 233486 92898 243490 93134
rect 243726 92898 253730 93134
rect 253966 92898 263970 93134
rect 264206 92898 274210 93134
rect 274446 92898 284450 93134
rect 284686 92898 294690 93134
rect 294926 92898 304930 93134
rect 305166 92898 315170 93134
rect 315406 92898 325410 93134
rect 325646 92898 335650 93134
rect 335886 92898 345890 93134
rect 346126 92898 356130 93134
rect 356366 92898 366370 93134
rect 366606 92898 376610 93134
rect 376846 92898 386850 93134
rect 387086 92898 397090 93134
rect 397326 92898 407330 93134
rect 407566 92898 417570 93134
rect 417806 92898 427810 93134
rect 428046 92898 438050 93134
rect 438286 92898 448290 93134
rect 448526 92898 458530 93134
rect 458766 92898 468770 93134
rect 469006 92898 479010 93134
rect 479246 92898 489250 93134
rect 489486 92898 499490 93134
rect 499726 92898 509730 93134
rect 509966 92898 519970 93134
rect 520206 92898 530210 93134
rect 530446 92898 549666 93134
rect 549902 92898 549986 93134
rect 550222 92898 559906 93134
rect 560142 92898 560226 93134
rect 560462 92898 570146 93134
rect 570382 92898 570466 93134
rect 570702 92898 580386 93134
rect 580622 92898 580706 93134
rect 580942 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 545466 86614
rect 545702 86378 545786 86614
rect 546022 86378 555706 86614
rect 555942 86378 556026 86614
rect 556262 86378 565946 86614
rect 566182 86378 566266 86614
rect 566502 86378 576186 86614
rect 576422 86378 576506 86614
rect 576742 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 545466 86294
rect 545702 86058 545786 86294
rect 546022 86058 555706 86294
rect 555942 86058 556026 86294
rect 556262 86058 565946 86294
rect 566182 86058 566266 86294
rect 566502 86058 576186 86294
rect 576422 86058 576506 86294
rect 576742 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 541746 82894
rect 541982 82658 542066 82894
rect 542302 82658 551986 82894
rect 552222 82658 552306 82894
rect 552542 82658 562226 82894
rect 562462 82658 562546 82894
rect 562782 82658 572466 82894
rect 572702 82658 572786 82894
rect 573022 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 541746 82574
rect 541982 82338 542066 82574
rect 542302 82338 551986 82574
rect 552222 82338 552306 82574
rect 552542 82338 562226 82574
rect 562462 82338 562546 82574
rect 562782 82338 572466 82574
rect 572702 82338 572786 82574
rect 573022 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 15786 79174
rect 16022 78938 16106 79174
rect 16342 78938 548266 79174
rect 548502 78938 548586 79174
rect 548822 78938 558506 79174
rect 558742 78938 558826 79174
rect 559062 78938 568746 79174
rect 568982 78938 569066 79174
rect 569302 78938 578986 79174
rect 579222 78938 579306 79174
rect 579542 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 15786 78854
rect 16022 78618 16106 78854
rect 16342 78618 548266 78854
rect 548502 78618 548586 78854
rect 548822 78618 558506 78854
rect 558742 78618 558826 78854
rect 559062 78618 568746 78854
rect 568982 78618 569066 78854
rect 569302 78618 578986 78854
rect 579222 78618 579306 78854
rect 579542 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 12066 75454
rect 12302 75218 12386 75454
rect 12622 75218 23330 75454
rect 23566 75218 33570 75454
rect 33806 75218 43810 75454
rect 44046 75218 54050 75454
rect 54286 75218 64290 75454
rect 64526 75218 74530 75454
rect 74766 75218 84770 75454
rect 85006 75218 95010 75454
rect 95246 75218 105250 75454
rect 105486 75218 115490 75454
rect 115726 75218 125730 75454
rect 125966 75218 135970 75454
rect 136206 75218 146210 75454
rect 146446 75218 156450 75454
rect 156686 75218 166690 75454
rect 166926 75218 176930 75454
rect 177166 75218 187170 75454
rect 187406 75218 197410 75454
rect 197646 75218 207650 75454
rect 207886 75218 217890 75454
rect 218126 75218 228130 75454
rect 228366 75218 238370 75454
rect 238606 75218 248610 75454
rect 248846 75218 258850 75454
rect 259086 75218 269090 75454
rect 269326 75218 279330 75454
rect 279566 75218 289570 75454
rect 289806 75218 299810 75454
rect 300046 75218 310050 75454
rect 310286 75218 320290 75454
rect 320526 75218 330530 75454
rect 330766 75218 340770 75454
rect 341006 75218 351010 75454
rect 351246 75218 361250 75454
rect 361486 75218 371490 75454
rect 371726 75218 381730 75454
rect 381966 75218 391970 75454
rect 392206 75218 402210 75454
rect 402446 75218 412450 75454
rect 412686 75218 422690 75454
rect 422926 75218 432930 75454
rect 433166 75218 443170 75454
rect 443406 75218 453410 75454
rect 453646 75218 463650 75454
rect 463886 75218 473890 75454
rect 474126 75218 484130 75454
rect 484366 75218 494370 75454
rect 494606 75218 504610 75454
rect 504846 75218 514850 75454
rect 515086 75218 525090 75454
rect 525326 75218 535330 75454
rect 535566 75218 544546 75454
rect 544782 75218 544866 75454
rect 545102 75218 554786 75454
rect 555022 75218 555106 75454
rect 555342 75218 565026 75454
rect 565262 75218 565346 75454
rect 565582 75218 575266 75454
rect 575502 75218 575586 75454
rect 575822 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 12066 75134
rect 12302 74898 12386 75134
rect 12622 74898 23330 75134
rect 23566 74898 33570 75134
rect 33806 74898 43810 75134
rect 44046 74898 54050 75134
rect 54286 74898 64290 75134
rect 64526 74898 74530 75134
rect 74766 74898 84770 75134
rect 85006 74898 95010 75134
rect 95246 74898 105250 75134
rect 105486 74898 115490 75134
rect 115726 74898 125730 75134
rect 125966 74898 135970 75134
rect 136206 74898 146210 75134
rect 146446 74898 156450 75134
rect 156686 74898 166690 75134
rect 166926 74898 176930 75134
rect 177166 74898 187170 75134
rect 187406 74898 197410 75134
rect 197646 74898 207650 75134
rect 207886 74898 217890 75134
rect 218126 74898 228130 75134
rect 228366 74898 238370 75134
rect 238606 74898 248610 75134
rect 248846 74898 258850 75134
rect 259086 74898 269090 75134
rect 269326 74898 279330 75134
rect 279566 74898 289570 75134
rect 289806 74898 299810 75134
rect 300046 74898 310050 75134
rect 310286 74898 320290 75134
rect 320526 74898 330530 75134
rect 330766 74898 340770 75134
rect 341006 74898 351010 75134
rect 351246 74898 361250 75134
rect 361486 74898 371490 75134
rect 371726 74898 381730 75134
rect 381966 74898 391970 75134
rect 392206 74898 402210 75134
rect 402446 74898 412450 75134
rect 412686 74898 422690 75134
rect 422926 74898 432930 75134
rect 433166 74898 443170 75134
rect 443406 74898 453410 75134
rect 453646 74898 463650 75134
rect 463886 74898 473890 75134
rect 474126 74898 484130 75134
rect 484366 74898 494370 75134
rect 494606 74898 504610 75134
rect 504846 74898 514850 75134
rect 515086 74898 525090 75134
rect 525326 74898 535330 75134
rect 535566 74898 544546 75134
rect 544782 74898 544866 75134
rect 545102 74898 554786 75134
rect 555022 74898 555106 75134
rect 555342 74898 565026 75134
rect 565262 74898 565346 75134
rect 565582 74898 575266 75134
rect 575502 74898 575586 75134
rect 575822 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 550586 68614
rect 550822 68378 550906 68614
rect 551142 68378 560826 68614
rect 561062 68378 561146 68614
rect 561382 68378 571066 68614
rect 571302 68378 571386 68614
rect 571622 68378 581306 68614
rect 581542 68378 581626 68614
rect 581862 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 550586 68294
rect 550822 68058 550906 68294
rect 551142 68058 560826 68294
rect 561062 68058 561146 68294
rect 561382 68058 571066 68294
rect 571302 68058 571386 68294
rect 571622 68058 581306 68294
rect 581542 68058 581626 68294
rect 581862 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 14386 64894
rect 14622 64658 14706 64894
rect 14942 64658 546866 64894
rect 547102 64658 547186 64894
rect 547422 64658 557106 64894
rect 557342 64658 557426 64894
rect 557662 64658 567346 64894
rect 567582 64658 567666 64894
rect 567902 64658 577586 64894
rect 577822 64658 577906 64894
rect 578142 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 14386 64574
rect 14622 64338 14706 64574
rect 14942 64338 546866 64574
rect 547102 64338 547186 64574
rect 547422 64338 557106 64574
rect 557342 64338 557426 64574
rect 557662 64338 567346 64574
rect 567582 64338 567666 64574
rect 567902 64338 577586 64574
rect 577822 64338 577906 64574
rect 578142 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 10666 61174
rect 10902 60938 10986 61174
rect 11222 60938 543146 61174
rect 543382 60938 543466 61174
rect 543702 60938 553386 61174
rect 553622 60938 553706 61174
rect 553942 60938 563626 61174
rect 563862 60938 563946 61174
rect 564182 60938 573866 61174
rect 574102 60938 574186 61174
rect 574422 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 10666 60854
rect 10902 60618 10986 60854
rect 11222 60618 543146 60854
rect 543382 60618 543466 60854
rect 543702 60618 553386 60854
rect 553622 60618 553706 60854
rect 553942 60618 563626 60854
rect 563862 60618 563946 60854
rect 564182 60618 573866 60854
rect 574102 60618 574186 60854
rect 574422 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 6946 57454
rect 7182 57218 7266 57454
rect 7502 57218 28450 57454
rect 28686 57218 38690 57454
rect 38926 57218 48930 57454
rect 49166 57218 59170 57454
rect 59406 57218 69410 57454
rect 69646 57218 79650 57454
rect 79886 57218 89890 57454
rect 90126 57218 100130 57454
rect 100366 57218 110370 57454
rect 110606 57218 120610 57454
rect 120846 57218 130850 57454
rect 131086 57218 141090 57454
rect 141326 57218 151330 57454
rect 151566 57218 161570 57454
rect 161806 57218 171810 57454
rect 172046 57218 182050 57454
rect 182286 57218 192290 57454
rect 192526 57218 202530 57454
rect 202766 57218 212770 57454
rect 213006 57218 223010 57454
rect 223246 57218 233250 57454
rect 233486 57218 243490 57454
rect 243726 57218 253730 57454
rect 253966 57218 263970 57454
rect 264206 57218 274210 57454
rect 274446 57218 284450 57454
rect 284686 57218 294690 57454
rect 294926 57218 304930 57454
rect 305166 57218 315170 57454
rect 315406 57218 325410 57454
rect 325646 57218 335650 57454
rect 335886 57218 345890 57454
rect 346126 57218 356130 57454
rect 356366 57218 366370 57454
rect 366606 57218 376610 57454
rect 376846 57218 386850 57454
rect 387086 57218 397090 57454
rect 397326 57218 407330 57454
rect 407566 57218 417570 57454
rect 417806 57218 427810 57454
rect 428046 57218 438050 57454
rect 438286 57218 448290 57454
rect 448526 57218 458530 57454
rect 458766 57218 468770 57454
rect 469006 57218 479010 57454
rect 479246 57218 489250 57454
rect 489486 57218 499490 57454
rect 499726 57218 509730 57454
rect 509966 57218 519970 57454
rect 520206 57218 530210 57454
rect 530446 57218 549666 57454
rect 549902 57218 549986 57454
rect 550222 57218 559906 57454
rect 560142 57218 560226 57454
rect 560462 57218 570146 57454
rect 570382 57218 570466 57454
rect 570702 57218 580386 57454
rect 580622 57218 580706 57454
rect 580942 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 6946 57134
rect 7182 56898 7266 57134
rect 7502 56898 28450 57134
rect 28686 56898 38690 57134
rect 38926 56898 48930 57134
rect 49166 56898 59170 57134
rect 59406 56898 69410 57134
rect 69646 56898 79650 57134
rect 79886 56898 89890 57134
rect 90126 56898 100130 57134
rect 100366 56898 110370 57134
rect 110606 56898 120610 57134
rect 120846 56898 130850 57134
rect 131086 56898 141090 57134
rect 141326 56898 151330 57134
rect 151566 56898 161570 57134
rect 161806 56898 171810 57134
rect 172046 56898 182050 57134
rect 182286 56898 192290 57134
rect 192526 56898 202530 57134
rect 202766 56898 212770 57134
rect 213006 56898 223010 57134
rect 223246 56898 233250 57134
rect 233486 56898 243490 57134
rect 243726 56898 253730 57134
rect 253966 56898 263970 57134
rect 264206 56898 274210 57134
rect 274446 56898 284450 57134
rect 284686 56898 294690 57134
rect 294926 56898 304930 57134
rect 305166 56898 315170 57134
rect 315406 56898 325410 57134
rect 325646 56898 335650 57134
rect 335886 56898 345890 57134
rect 346126 56898 356130 57134
rect 356366 56898 366370 57134
rect 366606 56898 376610 57134
rect 376846 56898 386850 57134
rect 387086 56898 397090 57134
rect 397326 56898 407330 57134
rect 407566 56898 417570 57134
rect 417806 56898 427810 57134
rect 428046 56898 438050 57134
rect 438286 56898 448290 57134
rect 448526 56898 458530 57134
rect 458766 56898 468770 57134
rect 469006 56898 479010 57134
rect 479246 56898 489250 57134
rect 489486 56898 499490 57134
rect 499726 56898 509730 57134
rect 509966 56898 519970 57134
rect 520206 56898 530210 57134
rect 530446 56898 549666 57134
rect 549902 56898 549986 57134
rect 550222 56898 559906 57134
rect 560142 56898 560226 57134
rect 560462 56898 570146 57134
rect 570382 56898 570466 57134
rect 570702 56898 580386 57134
rect 580622 56898 580706 57134
rect 580942 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 545466 50614
rect 545702 50378 545786 50614
rect 546022 50378 555706 50614
rect 555942 50378 556026 50614
rect 556262 50378 565946 50614
rect 566182 50378 566266 50614
rect 566502 50378 576186 50614
rect 576422 50378 576506 50614
rect 576742 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 545466 50294
rect 545702 50058 545786 50294
rect 546022 50058 555706 50294
rect 555942 50058 556026 50294
rect 556262 50058 565946 50294
rect 566182 50058 566266 50294
rect 566502 50058 576186 50294
rect 576422 50058 576506 50294
rect 576742 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 541746 46894
rect 541982 46658 542066 46894
rect 542302 46658 551986 46894
rect 552222 46658 552306 46894
rect 552542 46658 562226 46894
rect 562462 46658 562546 46894
rect 562782 46658 572466 46894
rect 572702 46658 572786 46894
rect 573022 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 541746 46574
rect 541982 46338 542066 46574
rect 542302 46338 551986 46574
rect 552222 46338 552306 46574
rect 552542 46338 562226 46574
rect 562462 46338 562546 46574
rect 562782 46338 572466 46574
rect 572702 46338 572786 46574
rect 573022 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 15786 43174
rect 16022 42938 16106 43174
rect 16342 42938 548266 43174
rect 548502 42938 548586 43174
rect 548822 42938 558506 43174
rect 558742 42938 558826 43174
rect 559062 42938 568746 43174
rect 568982 42938 569066 43174
rect 569302 42938 578986 43174
rect 579222 42938 579306 43174
rect 579542 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 15786 42854
rect 16022 42618 16106 42854
rect 16342 42618 548266 42854
rect 548502 42618 548586 42854
rect 548822 42618 558506 42854
rect 558742 42618 558826 42854
rect 559062 42618 568746 42854
rect 568982 42618 569066 42854
rect 569302 42618 578986 42854
rect 579222 42618 579306 42854
rect 579542 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 12066 39454
rect 12302 39218 12386 39454
rect 12622 39218 23330 39454
rect 23566 39218 33570 39454
rect 33806 39218 43810 39454
rect 44046 39218 54050 39454
rect 54286 39218 64290 39454
rect 64526 39218 74530 39454
rect 74766 39218 84770 39454
rect 85006 39218 95010 39454
rect 95246 39218 105250 39454
rect 105486 39218 115490 39454
rect 115726 39218 125730 39454
rect 125966 39218 135970 39454
rect 136206 39218 146210 39454
rect 146446 39218 156450 39454
rect 156686 39218 166690 39454
rect 166926 39218 176930 39454
rect 177166 39218 187170 39454
rect 187406 39218 197410 39454
rect 197646 39218 207650 39454
rect 207886 39218 217890 39454
rect 218126 39218 228130 39454
rect 228366 39218 238370 39454
rect 238606 39218 248610 39454
rect 248846 39218 258850 39454
rect 259086 39218 269090 39454
rect 269326 39218 279330 39454
rect 279566 39218 289570 39454
rect 289806 39218 299810 39454
rect 300046 39218 310050 39454
rect 310286 39218 320290 39454
rect 320526 39218 330530 39454
rect 330766 39218 340770 39454
rect 341006 39218 351010 39454
rect 351246 39218 361250 39454
rect 361486 39218 371490 39454
rect 371726 39218 381730 39454
rect 381966 39218 391970 39454
rect 392206 39218 402210 39454
rect 402446 39218 412450 39454
rect 412686 39218 422690 39454
rect 422926 39218 432930 39454
rect 433166 39218 443170 39454
rect 443406 39218 453410 39454
rect 453646 39218 463650 39454
rect 463886 39218 473890 39454
rect 474126 39218 484130 39454
rect 484366 39218 494370 39454
rect 494606 39218 504610 39454
rect 504846 39218 514850 39454
rect 515086 39218 525090 39454
rect 525326 39218 535330 39454
rect 535566 39218 544546 39454
rect 544782 39218 544866 39454
rect 545102 39218 554786 39454
rect 555022 39218 555106 39454
rect 555342 39218 565026 39454
rect 565262 39218 565346 39454
rect 565582 39218 575266 39454
rect 575502 39218 575586 39454
rect 575822 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 12066 39134
rect 12302 38898 12386 39134
rect 12622 38898 23330 39134
rect 23566 38898 33570 39134
rect 33806 38898 43810 39134
rect 44046 38898 54050 39134
rect 54286 38898 64290 39134
rect 64526 38898 74530 39134
rect 74766 38898 84770 39134
rect 85006 38898 95010 39134
rect 95246 38898 105250 39134
rect 105486 38898 115490 39134
rect 115726 38898 125730 39134
rect 125966 38898 135970 39134
rect 136206 38898 146210 39134
rect 146446 38898 156450 39134
rect 156686 38898 166690 39134
rect 166926 38898 176930 39134
rect 177166 38898 187170 39134
rect 187406 38898 197410 39134
rect 197646 38898 207650 39134
rect 207886 38898 217890 39134
rect 218126 38898 228130 39134
rect 228366 38898 238370 39134
rect 238606 38898 248610 39134
rect 248846 38898 258850 39134
rect 259086 38898 269090 39134
rect 269326 38898 279330 39134
rect 279566 38898 289570 39134
rect 289806 38898 299810 39134
rect 300046 38898 310050 39134
rect 310286 38898 320290 39134
rect 320526 38898 330530 39134
rect 330766 38898 340770 39134
rect 341006 38898 351010 39134
rect 351246 38898 361250 39134
rect 361486 38898 371490 39134
rect 371726 38898 381730 39134
rect 381966 38898 391970 39134
rect 392206 38898 402210 39134
rect 402446 38898 412450 39134
rect 412686 38898 422690 39134
rect 422926 38898 432930 39134
rect 433166 38898 443170 39134
rect 443406 38898 453410 39134
rect 453646 38898 463650 39134
rect 463886 38898 473890 39134
rect 474126 38898 484130 39134
rect 484366 38898 494370 39134
rect 494606 38898 504610 39134
rect 504846 38898 514850 39134
rect 515086 38898 525090 39134
rect 525326 38898 535330 39134
rect 535566 38898 544546 39134
rect 544782 38898 544866 39134
rect 545102 38898 554786 39134
rect 555022 38898 555106 39134
rect 555342 38898 565026 39134
rect 565262 38898 565346 39134
rect 565582 38898 575266 39134
rect 575502 38898 575586 39134
rect 575822 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 550586 32614
rect 550822 32378 550906 32614
rect 551142 32378 560826 32614
rect 561062 32378 561146 32614
rect 561382 32378 571066 32614
rect 571302 32378 571386 32614
rect 571622 32378 581306 32614
rect 581542 32378 581626 32614
rect 581862 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 550586 32294
rect 550822 32058 550906 32294
rect 551142 32058 560826 32294
rect 561062 32058 561146 32294
rect 561382 32058 571066 32294
rect 571302 32058 571386 32294
rect 571622 32058 581306 32294
rect 581542 32058 581626 32294
rect 581862 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 14386 28894
rect 14622 28658 14706 28894
rect 14942 28658 546866 28894
rect 547102 28658 547186 28894
rect 547422 28658 557106 28894
rect 557342 28658 557426 28894
rect 557662 28658 567346 28894
rect 567582 28658 567666 28894
rect 567902 28658 577586 28894
rect 577822 28658 577906 28894
rect 578142 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 14386 28574
rect 14622 28338 14706 28574
rect 14942 28338 546866 28574
rect 547102 28338 547186 28574
rect 547422 28338 557106 28574
rect 557342 28338 557426 28574
rect 557662 28338 567346 28574
rect 567582 28338 567666 28574
rect 567902 28338 577586 28574
rect 577822 28338 577906 28574
rect 578142 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 10666 25174
rect 10902 24938 10986 25174
rect 11222 24938 543146 25174
rect 543382 24938 543466 25174
rect 543702 24938 553386 25174
rect 553622 24938 553706 25174
rect 553942 24938 563626 25174
rect 563862 24938 563946 25174
rect 564182 24938 573866 25174
rect 574102 24938 574186 25174
rect 574422 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 10666 24854
rect 10902 24618 10986 24854
rect 11222 24618 543146 24854
rect 543382 24618 543466 24854
rect 543702 24618 553386 24854
rect 553622 24618 553706 24854
rect 553942 24618 563626 24854
rect 563862 24618 563946 24854
rect 564182 24618 573866 24854
rect 574102 24618 574186 24854
rect 574422 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 6946 21454
rect 7182 21218 7266 21454
rect 7502 21218 28450 21454
rect 28686 21218 38690 21454
rect 38926 21218 48930 21454
rect 49166 21218 59170 21454
rect 59406 21218 69410 21454
rect 69646 21218 79650 21454
rect 79886 21218 89890 21454
rect 90126 21218 100130 21454
rect 100366 21218 110370 21454
rect 110606 21218 120610 21454
rect 120846 21218 130850 21454
rect 131086 21218 141090 21454
rect 141326 21218 151330 21454
rect 151566 21218 161570 21454
rect 161806 21218 171810 21454
rect 172046 21218 182050 21454
rect 182286 21218 192290 21454
rect 192526 21218 202530 21454
rect 202766 21218 212770 21454
rect 213006 21218 223010 21454
rect 223246 21218 233250 21454
rect 233486 21218 243490 21454
rect 243726 21218 253730 21454
rect 253966 21218 263970 21454
rect 264206 21218 274210 21454
rect 274446 21218 284450 21454
rect 284686 21218 294690 21454
rect 294926 21218 304930 21454
rect 305166 21218 315170 21454
rect 315406 21218 325410 21454
rect 325646 21218 335650 21454
rect 335886 21218 345890 21454
rect 346126 21218 356130 21454
rect 356366 21218 366370 21454
rect 366606 21218 376610 21454
rect 376846 21218 386850 21454
rect 387086 21218 397090 21454
rect 397326 21218 407330 21454
rect 407566 21218 417570 21454
rect 417806 21218 427810 21454
rect 428046 21218 438050 21454
rect 438286 21218 448290 21454
rect 448526 21218 458530 21454
rect 458766 21218 468770 21454
rect 469006 21218 479010 21454
rect 479246 21218 489250 21454
rect 489486 21218 499490 21454
rect 499726 21218 509730 21454
rect 509966 21218 519970 21454
rect 520206 21218 530210 21454
rect 530446 21218 549666 21454
rect 549902 21218 549986 21454
rect 550222 21218 559906 21454
rect 560142 21218 560226 21454
rect 560462 21218 570146 21454
rect 570382 21218 570466 21454
rect 570702 21218 580386 21454
rect 580622 21218 580706 21454
rect 580942 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 6946 21134
rect 7182 20898 7266 21134
rect 7502 20898 28450 21134
rect 28686 20898 38690 21134
rect 38926 20898 48930 21134
rect 49166 20898 59170 21134
rect 59406 20898 69410 21134
rect 69646 20898 79650 21134
rect 79886 20898 89890 21134
rect 90126 20898 100130 21134
rect 100366 20898 110370 21134
rect 110606 20898 120610 21134
rect 120846 20898 130850 21134
rect 131086 20898 141090 21134
rect 141326 20898 151330 21134
rect 151566 20898 161570 21134
rect 161806 20898 171810 21134
rect 172046 20898 182050 21134
rect 182286 20898 192290 21134
rect 192526 20898 202530 21134
rect 202766 20898 212770 21134
rect 213006 20898 223010 21134
rect 223246 20898 233250 21134
rect 233486 20898 243490 21134
rect 243726 20898 253730 21134
rect 253966 20898 263970 21134
rect 264206 20898 274210 21134
rect 274446 20898 284450 21134
rect 284686 20898 294690 21134
rect 294926 20898 304930 21134
rect 305166 20898 315170 21134
rect 315406 20898 325410 21134
rect 325646 20898 335650 21134
rect 335886 20898 345890 21134
rect 346126 20898 356130 21134
rect 356366 20898 366370 21134
rect 366606 20898 376610 21134
rect 376846 20898 386850 21134
rect 387086 20898 397090 21134
rect 397326 20898 407330 21134
rect 407566 20898 417570 21134
rect 417806 20898 427810 21134
rect 428046 20898 438050 21134
rect 438286 20898 448290 21134
rect 448526 20898 458530 21134
rect 458766 20898 468770 21134
rect 469006 20898 479010 21134
rect 479246 20898 489250 21134
rect 489486 20898 499490 21134
rect 499726 20898 509730 21134
rect 509966 20898 519970 21134
rect 520206 20898 530210 21134
rect 530446 20898 549666 21134
rect 549902 20898 549986 21134
rect 550222 20898 559906 21134
rect 560142 20898 560226 21134
rect 560462 20898 570146 21134
rect 570382 20898 570466 21134
rect 570702 20898 580386 21134
rect 580622 20898 580706 21134
rect 580942 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 545466 14614
rect 545702 14378 545786 14614
rect 546022 14378 555706 14614
rect 555942 14378 556026 14614
rect 556262 14378 565946 14614
rect 566182 14378 566266 14614
rect 566502 14378 576186 14614
rect 576422 14378 576506 14614
rect 576742 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 545466 14294
rect 545702 14058 545786 14294
rect 546022 14058 555706 14294
rect 555942 14058 556026 14294
rect 556262 14058 565946 14294
rect 566182 14058 566266 14294
rect 566502 14058 576186 14294
rect 576422 14058 576506 14294
rect 576742 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 19506 10894
rect 19742 10658 19826 10894
rect 20062 10658 29746 10894
rect 29982 10658 30066 10894
rect 30302 10658 39986 10894
rect 40222 10658 40306 10894
rect 40542 10658 50226 10894
rect 50462 10658 50546 10894
rect 50782 10658 60466 10894
rect 60702 10658 60786 10894
rect 61022 10658 70706 10894
rect 70942 10658 71026 10894
rect 71262 10658 80946 10894
rect 81182 10658 81266 10894
rect 81502 10658 91186 10894
rect 91422 10658 91506 10894
rect 91742 10658 101426 10894
rect 101662 10658 101746 10894
rect 101982 10658 111666 10894
rect 111902 10658 111986 10894
rect 112222 10658 121906 10894
rect 122142 10658 122226 10894
rect 122462 10658 132146 10894
rect 132382 10658 132466 10894
rect 132702 10658 142386 10894
rect 142622 10658 142706 10894
rect 142942 10658 152626 10894
rect 152862 10658 152946 10894
rect 153182 10658 162866 10894
rect 163102 10658 163186 10894
rect 163422 10658 173106 10894
rect 173342 10658 173426 10894
rect 173662 10658 183346 10894
rect 183582 10658 183666 10894
rect 183902 10658 193586 10894
rect 193822 10658 193906 10894
rect 194142 10658 203826 10894
rect 204062 10658 204146 10894
rect 204382 10658 214066 10894
rect 214302 10658 214386 10894
rect 214622 10658 224306 10894
rect 224542 10658 224626 10894
rect 224862 10658 234546 10894
rect 234782 10658 234866 10894
rect 235102 10658 244786 10894
rect 245022 10658 245106 10894
rect 245342 10658 255026 10894
rect 255262 10658 255346 10894
rect 255582 10658 265266 10894
rect 265502 10658 265586 10894
rect 265822 10658 275506 10894
rect 275742 10658 275826 10894
rect 276062 10658 285746 10894
rect 285982 10658 286066 10894
rect 286302 10658 295986 10894
rect 296222 10658 296306 10894
rect 296542 10658 306226 10894
rect 306462 10658 306546 10894
rect 306782 10658 316466 10894
rect 316702 10658 316786 10894
rect 317022 10658 326706 10894
rect 326942 10658 327026 10894
rect 327262 10658 336946 10894
rect 337182 10658 337266 10894
rect 337502 10658 347186 10894
rect 347422 10658 347506 10894
rect 347742 10658 357426 10894
rect 357662 10658 357746 10894
rect 357982 10658 367666 10894
rect 367902 10658 367986 10894
rect 368222 10658 377906 10894
rect 378142 10658 378226 10894
rect 378462 10658 388146 10894
rect 388382 10658 388466 10894
rect 388702 10658 398386 10894
rect 398622 10658 398706 10894
rect 398942 10658 408626 10894
rect 408862 10658 408946 10894
rect 409182 10658 418866 10894
rect 419102 10658 419186 10894
rect 419422 10658 429106 10894
rect 429342 10658 429426 10894
rect 429662 10658 439346 10894
rect 439582 10658 439666 10894
rect 439902 10658 449586 10894
rect 449822 10658 449906 10894
rect 450142 10658 459826 10894
rect 460062 10658 460146 10894
rect 460382 10658 470066 10894
rect 470302 10658 470386 10894
rect 470622 10658 480306 10894
rect 480542 10658 480626 10894
rect 480862 10658 490546 10894
rect 490782 10658 490866 10894
rect 491102 10658 500786 10894
rect 501022 10658 501106 10894
rect 501342 10658 511026 10894
rect 511262 10658 511346 10894
rect 511582 10658 521266 10894
rect 521502 10658 521586 10894
rect 521822 10658 531506 10894
rect 531742 10658 531826 10894
rect 532062 10658 541746 10894
rect 541982 10658 542066 10894
rect 542302 10658 551986 10894
rect 552222 10658 552306 10894
rect 552542 10658 562226 10894
rect 562462 10658 562546 10894
rect 562782 10658 572466 10894
rect 572702 10658 572786 10894
rect 573022 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 19506 10574
rect 19742 10338 19826 10574
rect 20062 10338 29746 10574
rect 29982 10338 30066 10574
rect 30302 10338 39986 10574
rect 40222 10338 40306 10574
rect 40542 10338 50226 10574
rect 50462 10338 50546 10574
rect 50782 10338 60466 10574
rect 60702 10338 60786 10574
rect 61022 10338 70706 10574
rect 70942 10338 71026 10574
rect 71262 10338 80946 10574
rect 81182 10338 81266 10574
rect 81502 10338 91186 10574
rect 91422 10338 91506 10574
rect 91742 10338 101426 10574
rect 101662 10338 101746 10574
rect 101982 10338 111666 10574
rect 111902 10338 111986 10574
rect 112222 10338 121906 10574
rect 122142 10338 122226 10574
rect 122462 10338 132146 10574
rect 132382 10338 132466 10574
rect 132702 10338 142386 10574
rect 142622 10338 142706 10574
rect 142942 10338 152626 10574
rect 152862 10338 152946 10574
rect 153182 10338 162866 10574
rect 163102 10338 163186 10574
rect 163422 10338 173106 10574
rect 173342 10338 173426 10574
rect 173662 10338 183346 10574
rect 183582 10338 183666 10574
rect 183902 10338 193586 10574
rect 193822 10338 193906 10574
rect 194142 10338 203826 10574
rect 204062 10338 204146 10574
rect 204382 10338 214066 10574
rect 214302 10338 214386 10574
rect 214622 10338 224306 10574
rect 224542 10338 224626 10574
rect 224862 10338 234546 10574
rect 234782 10338 234866 10574
rect 235102 10338 244786 10574
rect 245022 10338 245106 10574
rect 245342 10338 255026 10574
rect 255262 10338 255346 10574
rect 255582 10338 265266 10574
rect 265502 10338 265586 10574
rect 265822 10338 275506 10574
rect 275742 10338 275826 10574
rect 276062 10338 285746 10574
rect 285982 10338 286066 10574
rect 286302 10338 295986 10574
rect 296222 10338 296306 10574
rect 296542 10338 306226 10574
rect 306462 10338 306546 10574
rect 306782 10338 316466 10574
rect 316702 10338 316786 10574
rect 317022 10338 326706 10574
rect 326942 10338 327026 10574
rect 327262 10338 336946 10574
rect 337182 10338 337266 10574
rect 337502 10338 347186 10574
rect 347422 10338 347506 10574
rect 347742 10338 357426 10574
rect 357662 10338 357746 10574
rect 357982 10338 367666 10574
rect 367902 10338 367986 10574
rect 368222 10338 377906 10574
rect 378142 10338 378226 10574
rect 378462 10338 388146 10574
rect 388382 10338 388466 10574
rect 388702 10338 398386 10574
rect 398622 10338 398706 10574
rect 398942 10338 408626 10574
rect 408862 10338 408946 10574
rect 409182 10338 418866 10574
rect 419102 10338 419186 10574
rect 419422 10338 429106 10574
rect 429342 10338 429426 10574
rect 429662 10338 439346 10574
rect 439582 10338 439666 10574
rect 439902 10338 449586 10574
rect 449822 10338 449906 10574
rect 450142 10338 459826 10574
rect 460062 10338 460146 10574
rect 460382 10338 470066 10574
rect 470302 10338 470386 10574
rect 470622 10338 480306 10574
rect 480542 10338 480626 10574
rect 480862 10338 490546 10574
rect 490782 10338 490866 10574
rect 491102 10338 500786 10574
rect 501022 10338 501106 10574
rect 501342 10338 511026 10574
rect 511262 10338 511346 10574
rect 511582 10338 521266 10574
rect 521502 10338 521586 10574
rect 521822 10338 531506 10574
rect 531742 10338 531826 10574
rect 532062 10338 541746 10574
rect 541982 10338 542066 10574
rect 542302 10338 551986 10574
rect 552222 10338 552306 10574
rect 552542 10338 562226 10574
rect 562462 10338 562546 10574
rect 562782 10338 572466 10574
rect 572702 10338 572786 10574
rect 573022 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 15786 7174
rect 16022 6938 16106 7174
rect 16342 6938 26026 7174
rect 26262 6938 26346 7174
rect 26582 6938 36266 7174
rect 36502 6938 36586 7174
rect 36822 6938 46506 7174
rect 46742 6938 46826 7174
rect 47062 6938 56746 7174
rect 56982 6938 57066 7174
rect 57302 6938 66986 7174
rect 67222 6938 67306 7174
rect 67542 6938 77226 7174
rect 77462 6938 77546 7174
rect 77782 6938 87466 7174
rect 87702 6938 87786 7174
rect 88022 6938 97706 7174
rect 97942 6938 98026 7174
rect 98262 6938 107946 7174
rect 108182 6938 108266 7174
rect 108502 6938 118186 7174
rect 118422 6938 118506 7174
rect 118742 6938 128426 7174
rect 128662 6938 128746 7174
rect 128982 6938 138666 7174
rect 138902 6938 138986 7174
rect 139222 6938 148906 7174
rect 149142 6938 149226 7174
rect 149462 6938 159146 7174
rect 159382 6938 159466 7174
rect 159702 6938 169386 7174
rect 169622 6938 169706 7174
rect 169942 6938 179626 7174
rect 179862 6938 179946 7174
rect 180182 6938 189866 7174
rect 190102 6938 190186 7174
rect 190422 6938 200106 7174
rect 200342 6938 200426 7174
rect 200662 6938 210346 7174
rect 210582 6938 210666 7174
rect 210902 6938 220586 7174
rect 220822 6938 220906 7174
rect 221142 6938 230826 7174
rect 231062 6938 231146 7174
rect 231382 6938 241066 7174
rect 241302 6938 241386 7174
rect 241622 6938 251306 7174
rect 251542 6938 251626 7174
rect 251862 6938 261546 7174
rect 261782 6938 261866 7174
rect 262102 6938 271786 7174
rect 272022 6938 272106 7174
rect 272342 6938 282026 7174
rect 282262 6938 282346 7174
rect 282582 6938 292266 7174
rect 292502 6938 292586 7174
rect 292822 6938 302506 7174
rect 302742 6938 302826 7174
rect 303062 6938 312746 7174
rect 312982 6938 313066 7174
rect 313302 6938 322986 7174
rect 323222 6938 323306 7174
rect 323542 6938 333226 7174
rect 333462 6938 333546 7174
rect 333782 6938 343466 7174
rect 343702 6938 343786 7174
rect 344022 6938 353706 7174
rect 353942 6938 354026 7174
rect 354262 6938 363946 7174
rect 364182 6938 364266 7174
rect 364502 6938 374186 7174
rect 374422 6938 374506 7174
rect 374742 6938 384426 7174
rect 384662 6938 384746 7174
rect 384982 6938 394666 7174
rect 394902 6938 394986 7174
rect 395222 6938 404906 7174
rect 405142 6938 405226 7174
rect 405462 6938 415146 7174
rect 415382 6938 415466 7174
rect 415702 6938 425386 7174
rect 425622 6938 425706 7174
rect 425942 6938 435626 7174
rect 435862 6938 435946 7174
rect 436182 6938 445866 7174
rect 446102 6938 446186 7174
rect 446422 6938 456106 7174
rect 456342 6938 456426 7174
rect 456662 6938 466346 7174
rect 466582 6938 466666 7174
rect 466902 6938 476586 7174
rect 476822 6938 476906 7174
rect 477142 6938 486826 7174
rect 487062 6938 487146 7174
rect 487382 6938 497066 7174
rect 497302 6938 497386 7174
rect 497622 6938 507306 7174
rect 507542 6938 507626 7174
rect 507862 6938 517546 7174
rect 517782 6938 517866 7174
rect 518102 6938 527786 7174
rect 528022 6938 528106 7174
rect 528342 6938 538026 7174
rect 538262 6938 538346 7174
rect 538582 6938 548266 7174
rect 548502 6938 548586 7174
rect 548822 6938 558506 7174
rect 558742 6938 558826 7174
rect 559062 6938 568746 7174
rect 568982 6938 569066 7174
rect 569302 6938 578986 7174
rect 579222 6938 579306 7174
rect 579542 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 15786 6854
rect 16022 6618 16106 6854
rect 16342 6618 26026 6854
rect 26262 6618 26346 6854
rect 26582 6618 36266 6854
rect 36502 6618 36586 6854
rect 36822 6618 46506 6854
rect 46742 6618 46826 6854
rect 47062 6618 56746 6854
rect 56982 6618 57066 6854
rect 57302 6618 66986 6854
rect 67222 6618 67306 6854
rect 67542 6618 77226 6854
rect 77462 6618 77546 6854
rect 77782 6618 87466 6854
rect 87702 6618 87786 6854
rect 88022 6618 97706 6854
rect 97942 6618 98026 6854
rect 98262 6618 107946 6854
rect 108182 6618 108266 6854
rect 108502 6618 118186 6854
rect 118422 6618 118506 6854
rect 118742 6618 128426 6854
rect 128662 6618 128746 6854
rect 128982 6618 138666 6854
rect 138902 6618 138986 6854
rect 139222 6618 148906 6854
rect 149142 6618 149226 6854
rect 149462 6618 159146 6854
rect 159382 6618 159466 6854
rect 159702 6618 169386 6854
rect 169622 6618 169706 6854
rect 169942 6618 179626 6854
rect 179862 6618 179946 6854
rect 180182 6618 189866 6854
rect 190102 6618 190186 6854
rect 190422 6618 200106 6854
rect 200342 6618 200426 6854
rect 200662 6618 210346 6854
rect 210582 6618 210666 6854
rect 210902 6618 220586 6854
rect 220822 6618 220906 6854
rect 221142 6618 230826 6854
rect 231062 6618 231146 6854
rect 231382 6618 241066 6854
rect 241302 6618 241386 6854
rect 241622 6618 251306 6854
rect 251542 6618 251626 6854
rect 251862 6618 261546 6854
rect 261782 6618 261866 6854
rect 262102 6618 271786 6854
rect 272022 6618 272106 6854
rect 272342 6618 282026 6854
rect 282262 6618 282346 6854
rect 282582 6618 292266 6854
rect 292502 6618 292586 6854
rect 292822 6618 302506 6854
rect 302742 6618 302826 6854
rect 303062 6618 312746 6854
rect 312982 6618 313066 6854
rect 313302 6618 322986 6854
rect 323222 6618 323306 6854
rect 323542 6618 333226 6854
rect 333462 6618 333546 6854
rect 333782 6618 343466 6854
rect 343702 6618 343786 6854
rect 344022 6618 353706 6854
rect 353942 6618 354026 6854
rect 354262 6618 363946 6854
rect 364182 6618 364266 6854
rect 364502 6618 374186 6854
rect 374422 6618 374506 6854
rect 374742 6618 384426 6854
rect 384662 6618 384746 6854
rect 384982 6618 394666 6854
rect 394902 6618 394986 6854
rect 395222 6618 404906 6854
rect 405142 6618 405226 6854
rect 405462 6618 415146 6854
rect 415382 6618 415466 6854
rect 415702 6618 425386 6854
rect 425622 6618 425706 6854
rect 425942 6618 435626 6854
rect 435862 6618 435946 6854
rect 436182 6618 445866 6854
rect 446102 6618 446186 6854
rect 446422 6618 456106 6854
rect 456342 6618 456426 6854
rect 456662 6618 466346 6854
rect 466582 6618 466666 6854
rect 466902 6618 476586 6854
rect 476822 6618 476906 6854
rect 477142 6618 486826 6854
rect 487062 6618 487146 6854
rect 487382 6618 497066 6854
rect 497302 6618 497386 6854
rect 497622 6618 507306 6854
rect 507542 6618 507626 6854
rect 507862 6618 517546 6854
rect 517782 6618 517866 6854
rect 518102 6618 527786 6854
rect 528022 6618 528106 6854
rect 528342 6618 538026 6854
rect 538262 6618 538346 6854
rect 538582 6618 548266 6854
rect 548502 6618 548586 6854
rect 548822 6618 558506 6854
rect 558742 6618 558826 6854
rect 559062 6618 568746 6854
rect 568982 6618 569066 6854
rect 569302 6618 578986 6854
rect 579222 6618 579306 6854
rect 579542 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 12066 3454
rect 12302 3218 12386 3454
rect 12622 3218 22306 3454
rect 22542 3218 22626 3454
rect 22862 3218 32546 3454
rect 32782 3218 32866 3454
rect 33102 3218 42786 3454
rect 43022 3218 43106 3454
rect 43342 3218 53026 3454
rect 53262 3218 53346 3454
rect 53582 3218 63266 3454
rect 63502 3218 63586 3454
rect 63822 3218 73506 3454
rect 73742 3218 73826 3454
rect 74062 3218 83746 3454
rect 83982 3218 84066 3454
rect 84302 3218 93986 3454
rect 94222 3218 94306 3454
rect 94542 3218 104226 3454
rect 104462 3218 104546 3454
rect 104782 3218 114466 3454
rect 114702 3218 114786 3454
rect 115022 3218 124706 3454
rect 124942 3218 125026 3454
rect 125262 3218 134946 3454
rect 135182 3218 135266 3454
rect 135502 3218 145186 3454
rect 145422 3218 145506 3454
rect 145742 3218 155426 3454
rect 155662 3218 155746 3454
rect 155982 3218 165666 3454
rect 165902 3218 165986 3454
rect 166222 3218 175906 3454
rect 176142 3218 176226 3454
rect 176462 3218 186146 3454
rect 186382 3218 186466 3454
rect 186702 3218 196386 3454
rect 196622 3218 196706 3454
rect 196942 3218 206626 3454
rect 206862 3218 206946 3454
rect 207182 3218 216866 3454
rect 217102 3218 217186 3454
rect 217422 3218 227106 3454
rect 227342 3218 227426 3454
rect 227662 3218 237346 3454
rect 237582 3218 237666 3454
rect 237902 3218 247586 3454
rect 247822 3218 247906 3454
rect 248142 3218 257826 3454
rect 258062 3218 258146 3454
rect 258382 3218 268066 3454
rect 268302 3218 268386 3454
rect 268622 3218 278306 3454
rect 278542 3218 278626 3454
rect 278862 3218 288546 3454
rect 288782 3218 288866 3454
rect 289102 3218 298786 3454
rect 299022 3218 299106 3454
rect 299342 3218 309026 3454
rect 309262 3218 309346 3454
rect 309582 3218 319266 3454
rect 319502 3218 319586 3454
rect 319822 3218 329506 3454
rect 329742 3218 329826 3454
rect 330062 3218 339746 3454
rect 339982 3218 340066 3454
rect 340302 3218 349986 3454
rect 350222 3218 350306 3454
rect 350542 3218 360226 3454
rect 360462 3218 360546 3454
rect 360782 3218 370466 3454
rect 370702 3218 370786 3454
rect 371022 3218 380706 3454
rect 380942 3218 381026 3454
rect 381262 3218 390946 3454
rect 391182 3218 391266 3454
rect 391502 3218 401186 3454
rect 401422 3218 401506 3454
rect 401742 3218 411426 3454
rect 411662 3218 411746 3454
rect 411982 3218 421666 3454
rect 421902 3218 421986 3454
rect 422222 3218 431906 3454
rect 432142 3218 432226 3454
rect 432462 3218 442146 3454
rect 442382 3218 442466 3454
rect 442702 3218 452386 3454
rect 452622 3218 452706 3454
rect 452942 3218 462626 3454
rect 462862 3218 462946 3454
rect 463182 3218 472866 3454
rect 473102 3218 473186 3454
rect 473422 3218 483106 3454
rect 483342 3218 483426 3454
rect 483662 3218 493346 3454
rect 493582 3218 493666 3454
rect 493902 3218 503586 3454
rect 503822 3218 503906 3454
rect 504142 3218 513826 3454
rect 514062 3218 514146 3454
rect 514382 3218 524066 3454
rect 524302 3218 524386 3454
rect 524622 3218 534306 3454
rect 534542 3218 534626 3454
rect 534862 3218 544546 3454
rect 544782 3218 544866 3454
rect 545102 3218 554786 3454
rect 555022 3218 555106 3454
rect 555342 3218 565026 3454
rect 565262 3218 565346 3454
rect 565582 3218 575266 3454
rect 575502 3218 575586 3454
rect 575822 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 12066 3134
rect 12302 2898 12386 3134
rect 12622 2898 22306 3134
rect 22542 2898 22626 3134
rect 22862 2898 32546 3134
rect 32782 2898 32866 3134
rect 33102 2898 42786 3134
rect 43022 2898 43106 3134
rect 43342 2898 53026 3134
rect 53262 2898 53346 3134
rect 53582 2898 63266 3134
rect 63502 2898 63586 3134
rect 63822 2898 73506 3134
rect 73742 2898 73826 3134
rect 74062 2898 83746 3134
rect 83982 2898 84066 3134
rect 84302 2898 93986 3134
rect 94222 2898 94306 3134
rect 94542 2898 104226 3134
rect 104462 2898 104546 3134
rect 104782 2898 114466 3134
rect 114702 2898 114786 3134
rect 115022 2898 124706 3134
rect 124942 2898 125026 3134
rect 125262 2898 134946 3134
rect 135182 2898 135266 3134
rect 135502 2898 145186 3134
rect 145422 2898 145506 3134
rect 145742 2898 155426 3134
rect 155662 2898 155746 3134
rect 155982 2898 165666 3134
rect 165902 2898 165986 3134
rect 166222 2898 175906 3134
rect 176142 2898 176226 3134
rect 176462 2898 186146 3134
rect 186382 2898 186466 3134
rect 186702 2898 196386 3134
rect 196622 2898 196706 3134
rect 196942 2898 206626 3134
rect 206862 2898 206946 3134
rect 207182 2898 216866 3134
rect 217102 2898 217186 3134
rect 217422 2898 227106 3134
rect 227342 2898 227426 3134
rect 227662 2898 237346 3134
rect 237582 2898 237666 3134
rect 237902 2898 247586 3134
rect 247822 2898 247906 3134
rect 248142 2898 257826 3134
rect 258062 2898 258146 3134
rect 258382 2898 268066 3134
rect 268302 2898 268386 3134
rect 268622 2898 278306 3134
rect 278542 2898 278626 3134
rect 278862 2898 288546 3134
rect 288782 2898 288866 3134
rect 289102 2898 298786 3134
rect 299022 2898 299106 3134
rect 299342 2898 309026 3134
rect 309262 2898 309346 3134
rect 309582 2898 319266 3134
rect 319502 2898 319586 3134
rect 319822 2898 329506 3134
rect 329742 2898 329826 3134
rect 330062 2898 339746 3134
rect 339982 2898 340066 3134
rect 340302 2898 349986 3134
rect 350222 2898 350306 3134
rect 350542 2898 360226 3134
rect 360462 2898 360546 3134
rect 360782 2898 370466 3134
rect 370702 2898 370786 3134
rect 371022 2898 380706 3134
rect 380942 2898 381026 3134
rect 381262 2898 390946 3134
rect 391182 2898 391266 3134
rect 391502 2898 401186 3134
rect 401422 2898 401506 3134
rect 401742 2898 411426 3134
rect 411662 2898 411746 3134
rect 411982 2898 421666 3134
rect 421902 2898 421986 3134
rect 422222 2898 431906 3134
rect 432142 2898 432226 3134
rect 432462 2898 442146 3134
rect 442382 2898 442466 3134
rect 442702 2898 452386 3134
rect 452622 2898 452706 3134
rect 452942 2898 462626 3134
rect 462862 2898 462946 3134
rect 463182 2898 472866 3134
rect 473102 2898 473186 3134
rect 473422 2898 483106 3134
rect 483342 2898 483426 3134
rect 483662 2898 493346 3134
rect 493582 2898 493666 3134
rect 493902 2898 503586 3134
rect 503822 2898 503906 3134
rect 504142 2898 513826 3134
rect 514062 2898 514146 3134
rect 514382 2898 524066 3134
rect 524302 2898 524386 3134
rect 524622 2898 534306 3134
rect 534542 2898 534626 3134
rect 534862 2898 544546 3134
rect 544782 2898 544866 3134
rect 545102 2898 554786 3134
rect 555022 2898 555106 3134
rect 555342 2898 565026 3134
rect 565262 2898 565346 3134
rect 565582 2898 575266 3134
rect 575502 2898 575586 3134
rect 575822 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 12066 -346
rect 12302 -582 12386 -346
rect 12622 -582 22306 -346
rect 22542 -582 22626 -346
rect 22862 -582 32546 -346
rect 32782 -582 32866 -346
rect 33102 -582 42786 -346
rect 43022 -582 43106 -346
rect 43342 -582 53026 -346
rect 53262 -582 53346 -346
rect 53582 -582 63266 -346
rect 63502 -582 63586 -346
rect 63822 -582 73506 -346
rect 73742 -582 73826 -346
rect 74062 -582 83746 -346
rect 83982 -582 84066 -346
rect 84302 -582 93986 -346
rect 94222 -582 94306 -346
rect 94542 -582 104226 -346
rect 104462 -582 104546 -346
rect 104782 -582 114466 -346
rect 114702 -582 114786 -346
rect 115022 -582 124706 -346
rect 124942 -582 125026 -346
rect 125262 -582 134946 -346
rect 135182 -582 135266 -346
rect 135502 -582 145186 -346
rect 145422 -582 145506 -346
rect 145742 -582 155426 -346
rect 155662 -582 155746 -346
rect 155982 -582 165666 -346
rect 165902 -582 165986 -346
rect 166222 -582 175906 -346
rect 176142 -582 176226 -346
rect 176462 -582 186146 -346
rect 186382 -582 186466 -346
rect 186702 -582 196386 -346
rect 196622 -582 196706 -346
rect 196942 -582 206626 -346
rect 206862 -582 206946 -346
rect 207182 -582 216866 -346
rect 217102 -582 217186 -346
rect 217422 -582 227106 -346
rect 227342 -582 227426 -346
rect 227662 -582 237346 -346
rect 237582 -582 237666 -346
rect 237902 -582 247586 -346
rect 247822 -582 247906 -346
rect 248142 -582 257826 -346
rect 258062 -582 258146 -346
rect 258382 -582 268066 -346
rect 268302 -582 268386 -346
rect 268622 -582 278306 -346
rect 278542 -582 278626 -346
rect 278862 -582 288546 -346
rect 288782 -582 288866 -346
rect 289102 -582 298786 -346
rect 299022 -582 299106 -346
rect 299342 -582 309026 -346
rect 309262 -582 309346 -346
rect 309582 -582 319266 -346
rect 319502 -582 319586 -346
rect 319822 -582 329506 -346
rect 329742 -582 329826 -346
rect 330062 -582 339746 -346
rect 339982 -582 340066 -346
rect 340302 -582 349986 -346
rect 350222 -582 350306 -346
rect 350542 -582 360226 -346
rect 360462 -582 360546 -346
rect 360782 -582 370466 -346
rect 370702 -582 370786 -346
rect 371022 -582 380706 -346
rect 380942 -582 381026 -346
rect 381262 -582 390946 -346
rect 391182 -582 391266 -346
rect 391502 -582 401186 -346
rect 401422 -582 401506 -346
rect 401742 -582 411426 -346
rect 411662 -582 411746 -346
rect 411982 -582 421666 -346
rect 421902 -582 421986 -346
rect 422222 -582 431906 -346
rect 432142 -582 432226 -346
rect 432462 -582 442146 -346
rect 442382 -582 442466 -346
rect 442702 -582 452386 -346
rect 452622 -582 452706 -346
rect 452942 -582 462626 -346
rect 462862 -582 462946 -346
rect 463182 -582 472866 -346
rect 473102 -582 473186 -346
rect 473422 -582 483106 -346
rect 483342 -582 483426 -346
rect 483662 -582 493346 -346
rect 493582 -582 493666 -346
rect 493902 -582 503586 -346
rect 503822 -582 503906 -346
rect 504142 -582 513826 -346
rect 514062 -582 514146 -346
rect 514382 -582 524066 -346
rect 524302 -582 524386 -346
rect 524622 -582 534306 -346
rect 534542 -582 534626 -346
rect 534862 -582 544546 -346
rect 544782 -582 544866 -346
rect 545102 -582 554786 -346
rect 555022 -582 555106 -346
rect 555342 -582 565026 -346
rect 565262 -582 565346 -346
rect 565582 -582 575266 -346
rect 575502 -582 575586 -346
rect 575822 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 12066 -666
rect 12302 -902 12386 -666
rect 12622 -902 22306 -666
rect 22542 -902 22626 -666
rect 22862 -902 32546 -666
rect 32782 -902 32866 -666
rect 33102 -902 42786 -666
rect 43022 -902 43106 -666
rect 43342 -902 53026 -666
rect 53262 -902 53346 -666
rect 53582 -902 63266 -666
rect 63502 -902 63586 -666
rect 63822 -902 73506 -666
rect 73742 -902 73826 -666
rect 74062 -902 83746 -666
rect 83982 -902 84066 -666
rect 84302 -902 93986 -666
rect 94222 -902 94306 -666
rect 94542 -902 104226 -666
rect 104462 -902 104546 -666
rect 104782 -902 114466 -666
rect 114702 -902 114786 -666
rect 115022 -902 124706 -666
rect 124942 -902 125026 -666
rect 125262 -902 134946 -666
rect 135182 -902 135266 -666
rect 135502 -902 145186 -666
rect 145422 -902 145506 -666
rect 145742 -902 155426 -666
rect 155662 -902 155746 -666
rect 155982 -902 165666 -666
rect 165902 -902 165986 -666
rect 166222 -902 175906 -666
rect 176142 -902 176226 -666
rect 176462 -902 186146 -666
rect 186382 -902 186466 -666
rect 186702 -902 196386 -666
rect 196622 -902 196706 -666
rect 196942 -902 206626 -666
rect 206862 -902 206946 -666
rect 207182 -902 216866 -666
rect 217102 -902 217186 -666
rect 217422 -902 227106 -666
rect 227342 -902 227426 -666
rect 227662 -902 237346 -666
rect 237582 -902 237666 -666
rect 237902 -902 247586 -666
rect 247822 -902 247906 -666
rect 248142 -902 257826 -666
rect 258062 -902 258146 -666
rect 258382 -902 268066 -666
rect 268302 -902 268386 -666
rect 268622 -902 278306 -666
rect 278542 -902 278626 -666
rect 278862 -902 288546 -666
rect 288782 -902 288866 -666
rect 289102 -902 298786 -666
rect 299022 -902 299106 -666
rect 299342 -902 309026 -666
rect 309262 -902 309346 -666
rect 309582 -902 319266 -666
rect 319502 -902 319586 -666
rect 319822 -902 329506 -666
rect 329742 -902 329826 -666
rect 330062 -902 339746 -666
rect 339982 -902 340066 -666
rect 340302 -902 349986 -666
rect 350222 -902 350306 -666
rect 350542 -902 360226 -666
rect 360462 -902 360546 -666
rect 360782 -902 370466 -666
rect 370702 -902 370786 -666
rect 371022 -902 380706 -666
rect 380942 -902 381026 -666
rect 381262 -902 390946 -666
rect 391182 -902 391266 -666
rect 391502 -902 401186 -666
rect 401422 -902 401506 -666
rect 401742 -902 411426 -666
rect 411662 -902 411746 -666
rect 411982 -902 421666 -666
rect 421902 -902 421986 -666
rect 422222 -902 431906 -666
rect 432142 -902 432226 -666
rect 432462 -902 442146 -666
rect 442382 -902 442466 -666
rect 442702 -902 452386 -666
rect 452622 -902 452706 -666
rect 452942 -902 462626 -666
rect 462862 -902 462946 -666
rect 463182 -902 472866 -666
rect 473102 -902 473186 -666
rect 473422 -902 483106 -666
rect 483342 -902 483426 -666
rect 483662 -902 493346 -666
rect 493582 -902 493666 -666
rect 493902 -902 503586 -666
rect 503822 -902 503906 -666
rect 504142 -902 513826 -666
rect 514062 -902 514146 -666
rect 514382 -902 524066 -666
rect 524302 -902 524386 -666
rect 524622 -902 534306 -666
rect 534542 -902 534626 -666
rect 534862 -902 544546 -666
rect 544782 -902 544866 -666
rect 545102 -902 554786 -666
rect 555022 -902 555106 -666
rect 555342 -902 565026 -666
rect 565262 -902 565346 -666
rect 565582 -902 575266 -666
rect 575502 -902 575586 -666
rect 575822 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6946 -1306
rect 7182 -1542 7266 -1306
rect 7502 -1542 17186 -1306
rect 17422 -1542 17506 -1306
rect 17742 -1542 27426 -1306
rect 27662 -1542 27746 -1306
rect 27982 -1542 37666 -1306
rect 37902 -1542 37986 -1306
rect 38222 -1542 47906 -1306
rect 48142 -1542 48226 -1306
rect 48462 -1542 58146 -1306
rect 58382 -1542 58466 -1306
rect 58702 -1542 68386 -1306
rect 68622 -1542 68706 -1306
rect 68942 -1542 78626 -1306
rect 78862 -1542 78946 -1306
rect 79182 -1542 88866 -1306
rect 89102 -1542 89186 -1306
rect 89422 -1542 99106 -1306
rect 99342 -1542 99426 -1306
rect 99662 -1542 109346 -1306
rect 109582 -1542 109666 -1306
rect 109902 -1542 119586 -1306
rect 119822 -1542 119906 -1306
rect 120142 -1542 129826 -1306
rect 130062 -1542 130146 -1306
rect 130382 -1542 140066 -1306
rect 140302 -1542 140386 -1306
rect 140622 -1542 150306 -1306
rect 150542 -1542 150626 -1306
rect 150862 -1542 160546 -1306
rect 160782 -1542 160866 -1306
rect 161102 -1542 170786 -1306
rect 171022 -1542 171106 -1306
rect 171342 -1542 181026 -1306
rect 181262 -1542 181346 -1306
rect 181582 -1542 191266 -1306
rect 191502 -1542 191586 -1306
rect 191822 -1542 201506 -1306
rect 201742 -1542 201826 -1306
rect 202062 -1542 211746 -1306
rect 211982 -1542 212066 -1306
rect 212302 -1542 221986 -1306
rect 222222 -1542 222306 -1306
rect 222542 -1542 232226 -1306
rect 232462 -1542 232546 -1306
rect 232782 -1542 242466 -1306
rect 242702 -1542 242786 -1306
rect 243022 -1542 252706 -1306
rect 252942 -1542 253026 -1306
rect 253262 -1542 262946 -1306
rect 263182 -1542 263266 -1306
rect 263502 -1542 273186 -1306
rect 273422 -1542 273506 -1306
rect 273742 -1542 283426 -1306
rect 283662 -1542 283746 -1306
rect 283982 -1542 293666 -1306
rect 293902 -1542 293986 -1306
rect 294222 -1542 303906 -1306
rect 304142 -1542 304226 -1306
rect 304462 -1542 314146 -1306
rect 314382 -1542 314466 -1306
rect 314702 -1542 324386 -1306
rect 324622 -1542 324706 -1306
rect 324942 -1542 334626 -1306
rect 334862 -1542 334946 -1306
rect 335182 -1542 344866 -1306
rect 345102 -1542 345186 -1306
rect 345422 -1542 355106 -1306
rect 355342 -1542 355426 -1306
rect 355662 -1542 365346 -1306
rect 365582 -1542 365666 -1306
rect 365902 -1542 375586 -1306
rect 375822 -1542 375906 -1306
rect 376142 -1542 385826 -1306
rect 386062 -1542 386146 -1306
rect 386382 -1542 396066 -1306
rect 396302 -1542 396386 -1306
rect 396622 -1542 406306 -1306
rect 406542 -1542 406626 -1306
rect 406862 -1542 416546 -1306
rect 416782 -1542 416866 -1306
rect 417102 -1542 426786 -1306
rect 427022 -1542 427106 -1306
rect 427342 -1542 437026 -1306
rect 437262 -1542 437346 -1306
rect 437582 -1542 447266 -1306
rect 447502 -1542 447586 -1306
rect 447822 -1542 457506 -1306
rect 457742 -1542 457826 -1306
rect 458062 -1542 467746 -1306
rect 467982 -1542 468066 -1306
rect 468302 -1542 477986 -1306
rect 478222 -1542 478306 -1306
rect 478542 -1542 488226 -1306
rect 488462 -1542 488546 -1306
rect 488782 -1542 498466 -1306
rect 498702 -1542 498786 -1306
rect 499022 -1542 508706 -1306
rect 508942 -1542 509026 -1306
rect 509262 -1542 518946 -1306
rect 519182 -1542 519266 -1306
rect 519502 -1542 529186 -1306
rect 529422 -1542 529506 -1306
rect 529742 -1542 539426 -1306
rect 539662 -1542 539746 -1306
rect 539982 -1542 549666 -1306
rect 549902 -1542 549986 -1306
rect 550222 -1542 559906 -1306
rect 560142 -1542 560226 -1306
rect 560462 -1542 570146 -1306
rect 570382 -1542 570466 -1306
rect 570702 -1542 580386 -1306
rect 580622 -1542 580706 -1306
rect 580942 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6946 -1626
rect 7182 -1862 7266 -1626
rect 7502 -1862 17186 -1626
rect 17422 -1862 17506 -1626
rect 17742 -1862 27426 -1626
rect 27662 -1862 27746 -1626
rect 27982 -1862 37666 -1626
rect 37902 -1862 37986 -1626
rect 38222 -1862 47906 -1626
rect 48142 -1862 48226 -1626
rect 48462 -1862 58146 -1626
rect 58382 -1862 58466 -1626
rect 58702 -1862 68386 -1626
rect 68622 -1862 68706 -1626
rect 68942 -1862 78626 -1626
rect 78862 -1862 78946 -1626
rect 79182 -1862 88866 -1626
rect 89102 -1862 89186 -1626
rect 89422 -1862 99106 -1626
rect 99342 -1862 99426 -1626
rect 99662 -1862 109346 -1626
rect 109582 -1862 109666 -1626
rect 109902 -1862 119586 -1626
rect 119822 -1862 119906 -1626
rect 120142 -1862 129826 -1626
rect 130062 -1862 130146 -1626
rect 130382 -1862 140066 -1626
rect 140302 -1862 140386 -1626
rect 140622 -1862 150306 -1626
rect 150542 -1862 150626 -1626
rect 150862 -1862 160546 -1626
rect 160782 -1862 160866 -1626
rect 161102 -1862 170786 -1626
rect 171022 -1862 171106 -1626
rect 171342 -1862 181026 -1626
rect 181262 -1862 181346 -1626
rect 181582 -1862 191266 -1626
rect 191502 -1862 191586 -1626
rect 191822 -1862 201506 -1626
rect 201742 -1862 201826 -1626
rect 202062 -1862 211746 -1626
rect 211982 -1862 212066 -1626
rect 212302 -1862 221986 -1626
rect 222222 -1862 222306 -1626
rect 222542 -1862 232226 -1626
rect 232462 -1862 232546 -1626
rect 232782 -1862 242466 -1626
rect 242702 -1862 242786 -1626
rect 243022 -1862 252706 -1626
rect 252942 -1862 253026 -1626
rect 253262 -1862 262946 -1626
rect 263182 -1862 263266 -1626
rect 263502 -1862 273186 -1626
rect 273422 -1862 273506 -1626
rect 273742 -1862 283426 -1626
rect 283662 -1862 283746 -1626
rect 283982 -1862 293666 -1626
rect 293902 -1862 293986 -1626
rect 294222 -1862 303906 -1626
rect 304142 -1862 304226 -1626
rect 304462 -1862 314146 -1626
rect 314382 -1862 314466 -1626
rect 314702 -1862 324386 -1626
rect 324622 -1862 324706 -1626
rect 324942 -1862 334626 -1626
rect 334862 -1862 334946 -1626
rect 335182 -1862 344866 -1626
rect 345102 -1862 345186 -1626
rect 345422 -1862 355106 -1626
rect 355342 -1862 355426 -1626
rect 355662 -1862 365346 -1626
rect 365582 -1862 365666 -1626
rect 365902 -1862 375586 -1626
rect 375822 -1862 375906 -1626
rect 376142 -1862 385826 -1626
rect 386062 -1862 386146 -1626
rect 386382 -1862 396066 -1626
rect 396302 -1862 396386 -1626
rect 396622 -1862 406306 -1626
rect 406542 -1862 406626 -1626
rect 406862 -1862 416546 -1626
rect 416782 -1862 416866 -1626
rect 417102 -1862 426786 -1626
rect 427022 -1862 427106 -1626
rect 427342 -1862 437026 -1626
rect 437262 -1862 437346 -1626
rect 437582 -1862 447266 -1626
rect 447502 -1862 447586 -1626
rect 447822 -1862 457506 -1626
rect 457742 -1862 457826 -1626
rect 458062 -1862 467746 -1626
rect 467982 -1862 468066 -1626
rect 468302 -1862 477986 -1626
rect 478222 -1862 478306 -1626
rect 478542 -1862 488226 -1626
rect 488462 -1862 488546 -1626
rect 488782 -1862 498466 -1626
rect 498702 -1862 498786 -1626
rect 499022 -1862 508706 -1626
rect 508942 -1862 509026 -1626
rect 509262 -1862 518946 -1626
rect 519182 -1862 519266 -1626
rect 519502 -1862 529186 -1626
rect 529422 -1862 529506 -1626
rect 529742 -1862 539426 -1626
rect 539662 -1862 539746 -1626
rect 539982 -1862 549666 -1626
rect 549902 -1862 549986 -1626
rect 550222 -1862 559906 -1626
rect 560142 -1862 560226 -1626
rect 560462 -1862 570146 -1626
rect 570382 -1862 570466 -1626
rect 570702 -1862 580386 -1626
rect 580622 -1862 580706 -1626
rect 580942 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 15786 -2266
rect 16022 -2502 16106 -2266
rect 16342 -2502 26026 -2266
rect 26262 -2502 26346 -2266
rect 26582 -2502 36266 -2266
rect 36502 -2502 36586 -2266
rect 36822 -2502 46506 -2266
rect 46742 -2502 46826 -2266
rect 47062 -2502 56746 -2266
rect 56982 -2502 57066 -2266
rect 57302 -2502 66986 -2266
rect 67222 -2502 67306 -2266
rect 67542 -2502 77226 -2266
rect 77462 -2502 77546 -2266
rect 77782 -2502 87466 -2266
rect 87702 -2502 87786 -2266
rect 88022 -2502 97706 -2266
rect 97942 -2502 98026 -2266
rect 98262 -2502 107946 -2266
rect 108182 -2502 108266 -2266
rect 108502 -2502 118186 -2266
rect 118422 -2502 118506 -2266
rect 118742 -2502 128426 -2266
rect 128662 -2502 128746 -2266
rect 128982 -2502 138666 -2266
rect 138902 -2502 138986 -2266
rect 139222 -2502 148906 -2266
rect 149142 -2502 149226 -2266
rect 149462 -2502 159146 -2266
rect 159382 -2502 159466 -2266
rect 159702 -2502 169386 -2266
rect 169622 -2502 169706 -2266
rect 169942 -2502 179626 -2266
rect 179862 -2502 179946 -2266
rect 180182 -2502 189866 -2266
rect 190102 -2502 190186 -2266
rect 190422 -2502 200106 -2266
rect 200342 -2502 200426 -2266
rect 200662 -2502 210346 -2266
rect 210582 -2502 210666 -2266
rect 210902 -2502 220586 -2266
rect 220822 -2502 220906 -2266
rect 221142 -2502 230826 -2266
rect 231062 -2502 231146 -2266
rect 231382 -2502 241066 -2266
rect 241302 -2502 241386 -2266
rect 241622 -2502 251306 -2266
rect 251542 -2502 251626 -2266
rect 251862 -2502 261546 -2266
rect 261782 -2502 261866 -2266
rect 262102 -2502 271786 -2266
rect 272022 -2502 272106 -2266
rect 272342 -2502 282026 -2266
rect 282262 -2502 282346 -2266
rect 282582 -2502 292266 -2266
rect 292502 -2502 292586 -2266
rect 292822 -2502 302506 -2266
rect 302742 -2502 302826 -2266
rect 303062 -2502 312746 -2266
rect 312982 -2502 313066 -2266
rect 313302 -2502 322986 -2266
rect 323222 -2502 323306 -2266
rect 323542 -2502 333226 -2266
rect 333462 -2502 333546 -2266
rect 333782 -2502 343466 -2266
rect 343702 -2502 343786 -2266
rect 344022 -2502 353706 -2266
rect 353942 -2502 354026 -2266
rect 354262 -2502 363946 -2266
rect 364182 -2502 364266 -2266
rect 364502 -2502 374186 -2266
rect 374422 -2502 374506 -2266
rect 374742 -2502 384426 -2266
rect 384662 -2502 384746 -2266
rect 384982 -2502 394666 -2266
rect 394902 -2502 394986 -2266
rect 395222 -2502 404906 -2266
rect 405142 -2502 405226 -2266
rect 405462 -2502 415146 -2266
rect 415382 -2502 415466 -2266
rect 415702 -2502 425386 -2266
rect 425622 -2502 425706 -2266
rect 425942 -2502 435626 -2266
rect 435862 -2502 435946 -2266
rect 436182 -2502 445866 -2266
rect 446102 -2502 446186 -2266
rect 446422 -2502 456106 -2266
rect 456342 -2502 456426 -2266
rect 456662 -2502 466346 -2266
rect 466582 -2502 466666 -2266
rect 466902 -2502 476586 -2266
rect 476822 -2502 476906 -2266
rect 477142 -2502 486826 -2266
rect 487062 -2502 487146 -2266
rect 487382 -2502 497066 -2266
rect 497302 -2502 497386 -2266
rect 497622 -2502 507306 -2266
rect 507542 -2502 507626 -2266
rect 507862 -2502 517546 -2266
rect 517782 -2502 517866 -2266
rect 518102 -2502 527786 -2266
rect 528022 -2502 528106 -2266
rect 528342 -2502 538026 -2266
rect 538262 -2502 538346 -2266
rect 538582 -2502 548266 -2266
rect 548502 -2502 548586 -2266
rect 548822 -2502 558506 -2266
rect 558742 -2502 558826 -2266
rect 559062 -2502 568746 -2266
rect 568982 -2502 569066 -2266
rect 569302 -2502 578986 -2266
rect 579222 -2502 579306 -2266
rect 579542 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 15786 -2586
rect 16022 -2822 16106 -2586
rect 16342 -2822 26026 -2586
rect 26262 -2822 26346 -2586
rect 26582 -2822 36266 -2586
rect 36502 -2822 36586 -2586
rect 36822 -2822 46506 -2586
rect 46742 -2822 46826 -2586
rect 47062 -2822 56746 -2586
rect 56982 -2822 57066 -2586
rect 57302 -2822 66986 -2586
rect 67222 -2822 67306 -2586
rect 67542 -2822 77226 -2586
rect 77462 -2822 77546 -2586
rect 77782 -2822 87466 -2586
rect 87702 -2822 87786 -2586
rect 88022 -2822 97706 -2586
rect 97942 -2822 98026 -2586
rect 98262 -2822 107946 -2586
rect 108182 -2822 108266 -2586
rect 108502 -2822 118186 -2586
rect 118422 -2822 118506 -2586
rect 118742 -2822 128426 -2586
rect 128662 -2822 128746 -2586
rect 128982 -2822 138666 -2586
rect 138902 -2822 138986 -2586
rect 139222 -2822 148906 -2586
rect 149142 -2822 149226 -2586
rect 149462 -2822 159146 -2586
rect 159382 -2822 159466 -2586
rect 159702 -2822 169386 -2586
rect 169622 -2822 169706 -2586
rect 169942 -2822 179626 -2586
rect 179862 -2822 179946 -2586
rect 180182 -2822 189866 -2586
rect 190102 -2822 190186 -2586
rect 190422 -2822 200106 -2586
rect 200342 -2822 200426 -2586
rect 200662 -2822 210346 -2586
rect 210582 -2822 210666 -2586
rect 210902 -2822 220586 -2586
rect 220822 -2822 220906 -2586
rect 221142 -2822 230826 -2586
rect 231062 -2822 231146 -2586
rect 231382 -2822 241066 -2586
rect 241302 -2822 241386 -2586
rect 241622 -2822 251306 -2586
rect 251542 -2822 251626 -2586
rect 251862 -2822 261546 -2586
rect 261782 -2822 261866 -2586
rect 262102 -2822 271786 -2586
rect 272022 -2822 272106 -2586
rect 272342 -2822 282026 -2586
rect 282262 -2822 282346 -2586
rect 282582 -2822 292266 -2586
rect 292502 -2822 292586 -2586
rect 292822 -2822 302506 -2586
rect 302742 -2822 302826 -2586
rect 303062 -2822 312746 -2586
rect 312982 -2822 313066 -2586
rect 313302 -2822 322986 -2586
rect 323222 -2822 323306 -2586
rect 323542 -2822 333226 -2586
rect 333462 -2822 333546 -2586
rect 333782 -2822 343466 -2586
rect 343702 -2822 343786 -2586
rect 344022 -2822 353706 -2586
rect 353942 -2822 354026 -2586
rect 354262 -2822 363946 -2586
rect 364182 -2822 364266 -2586
rect 364502 -2822 374186 -2586
rect 374422 -2822 374506 -2586
rect 374742 -2822 384426 -2586
rect 384662 -2822 384746 -2586
rect 384982 -2822 394666 -2586
rect 394902 -2822 394986 -2586
rect 395222 -2822 404906 -2586
rect 405142 -2822 405226 -2586
rect 405462 -2822 415146 -2586
rect 415382 -2822 415466 -2586
rect 415702 -2822 425386 -2586
rect 425622 -2822 425706 -2586
rect 425942 -2822 435626 -2586
rect 435862 -2822 435946 -2586
rect 436182 -2822 445866 -2586
rect 446102 -2822 446186 -2586
rect 446422 -2822 456106 -2586
rect 456342 -2822 456426 -2586
rect 456662 -2822 466346 -2586
rect 466582 -2822 466666 -2586
rect 466902 -2822 476586 -2586
rect 476822 -2822 476906 -2586
rect 477142 -2822 486826 -2586
rect 487062 -2822 487146 -2586
rect 487382 -2822 497066 -2586
rect 497302 -2822 497386 -2586
rect 497622 -2822 507306 -2586
rect 507542 -2822 507626 -2586
rect 507862 -2822 517546 -2586
rect 517782 -2822 517866 -2586
rect 518102 -2822 527786 -2586
rect 528022 -2822 528106 -2586
rect 528342 -2822 538026 -2586
rect 538262 -2822 538346 -2586
rect 538582 -2822 548266 -2586
rect 548502 -2822 548586 -2586
rect 548822 -2822 558506 -2586
rect 558742 -2822 558826 -2586
rect 559062 -2822 568746 -2586
rect 568982 -2822 569066 -2586
rect 569302 -2822 578986 -2586
rect 579222 -2822 579306 -2586
rect 579542 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 10666 -3226
rect 10902 -3462 10986 -3226
rect 11222 -3462 20906 -3226
rect 21142 -3462 21226 -3226
rect 21462 -3462 31146 -3226
rect 31382 -3462 31466 -3226
rect 31702 -3462 41386 -3226
rect 41622 -3462 41706 -3226
rect 41942 -3462 51626 -3226
rect 51862 -3462 51946 -3226
rect 52182 -3462 61866 -3226
rect 62102 -3462 62186 -3226
rect 62422 -3462 72106 -3226
rect 72342 -3462 72426 -3226
rect 72662 -3462 82346 -3226
rect 82582 -3462 82666 -3226
rect 82902 -3462 92586 -3226
rect 92822 -3462 92906 -3226
rect 93142 -3462 102826 -3226
rect 103062 -3462 103146 -3226
rect 103382 -3462 113066 -3226
rect 113302 -3462 113386 -3226
rect 113622 -3462 123306 -3226
rect 123542 -3462 123626 -3226
rect 123862 -3462 133546 -3226
rect 133782 -3462 133866 -3226
rect 134102 -3462 143786 -3226
rect 144022 -3462 144106 -3226
rect 144342 -3462 154026 -3226
rect 154262 -3462 154346 -3226
rect 154582 -3462 164266 -3226
rect 164502 -3462 164586 -3226
rect 164822 -3462 174506 -3226
rect 174742 -3462 174826 -3226
rect 175062 -3462 184746 -3226
rect 184982 -3462 185066 -3226
rect 185302 -3462 194986 -3226
rect 195222 -3462 195306 -3226
rect 195542 -3462 205226 -3226
rect 205462 -3462 205546 -3226
rect 205782 -3462 215466 -3226
rect 215702 -3462 215786 -3226
rect 216022 -3462 225706 -3226
rect 225942 -3462 226026 -3226
rect 226262 -3462 235946 -3226
rect 236182 -3462 236266 -3226
rect 236502 -3462 246186 -3226
rect 246422 -3462 246506 -3226
rect 246742 -3462 256426 -3226
rect 256662 -3462 256746 -3226
rect 256982 -3462 266666 -3226
rect 266902 -3462 266986 -3226
rect 267222 -3462 276906 -3226
rect 277142 -3462 277226 -3226
rect 277462 -3462 287146 -3226
rect 287382 -3462 287466 -3226
rect 287702 -3462 297386 -3226
rect 297622 -3462 297706 -3226
rect 297942 -3462 307626 -3226
rect 307862 -3462 307946 -3226
rect 308182 -3462 317866 -3226
rect 318102 -3462 318186 -3226
rect 318422 -3462 328106 -3226
rect 328342 -3462 328426 -3226
rect 328662 -3462 338346 -3226
rect 338582 -3462 338666 -3226
rect 338902 -3462 348586 -3226
rect 348822 -3462 348906 -3226
rect 349142 -3462 358826 -3226
rect 359062 -3462 359146 -3226
rect 359382 -3462 369066 -3226
rect 369302 -3462 369386 -3226
rect 369622 -3462 379306 -3226
rect 379542 -3462 379626 -3226
rect 379862 -3462 389546 -3226
rect 389782 -3462 389866 -3226
rect 390102 -3462 399786 -3226
rect 400022 -3462 400106 -3226
rect 400342 -3462 410026 -3226
rect 410262 -3462 410346 -3226
rect 410582 -3462 420266 -3226
rect 420502 -3462 420586 -3226
rect 420822 -3462 430506 -3226
rect 430742 -3462 430826 -3226
rect 431062 -3462 440746 -3226
rect 440982 -3462 441066 -3226
rect 441302 -3462 450986 -3226
rect 451222 -3462 451306 -3226
rect 451542 -3462 461226 -3226
rect 461462 -3462 461546 -3226
rect 461782 -3462 471466 -3226
rect 471702 -3462 471786 -3226
rect 472022 -3462 481706 -3226
rect 481942 -3462 482026 -3226
rect 482262 -3462 491946 -3226
rect 492182 -3462 492266 -3226
rect 492502 -3462 502186 -3226
rect 502422 -3462 502506 -3226
rect 502742 -3462 512426 -3226
rect 512662 -3462 512746 -3226
rect 512982 -3462 522666 -3226
rect 522902 -3462 522986 -3226
rect 523222 -3462 532906 -3226
rect 533142 -3462 533226 -3226
rect 533462 -3462 543146 -3226
rect 543382 -3462 543466 -3226
rect 543702 -3462 553386 -3226
rect 553622 -3462 553706 -3226
rect 553942 -3462 563626 -3226
rect 563862 -3462 563946 -3226
rect 564182 -3462 573866 -3226
rect 574102 -3462 574186 -3226
rect 574422 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 10666 -3546
rect 10902 -3782 10986 -3546
rect 11222 -3782 20906 -3546
rect 21142 -3782 21226 -3546
rect 21462 -3782 31146 -3546
rect 31382 -3782 31466 -3546
rect 31702 -3782 41386 -3546
rect 41622 -3782 41706 -3546
rect 41942 -3782 51626 -3546
rect 51862 -3782 51946 -3546
rect 52182 -3782 61866 -3546
rect 62102 -3782 62186 -3546
rect 62422 -3782 72106 -3546
rect 72342 -3782 72426 -3546
rect 72662 -3782 82346 -3546
rect 82582 -3782 82666 -3546
rect 82902 -3782 92586 -3546
rect 92822 -3782 92906 -3546
rect 93142 -3782 102826 -3546
rect 103062 -3782 103146 -3546
rect 103382 -3782 113066 -3546
rect 113302 -3782 113386 -3546
rect 113622 -3782 123306 -3546
rect 123542 -3782 123626 -3546
rect 123862 -3782 133546 -3546
rect 133782 -3782 133866 -3546
rect 134102 -3782 143786 -3546
rect 144022 -3782 144106 -3546
rect 144342 -3782 154026 -3546
rect 154262 -3782 154346 -3546
rect 154582 -3782 164266 -3546
rect 164502 -3782 164586 -3546
rect 164822 -3782 174506 -3546
rect 174742 -3782 174826 -3546
rect 175062 -3782 184746 -3546
rect 184982 -3782 185066 -3546
rect 185302 -3782 194986 -3546
rect 195222 -3782 195306 -3546
rect 195542 -3782 205226 -3546
rect 205462 -3782 205546 -3546
rect 205782 -3782 215466 -3546
rect 215702 -3782 215786 -3546
rect 216022 -3782 225706 -3546
rect 225942 -3782 226026 -3546
rect 226262 -3782 235946 -3546
rect 236182 -3782 236266 -3546
rect 236502 -3782 246186 -3546
rect 246422 -3782 246506 -3546
rect 246742 -3782 256426 -3546
rect 256662 -3782 256746 -3546
rect 256982 -3782 266666 -3546
rect 266902 -3782 266986 -3546
rect 267222 -3782 276906 -3546
rect 277142 -3782 277226 -3546
rect 277462 -3782 287146 -3546
rect 287382 -3782 287466 -3546
rect 287702 -3782 297386 -3546
rect 297622 -3782 297706 -3546
rect 297942 -3782 307626 -3546
rect 307862 -3782 307946 -3546
rect 308182 -3782 317866 -3546
rect 318102 -3782 318186 -3546
rect 318422 -3782 328106 -3546
rect 328342 -3782 328426 -3546
rect 328662 -3782 338346 -3546
rect 338582 -3782 338666 -3546
rect 338902 -3782 348586 -3546
rect 348822 -3782 348906 -3546
rect 349142 -3782 358826 -3546
rect 359062 -3782 359146 -3546
rect 359382 -3782 369066 -3546
rect 369302 -3782 369386 -3546
rect 369622 -3782 379306 -3546
rect 379542 -3782 379626 -3546
rect 379862 -3782 389546 -3546
rect 389782 -3782 389866 -3546
rect 390102 -3782 399786 -3546
rect 400022 -3782 400106 -3546
rect 400342 -3782 410026 -3546
rect 410262 -3782 410346 -3546
rect 410582 -3782 420266 -3546
rect 420502 -3782 420586 -3546
rect 420822 -3782 430506 -3546
rect 430742 -3782 430826 -3546
rect 431062 -3782 440746 -3546
rect 440982 -3782 441066 -3546
rect 441302 -3782 450986 -3546
rect 451222 -3782 451306 -3546
rect 451542 -3782 461226 -3546
rect 461462 -3782 461546 -3546
rect 461782 -3782 471466 -3546
rect 471702 -3782 471786 -3546
rect 472022 -3782 481706 -3546
rect 481942 -3782 482026 -3546
rect 482262 -3782 491946 -3546
rect 492182 -3782 492266 -3546
rect 492502 -3782 502186 -3546
rect 502422 -3782 502506 -3546
rect 502742 -3782 512426 -3546
rect 512662 -3782 512746 -3546
rect 512982 -3782 522666 -3546
rect 522902 -3782 522986 -3546
rect 523222 -3782 532906 -3546
rect 533142 -3782 533226 -3546
rect 533462 -3782 543146 -3546
rect 543382 -3782 543466 -3546
rect 543702 -3782 553386 -3546
rect 553622 -3782 553706 -3546
rect 553942 -3782 563626 -3546
rect 563862 -3782 563946 -3546
rect 564182 -3782 573866 -3546
rect 574102 -3782 574186 -3546
rect 574422 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 19506 -4186
rect 19742 -4422 19826 -4186
rect 20062 -4422 29746 -4186
rect 29982 -4422 30066 -4186
rect 30302 -4422 39986 -4186
rect 40222 -4422 40306 -4186
rect 40542 -4422 50226 -4186
rect 50462 -4422 50546 -4186
rect 50782 -4422 60466 -4186
rect 60702 -4422 60786 -4186
rect 61022 -4422 70706 -4186
rect 70942 -4422 71026 -4186
rect 71262 -4422 80946 -4186
rect 81182 -4422 81266 -4186
rect 81502 -4422 91186 -4186
rect 91422 -4422 91506 -4186
rect 91742 -4422 101426 -4186
rect 101662 -4422 101746 -4186
rect 101982 -4422 111666 -4186
rect 111902 -4422 111986 -4186
rect 112222 -4422 121906 -4186
rect 122142 -4422 122226 -4186
rect 122462 -4422 132146 -4186
rect 132382 -4422 132466 -4186
rect 132702 -4422 142386 -4186
rect 142622 -4422 142706 -4186
rect 142942 -4422 152626 -4186
rect 152862 -4422 152946 -4186
rect 153182 -4422 162866 -4186
rect 163102 -4422 163186 -4186
rect 163422 -4422 173106 -4186
rect 173342 -4422 173426 -4186
rect 173662 -4422 183346 -4186
rect 183582 -4422 183666 -4186
rect 183902 -4422 193586 -4186
rect 193822 -4422 193906 -4186
rect 194142 -4422 203826 -4186
rect 204062 -4422 204146 -4186
rect 204382 -4422 214066 -4186
rect 214302 -4422 214386 -4186
rect 214622 -4422 224306 -4186
rect 224542 -4422 224626 -4186
rect 224862 -4422 234546 -4186
rect 234782 -4422 234866 -4186
rect 235102 -4422 244786 -4186
rect 245022 -4422 245106 -4186
rect 245342 -4422 255026 -4186
rect 255262 -4422 255346 -4186
rect 255582 -4422 265266 -4186
rect 265502 -4422 265586 -4186
rect 265822 -4422 275506 -4186
rect 275742 -4422 275826 -4186
rect 276062 -4422 285746 -4186
rect 285982 -4422 286066 -4186
rect 286302 -4422 295986 -4186
rect 296222 -4422 296306 -4186
rect 296542 -4422 306226 -4186
rect 306462 -4422 306546 -4186
rect 306782 -4422 316466 -4186
rect 316702 -4422 316786 -4186
rect 317022 -4422 326706 -4186
rect 326942 -4422 327026 -4186
rect 327262 -4422 336946 -4186
rect 337182 -4422 337266 -4186
rect 337502 -4422 347186 -4186
rect 347422 -4422 347506 -4186
rect 347742 -4422 357426 -4186
rect 357662 -4422 357746 -4186
rect 357982 -4422 367666 -4186
rect 367902 -4422 367986 -4186
rect 368222 -4422 377906 -4186
rect 378142 -4422 378226 -4186
rect 378462 -4422 388146 -4186
rect 388382 -4422 388466 -4186
rect 388702 -4422 398386 -4186
rect 398622 -4422 398706 -4186
rect 398942 -4422 408626 -4186
rect 408862 -4422 408946 -4186
rect 409182 -4422 418866 -4186
rect 419102 -4422 419186 -4186
rect 419422 -4422 429106 -4186
rect 429342 -4422 429426 -4186
rect 429662 -4422 439346 -4186
rect 439582 -4422 439666 -4186
rect 439902 -4422 449586 -4186
rect 449822 -4422 449906 -4186
rect 450142 -4422 459826 -4186
rect 460062 -4422 460146 -4186
rect 460382 -4422 470066 -4186
rect 470302 -4422 470386 -4186
rect 470622 -4422 480306 -4186
rect 480542 -4422 480626 -4186
rect 480862 -4422 490546 -4186
rect 490782 -4422 490866 -4186
rect 491102 -4422 500786 -4186
rect 501022 -4422 501106 -4186
rect 501342 -4422 511026 -4186
rect 511262 -4422 511346 -4186
rect 511582 -4422 521266 -4186
rect 521502 -4422 521586 -4186
rect 521822 -4422 531506 -4186
rect 531742 -4422 531826 -4186
rect 532062 -4422 541746 -4186
rect 541982 -4422 542066 -4186
rect 542302 -4422 551986 -4186
rect 552222 -4422 552306 -4186
rect 552542 -4422 562226 -4186
rect 562462 -4422 562546 -4186
rect 562782 -4422 572466 -4186
rect 572702 -4422 572786 -4186
rect 573022 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 19506 -4506
rect 19742 -4742 19826 -4506
rect 20062 -4742 29746 -4506
rect 29982 -4742 30066 -4506
rect 30302 -4742 39986 -4506
rect 40222 -4742 40306 -4506
rect 40542 -4742 50226 -4506
rect 50462 -4742 50546 -4506
rect 50782 -4742 60466 -4506
rect 60702 -4742 60786 -4506
rect 61022 -4742 70706 -4506
rect 70942 -4742 71026 -4506
rect 71262 -4742 80946 -4506
rect 81182 -4742 81266 -4506
rect 81502 -4742 91186 -4506
rect 91422 -4742 91506 -4506
rect 91742 -4742 101426 -4506
rect 101662 -4742 101746 -4506
rect 101982 -4742 111666 -4506
rect 111902 -4742 111986 -4506
rect 112222 -4742 121906 -4506
rect 122142 -4742 122226 -4506
rect 122462 -4742 132146 -4506
rect 132382 -4742 132466 -4506
rect 132702 -4742 142386 -4506
rect 142622 -4742 142706 -4506
rect 142942 -4742 152626 -4506
rect 152862 -4742 152946 -4506
rect 153182 -4742 162866 -4506
rect 163102 -4742 163186 -4506
rect 163422 -4742 173106 -4506
rect 173342 -4742 173426 -4506
rect 173662 -4742 183346 -4506
rect 183582 -4742 183666 -4506
rect 183902 -4742 193586 -4506
rect 193822 -4742 193906 -4506
rect 194142 -4742 203826 -4506
rect 204062 -4742 204146 -4506
rect 204382 -4742 214066 -4506
rect 214302 -4742 214386 -4506
rect 214622 -4742 224306 -4506
rect 224542 -4742 224626 -4506
rect 224862 -4742 234546 -4506
rect 234782 -4742 234866 -4506
rect 235102 -4742 244786 -4506
rect 245022 -4742 245106 -4506
rect 245342 -4742 255026 -4506
rect 255262 -4742 255346 -4506
rect 255582 -4742 265266 -4506
rect 265502 -4742 265586 -4506
rect 265822 -4742 275506 -4506
rect 275742 -4742 275826 -4506
rect 276062 -4742 285746 -4506
rect 285982 -4742 286066 -4506
rect 286302 -4742 295986 -4506
rect 296222 -4742 296306 -4506
rect 296542 -4742 306226 -4506
rect 306462 -4742 306546 -4506
rect 306782 -4742 316466 -4506
rect 316702 -4742 316786 -4506
rect 317022 -4742 326706 -4506
rect 326942 -4742 327026 -4506
rect 327262 -4742 336946 -4506
rect 337182 -4742 337266 -4506
rect 337502 -4742 347186 -4506
rect 347422 -4742 347506 -4506
rect 347742 -4742 357426 -4506
rect 357662 -4742 357746 -4506
rect 357982 -4742 367666 -4506
rect 367902 -4742 367986 -4506
rect 368222 -4742 377906 -4506
rect 378142 -4742 378226 -4506
rect 378462 -4742 388146 -4506
rect 388382 -4742 388466 -4506
rect 388702 -4742 398386 -4506
rect 398622 -4742 398706 -4506
rect 398942 -4742 408626 -4506
rect 408862 -4742 408946 -4506
rect 409182 -4742 418866 -4506
rect 419102 -4742 419186 -4506
rect 419422 -4742 429106 -4506
rect 429342 -4742 429426 -4506
rect 429662 -4742 439346 -4506
rect 439582 -4742 439666 -4506
rect 439902 -4742 449586 -4506
rect 449822 -4742 449906 -4506
rect 450142 -4742 459826 -4506
rect 460062 -4742 460146 -4506
rect 460382 -4742 470066 -4506
rect 470302 -4742 470386 -4506
rect 470622 -4742 480306 -4506
rect 480542 -4742 480626 -4506
rect 480862 -4742 490546 -4506
rect 490782 -4742 490866 -4506
rect 491102 -4742 500786 -4506
rect 501022 -4742 501106 -4506
rect 501342 -4742 511026 -4506
rect 511262 -4742 511346 -4506
rect 511582 -4742 521266 -4506
rect 521502 -4742 521586 -4506
rect 521822 -4742 531506 -4506
rect 531742 -4742 531826 -4506
rect 532062 -4742 541746 -4506
rect 541982 -4742 542066 -4506
rect 542302 -4742 551986 -4506
rect 552222 -4742 552306 -4506
rect 552542 -4742 562226 -4506
rect 562462 -4742 562546 -4506
rect 562782 -4742 572466 -4506
rect 572702 -4742 572786 -4506
rect 573022 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 14386 -5146
rect 14622 -5382 14706 -5146
rect 14942 -5382 24626 -5146
rect 24862 -5382 24946 -5146
rect 25182 -5382 34866 -5146
rect 35102 -5382 35186 -5146
rect 35422 -5382 45106 -5146
rect 45342 -5382 45426 -5146
rect 45662 -5382 55346 -5146
rect 55582 -5382 55666 -5146
rect 55902 -5382 65586 -5146
rect 65822 -5382 65906 -5146
rect 66142 -5382 75826 -5146
rect 76062 -5382 76146 -5146
rect 76382 -5382 86066 -5146
rect 86302 -5382 86386 -5146
rect 86622 -5382 96306 -5146
rect 96542 -5382 96626 -5146
rect 96862 -5382 106546 -5146
rect 106782 -5382 106866 -5146
rect 107102 -5382 116786 -5146
rect 117022 -5382 117106 -5146
rect 117342 -5382 127026 -5146
rect 127262 -5382 127346 -5146
rect 127582 -5382 137266 -5146
rect 137502 -5382 137586 -5146
rect 137822 -5382 147506 -5146
rect 147742 -5382 147826 -5146
rect 148062 -5382 157746 -5146
rect 157982 -5382 158066 -5146
rect 158302 -5382 167986 -5146
rect 168222 -5382 168306 -5146
rect 168542 -5382 178226 -5146
rect 178462 -5382 178546 -5146
rect 178782 -5382 188466 -5146
rect 188702 -5382 188786 -5146
rect 189022 -5382 198706 -5146
rect 198942 -5382 199026 -5146
rect 199262 -5382 208946 -5146
rect 209182 -5382 209266 -5146
rect 209502 -5382 219186 -5146
rect 219422 -5382 219506 -5146
rect 219742 -5382 229426 -5146
rect 229662 -5382 229746 -5146
rect 229982 -5382 239666 -5146
rect 239902 -5382 239986 -5146
rect 240222 -5382 249906 -5146
rect 250142 -5382 250226 -5146
rect 250462 -5382 260146 -5146
rect 260382 -5382 260466 -5146
rect 260702 -5382 270386 -5146
rect 270622 -5382 270706 -5146
rect 270942 -5382 280626 -5146
rect 280862 -5382 280946 -5146
rect 281182 -5382 290866 -5146
rect 291102 -5382 291186 -5146
rect 291422 -5382 301106 -5146
rect 301342 -5382 301426 -5146
rect 301662 -5382 311346 -5146
rect 311582 -5382 311666 -5146
rect 311902 -5382 321586 -5146
rect 321822 -5382 321906 -5146
rect 322142 -5382 331826 -5146
rect 332062 -5382 332146 -5146
rect 332382 -5382 342066 -5146
rect 342302 -5382 342386 -5146
rect 342622 -5382 352306 -5146
rect 352542 -5382 352626 -5146
rect 352862 -5382 362546 -5146
rect 362782 -5382 362866 -5146
rect 363102 -5382 372786 -5146
rect 373022 -5382 373106 -5146
rect 373342 -5382 383026 -5146
rect 383262 -5382 383346 -5146
rect 383582 -5382 393266 -5146
rect 393502 -5382 393586 -5146
rect 393822 -5382 403506 -5146
rect 403742 -5382 403826 -5146
rect 404062 -5382 413746 -5146
rect 413982 -5382 414066 -5146
rect 414302 -5382 423986 -5146
rect 424222 -5382 424306 -5146
rect 424542 -5382 434226 -5146
rect 434462 -5382 434546 -5146
rect 434782 -5382 444466 -5146
rect 444702 -5382 444786 -5146
rect 445022 -5382 454706 -5146
rect 454942 -5382 455026 -5146
rect 455262 -5382 464946 -5146
rect 465182 -5382 465266 -5146
rect 465502 -5382 475186 -5146
rect 475422 -5382 475506 -5146
rect 475742 -5382 485426 -5146
rect 485662 -5382 485746 -5146
rect 485982 -5382 495666 -5146
rect 495902 -5382 495986 -5146
rect 496222 -5382 505906 -5146
rect 506142 -5382 506226 -5146
rect 506462 -5382 516146 -5146
rect 516382 -5382 516466 -5146
rect 516702 -5382 526386 -5146
rect 526622 -5382 526706 -5146
rect 526942 -5382 536626 -5146
rect 536862 -5382 536946 -5146
rect 537182 -5382 546866 -5146
rect 547102 -5382 547186 -5146
rect 547422 -5382 557106 -5146
rect 557342 -5382 557426 -5146
rect 557662 -5382 567346 -5146
rect 567582 -5382 567666 -5146
rect 567902 -5382 577586 -5146
rect 577822 -5382 577906 -5146
rect 578142 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 14386 -5466
rect 14622 -5702 14706 -5466
rect 14942 -5702 24626 -5466
rect 24862 -5702 24946 -5466
rect 25182 -5702 34866 -5466
rect 35102 -5702 35186 -5466
rect 35422 -5702 45106 -5466
rect 45342 -5702 45426 -5466
rect 45662 -5702 55346 -5466
rect 55582 -5702 55666 -5466
rect 55902 -5702 65586 -5466
rect 65822 -5702 65906 -5466
rect 66142 -5702 75826 -5466
rect 76062 -5702 76146 -5466
rect 76382 -5702 86066 -5466
rect 86302 -5702 86386 -5466
rect 86622 -5702 96306 -5466
rect 96542 -5702 96626 -5466
rect 96862 -5702 106546 -5466
rect 106782 -5702 106866 -5466
rect 107102 -5702 116786 -5466
rect 117022 -5702 117106 -5466
rect 117342 -5702 127026 -5466
rect 127262 -5702 127346 -5466
rect 127582 -5702 137266 -5466
rect 137502 -5702 137586 -5466
rect 137822 -5702 147506 -5466
rect 147742 -5702 147826 -5466
rect 148062 -5702 157746 -5466
rect 157982 -5702 158066 -5466
rect 158302 -5702 167986 -5466
rect 168222 -5702 168306 -5466
rect 168542 -5702 178226 -5466
rect 178462 -5702 178546 -5466
rect 178782 -5702 188466 -5466
rect 188702 -5702 188786 -5466
rect 189022 -5702 198706 -5466
rect 198942 -5702 199026 -5466
rect 199262 -5702 208946 -5466
rect 209182 -5702 209266 -5466
rect 209502 -5702 219186 -5466
rect 219422 -5702 219506 -5466
rect 219742 -5702 229426 -5466
rect 229662 -5702 229746 -5466
rect 229982 -5702 239666 -5466
rect 239902 -5702 239986 -5466
rect 240222 -5702 249906 -5466
rect 250142 -5702 250226 -5466
rect 250462 -5702 260146 -5466
rect 260382 -5702 260466 -5466
rect 260702 -5702 270386 -5466
rect 270622 -5702 270706 -5466
rect 270942 -5702 280626 -5466
rect 280862 -5702 280946 -5466
rect 281182 -5702 290866 -5466
rect 291102 -5702 291186 -5466
rect 291422 -5702 301106 -5466
rect 301342 -5702 301426 -5466
rect 301662 -5702 311346 -5466
rect 311582 -5702 311666 -5466
rect 311902 -5702 321586 -5466
rect 321822 -5702 321906 -5466
rect 322142 -5702 331826 -5466
rect 332062 -5702 332146 -5466
rect 332382 -5702 342066 -5466
rect 342302 -5702 342386 -5466
rect 342622 -5702 352306 -5466
rect 352542 -5702 352626 -5466
rect 352862 -5702 362546 -5466
rect 362782 -5702 362866 -5466
rect 363102 -5702 372786 -5466
rect 373022 -5702 373106 -5466
rect 373342 -5702 383026 -5466
rect 383262 -5702 383346 -5466
rect 383582 -5702 393266 -5466
rect 393502 -5702 393586 -5466
rect 393822 -5702 403506 -5466
rect 403742 -5702 403826 -5466
rect 404062 -5702 413746 -5466
rect 413982 -5702 414066 -5466
rect 414302 -5702 423986 -5466
rect 424222 -5702 424306 -5466
rect 424542 -5702 434226 -5466
rect 434462 -5702 434546 -5466
rect 434782 -5702 444466 -5466
rect 444702 -5702 444786 -5466
rect 445022 -5702 454706 -5466
rect 454942 -5702 455026 -5466
rect 455262 -5702 464946 -5466
rect 465182 -5702 465266 -5466
rect 465502 -5702 475186 -5466
rect 475422 -5702 475506 -5466
rect 475742 -5702 485426 -5466
rect 485662 -5702 485746 -5466
rect 485982 -5702 495666 -5466
rect 495902 -5702 495986 -5466
rect 496222 -5702 505906 -5466
rect 506142 -5702 506226 -5466
rect 506462 -5702 516146 -5466
rect 516382 -5702 516466 -5466
rect 516702 -5702 526386 -5466
rect 526622 -5702 526706 -5466
rect 526942 -5702 536626 -5466
rect 536862 -5702 536946 -5466
rect 537182 -5702 546866 -5466
rect 547102 -5702 547186 -5466
rect 547422 -5702 557106 -5466
rect 557342 -5702 557426 -5466
rect 557662 -5702 567346 -5466
rect 567582 -5702 567666 -5466
rect 567902 -5702 577586 -5466
rect 577822 -5702 577906 -5466
rect 578142 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 23226 -6106
rect 23462 -6342 23546 -6106
rect 23782 -6342 33466 -6106
rect 33702 -6342 33786 -6106
rect 34022 -6342 43706 -6106
rect 43942 -6342 44026 -6106
rect 44262 -6342 53946 -6106
rect 54182 -6342 54266 -6106
rect 54502 -6342 64186 -6106
rect 64422 -6342 64506 -6106
rect 64742 -6342 74426 -6106
rect 74662 -6342 74746 -6106
rect 74982 -6342 84666 -6106
rect 84902 -6342 84986 -6106
rect 85222 -6342 94906 -6106
rect 95142 -6342 95226 -6106
rect 95462 -6342 105146 -6106
rect 105382 -6342 105466 -6106
rect 105702 -6342 115386 -6106
rect 115622 -6342 115706 -6106
rect 115942 -6342 125626 -6106
rect 125862 -6342 125946 -6106
rect 126182 -6342 135866 -6106
rect 136102 -6342 136186 -6106
rect 136422 -6342 146106 -6106
rect 146342 -6342 146426 -6106
rect 146662 -6342 156346 -6106
rect 156582 -6342 156666 -6106
rect 156902 -6342 166586 -6106
rect 166822 -6342 166906 -6106
rect 167142 -6342 176826 -6106
rect 177062 -6342 177146 -6106
rect 177382 -6342 187066 -6106
rect 187302 -6342 187386 -6106
rect 187622 -6342 197306 -6106
rect 197542 -6342 197626 -6106
rect 197862 -6342 207546 -6106
rect 207782 -6342 207866 -6106
rect 208102 -6342 217786 -6106
rect 218022 -6342 218106 -6106
rect 218342 -6342 228026 -6106
rect 228262 -6342 228346 -6106
rect 228582 -6342 238266 -6106
rect 238502 -6342 238586 -6106
rect 238822 -6342 248506 -6106
rect 248742 -6342 248826 -6106
rect 249062 -6342 258746 -6106
rect 258982 -6342 259066 -6106
rect 259302 -6342 268986 -6106
rect 269222 -6342 269306 -6106
rect 269542 -6342 279226 -6106
rect 279462 -6342 279546 -6106
rect 279782 -6342 289466 -6106
rect 289702 -6342 289786 -6106
rect 290022 -6342 299706 -6106
rect 299942 -6342 300026 -6106
rect 300262 -6342 309946 -6106
rect 310182 -6342 310266 -6106
rect 310502 -6342 320186 -6106
rect 320422 -6342 320506 -6106
rect 320742 -6342 330426 -6106
rect 330662 -6342 330746 -6106
rect 330982 -6342 340666 -6106
rect 340902 -6342 340986 -6106
rect 341222 -6342 350906 -6106
rect 351142 -6342 351226 -6106
rect 351462 -6342 361146 -6106
rect 361382 -6342 361466 -6106
rect 361702 -6342 371386 -6106
rect 371622 -6342 371706 -6106
rect 371942 -6342 381626 -6106
rect 381862 -6342 381946 -6106
rect 382182 -6342 391866 -6106
rect 392102 -6342 392186 -6106
rect 392422 -6342 402106 -6106
rect 402342 -6342 402426 -6106
rect 402662 -6342 412346 -6106
rect 412582 -6342 412666 -6106
rect 412902 -6342 422586 -6106
rect 422822 -6342 422906 -6106
rect 423142 -6342 432826 -6106
rect 433062 -6342 433146 -6106
rect 433382 -6342 443066 -6106
rect 443302 -6342 443386 -6106
rect 443622 -6342 453306 -6106
rect 453542 -6342 453626 -6106
rect 453862 -6342 463546 -6106
rect 463782 -6342 463866 -6106
rect 464102 -6342 473786 -6106
rect 474022 -6342 474106 -6106
rect 474342 -6342 484026 -6106
rect 484262 -6342 484346 -6106
rect 484582 -6342 494266 -6106
rect 494502 -6342 494586 -6106
rect 494822 -6342 504506 -6106
rect 504742 -6342 504826 -6106
rect 505062 -6342 514746 -6106
rect 514982 -6342 515066 -6106
rect 515302 -6342 524986 -6106
rect 525222 -6342 525306 -6106
rect 525542 -6342 535226 -6106
rect 535462 -6342 535546 -6106
rect 535782 -6342 545466 -6106
rect 545702 -6342 545786 -6106
rect 546022 -6342 555706 -6106
rect 555942 -6342 556026 -6106
rect 556262 -6342 565946 -6106
rect 566182 -6342 566266 -6106
rect 566502 -6342 576186 -6106
rect 576422 -6342 576506 -6106
rect 576742 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 23226 -6426
rect 23462 -6662 23546 -6426
rect 23782 -6662 33466 -6426
rect 33702 -6662 33786 -6426
rect 34022 -6662 43706 -6426
rect 43942 -6662 44026 -6426
rect 44262 -6662 53946 -6426
rect 54182 -6662 54266 -6426
rect 54502 -6662 64186 -6426
rect 64422 -6662 64506 -6426
rect 64742 -6662 74426 -6426
rect 74662 -6662 74746 -6426
rect 74982 -6662 84666 -6426
rect 84902 -6662 84986 -6426
rect 85222 -6662 94906 -6426
rect 95142 -6662 95226 -6426
rect 95462 -6662 105146 -6426
rect 105382 -6662 105466 -6426
rect 105702 -6662 115386 -6426
rect 115622 -6662 115706 -6426
rect 115942 -6662 125626 -6426
rect 125862 -6662 125946 -6426
rect 126182 -6662 135866 -6426
rect 136102 -6662 136186 -6426
rect 136422 -6662 146106 -6426
rect 146342 -6662 146426 -6426
rect 146662 -6662 156346 -6426
rect 156582 -6662 156666 -6426
rect 156902 -6662 166586 -6426
rect 166822 -6662 166906 -6426
rect 167142 -6662 176826 -6426
rect 177062 -6662 177146 -6426
rect 177382 -6662 187066 -6426
rect 187302 -6662 187386 -6426
rect 187622 -6662 197306 -6426
rect 197542 -6662 197626 -6426
rect 197862 -6662 207546 -6426
rect 207782 -6662 207866 -6426
rect 208102 -6662 217786 -6426
rect 218022 -6662 218106 -6426
rect 218342 -6662 228026 -6426
rect 228262 -6662 228346 -6426
rect 228582 -6662 238266 -6426
rect 238502 -6662 238586 -6426
rect 238822 -6662 248506 -6426
rect 248742 -6662 248826 -6426
rect 249062 -6662 258746 -6426
rect 258982 -6662 259066 -6426
rect 259302 -6662 268986 -6426
rect 269222 -6662 269306 -6426
rect 269542 -6662 279226 -6426
rect 279462 -6662 279546 -6426
rect 279782 -6662 289466 -6426
rect 289702 -6662 289786 -6426
rect 290022 -6662 299706 -6426
rect 299942 -6662 300026 -6426
rect 300262 -6662 309946 -6426
rect 310182 -6662 310266 -6426
rect 310502 -6662 320186 -6426
rect 320422 -6662 320506 -6426
rect 320742 -6662 330426 -6426
rect 330662 -6662 330746 -6426
rect 330982 -6662 340666 -6426
rect 340902 -6662 340986 -6426
rect 341222 -6662 350906 -6426
rect 351142 -6662 351226 -6426
rect 351462 -6662 361146 -6426
rect 361382 -6662 361466 -6426
rect 361702 -6662 371386 -6426
rect 371622 -6662 371706 -6426
rect 371942 -6662 381626 -6426
rect 381862 -6662 381946 -6426
rect 382182 -6662 391866 -6426
rect 392102 -6662 392186 -6426
rect 392422 -6662 402106 -6426
rect 402342 -6662 402426 -6426
rect 402662 -6662 412346 -6426
rect 412582 -6662 412666 -6426
rect 412902 -6662 422586 -6426
rect 422822 -6662 422906 -6426
rect 423142 -6662 432826 -6426
rect 433062 -6662 433146 -6426
rect 433382 -6662 443066 -6426
rect 443302 -6662 443386 -6426
rect 443622 -6662 453306 -6426
rect 453542 -6662 453626 -6426
rect 453862 -6662 463546 -6426
rect 463782 -6662 463866 -6426
rect 464102 -6662 473786 -6426
rect 474022 -6662 474106 -6426
rect 474342 -6662 484026 -6426
rect 484262 -6662 484346 -6426
rect 484582 -6662 494266 -6426
rect 494502 -6662 494586 -6426
rect 494822 -6662 504506 -6426
rect 504742 -6662 504826 -6426
rect 505062 -6662 514746 -6426
rect 514982 -6662 515066 -6426
rect 515302 -6662 524986 -6426
rect 525222 -6662 525306 -6426
rect 525542 -6662 535226 -6426
rect 535462 -6662 535546 -6426
rect 535782 -6662 545466 -6426
rect 545702 -6662 545786 -6426
rect 546022 -6662 555706 -6426
rect 555942 -6662 556026 -6426
rect 556262 -6662 565946 -6426
rect 566182 -6662 566266 -6426
rect 566502 -6662 576186 -6426
rect 576422 -6662 576506 -6426
rect 576742 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 18106 -7066
rect 18342 -7302 18426 -7066
rect 18662 -7302 28346 -7066
rect 28582 -7302 28666 -7066
rect 28902 -7302 38586 -7066
rect 38822 -7302 38906 -7066
rect 39142 -7302 48826 -7066
rect 49062 -7302 49146 -7066
rect 49382 -7302 59066 -7066
rect 59302 -7302 59386 -7066
rect 59622 -7302 69306 -7066
rect 69542 -7302 69626 -7066
rect 69862 -7302 79546 -7066
rect 79782 -7302 79866 -7066
rect 80102 -7302 89786 -7066
rect 90022 -7302 90106 -7066
rect 90342 -7302 100026 -7066
rect 100262 -7302 100346 -7066
rect 100582 -7302 110266 -7066
rect 110502 -7302 110586 -7066
rect 110822 -7302 120506 -7066
rect 120742 -7302 120826 -7066
rect 121062 -7302 130746 -7066
rect 130982 -7302 131066 -7066
rect 131302 -7302 140986 -7066
rect 141222 -7302 141306 -7066
rect 141542 -7302 151226 -7066
rect 151462 -7302 151546 -7066
rect 151782 -7302 161466 -7066
rect 161702 -7302 161786 -7066
rect 162022 -7302 171706 -7066
rect 171942 -7302 172026 -7066
rect 172262 -7302 181946 -7066
rect 182182 -7302 182266 -7066
rect 182502 -7302 192186 -7066
rect 192422 -7302 192506 -7066
rect 192742 -7302 202426 -7066
rect 202662 -7302 202746 -7066
rect 202982 -7302 212666 -7066
rect 212902 -7302 212986 -7066
rect 213222 -7302 222906 -7066
rect 223142 -7302 223226 -7066
rect 223462 -7302 233146 -7066
rect 233382 -7302 233466 -7066
rect 233702 -7302 243386 -7066
rect 243622 -7302 243706 -7066
rect 243942 -7302 253626 -7066
rect 253862 -7302 253946 -7066
rect 254182 -7302 263866 -7066
rect 264102 -7302 264186 -7066
rect 264422 -7302 274106 -7066
rect 274342 -7302 274426 -7066
rect 274662 -7302 284346 -7066
rect 284582 -7302 284666 -7066
rect 284902 -7302 294586 -7066
rect 294822 -7302 294906 -7066
rect 295142 -7302 304826 -7066
rect 305062 -7302 305146 -7066
rect 305382 -7302 315066 -7066
rect 315302 -7302 315386 -7066
rect 315622 -7302 325306 -7066
rect 325542 -7302 325626 -7066
rect 325862 -7302 335546 -7066
rect 335782 -7302 335866 -7066
rect 336102 -7302 345786 -7066
rect 346022 -7302 346106 -7066
rect 346342 -7302 356026 -7066
rect 356262 -7302 356346 -7066
rect 356582 -7302 366266 -7066
rect 366502 -7302 366586 -7066
rect 366822 -7302 376506 -7066
rect 376742 -7302 376826 -7066
rect 377062 -7302 386746 -7066
rect 386982 -7302 387066 -7066
rect 387302 -7302 396986 -7066
rect 397222 -7302 397306 -7066
rect 397542 -7302 407226 -7066
rect 407462 -7302 407546 -7066
rect 407782 -7302 417466 -7066
rect 417702 -7302 417786 -7066
rect 418022 -7302 427706 -7066
rect 427942 -7302 428026 -7066
rect 428262 -7302 437946 -7066
rect 438182 -7302 438266 -7066
rect 438502 -7302 448186 -7066
rect 448422 -7302 448506 -7066
rect 448742 -7302 458426 -7066
rect 458662 -7302 458746 -7066
rect 458982 -7302 468666 -7066
rect 468902 -7302 468986 -7066
rect 469222 -7302 478906 -7066
rect 479142 -7302 479226 -7066
rect 479462 -7302 489146 -7066
rect 489382 -7302 489466 -7066
rect 489702 -7302 499386 -7066
rect 499622 -7302 499706 -7066
rect 499942 -7302 509626 -7066
rect 509862 -7302 509946 -7066
rect 510182 -7302 519866 -7066
rect 520102 -7302 520186 -7066
rect 520422 -7302 530106 -7066
rect 530342 -7302 530426 -7066
rect 530662 -7302 540346 -7066
rect 540582 -7302 540666 -7066
rect 540902 -7302 550586 -7066
rect 550822 -7302 550906 -7066
rect 551142 -7302 560826 -7066
rect 561062 -7302 561146 -7066
rect 561382 -7302 571066 -7066
rect 571302 -7302 571386 -7066
rect 571622 -7302 581306 -7066
rect 581542 -7302 581626 -7066
rect 581862 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 18106 -7386
rect 18342 -7622 18426 -7386
rect 18662 -7622 28346 -7386
rect 28582 -7622 28666 -7386
rect 28902 -7622 38586 -7386
rect 38822 -7622 38906 -7386
rect 39142 -7622 48826 -7386
rect 49062 -7622 49146 -7386
rect 49382 -7622 59066 -7386
rect 59302 -7622 59386 -7386
rect 59622 -7622 69306 -7386
rect 69542 -7622 69626 -7386
rect 69862 -7622 79546 -7386
rect 79782 -7622 79866 -7386
rect 80102 -7622 89786 -7386
rect 90022 -7622 90106 -7386
rect 90342 -7622 100026 -7386
rect 100262 -7622 100346 -7386
rect 100582 -7622 110266 -7386
rect 110502 -7622 110586 -7386
rect 110822 -7622 120506 -7386
rect 120742 -7622 120826 -7386
rect 121062 -7622 130746 -7386
rect 130982 -7622 131066 -7386
rect 131302 -7622 140986 -7386
rect 141222 -7622 141306 -7386
rect 141542 -7622 151226 -7386
rect 151462 -7622 151546 -7386
rect 151782 -7622 161466 -7386
rect 161702 -7622 161786 -7386
rect 162022 -7622 171706 -7386
rect 171942 -7622 172026 -7386
rect 172262 -7622 181946 -7386
rect 182182 -7622 182266 -7386
rect 182502 -7622 192186 -7386
rect 192422 -7622 192506 -7386
rect 192742 -7622 202426 -7386
rect 202662 -7622 202746 -7386
rect 202982 -7622 212666 -7386
rect 212902 -7622 212986 -7386
rect 213222 -7622 222906 -7386
rect 223142 -7622 223226 -7386
rect 223462 -7622 233146 -7386
rect 233382 -7622 233466 -7386
rect 233702 -7622 243386 -7386
rect 243622 -7622 243706 -7386
rect 243942 -7622 253626 -7386
rect 253862 -7622 253946 -7386
rect 254182 -7622 263866 -7386
rect 264102 -7622 264186 -7386
rect 264422 -7622 274106 -7386
rect 274342 -7622 274426 -7386
rect 274662 -7622 284346 -7386
rect 284582 -7622 284666 -7386
rect 284902 -7622 294586 -7386
rect 294822 -7622 294906 -7386
rect 295142 -7622 304826 -7386
rect 305062 -7622 305146 -7386
rect 305382 -7622 315066 -7386
rect 315302 -7622 315386 -7386
rect 315622 -7622 325306 -7386
rect 325542 -7622 325626 -7386
rect 325862 -7622 335546 -7386
rect 335782 -7622 335866 -7386
rect 336102 -7622 345786 -7386
rect 346022 -7622 346106 -7386
rect 346342 -7622 356026 -7386
rect 356262 -7622 356346 -7386
rect 356582 -7622 366266 -7386
rect 366502 -7622 366586 -7386
rect 366822 -7622 376506 -7386
rect 376742 -7622 376826 -7386
rect 377062 -7622 386746 -7386
rect 386982 -7622 387066 -7386
rect 387302 -7622 396986 -7386
rect 397222 -7622 397306 -7386
rect 397542 -7622 407226 -7386
rect 407462 -7622 407546 -7386
rect 407782 -7622 417466 -7386
rect 417702 -7622 417786 -7386
rect 418022 -7622 427706 -7386
rect 427942 -7622 428026 -7386
rect 428262 -7622 437946 -7386
rect 438182 -7622 438266 -7386
rect 438502 -7622 448186 -7386
rect 448422 -7622 448506 -7386
rect 448742 -7622 458426 -7386
rect 458662 -7622 458746 -7386
rect 458982 -7622 468666 -7386
rect 468902 -7622 468986 -7386
rect 469222 -7622 478906 -7386
rect 479142 -7622 479226 -7386
rect 479462 -7622 489146 -7386
rect 489382 -7622 489466 -7386
rect 489702 -7622 499386 -7386
rect 499622 -7622 499706 -7386
rect 499942 -7622 509626 -7386
rect 509862 -7622 509946 -7386
rect 510182 -7622 519866 -7386
rect 520102 -7622 520186 -7386
rect 520422 -7622 530106 -7386
rect 530342 -7622 530426 -7386
rect 530662 -7622 540346 -7386
rect 540582 -7622 540666 -7386
rect 540902 -7622 550586 -7386
rect 550822 -7622 550906 -7386
rect 551142 -7622 560826 -7386
rect 561062 -7622 561146 -7386
rect 561382 -7622 571066 -7386
rect 571302 -7622 571386 -7386
rect 571622 -7622 581306 -7386
rect 581542 -7622 581626 -7386
rect 581862 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use top  dut
timestamp 0
transform 1 0 19080 0 1 15000
box 0 0 520000 640000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 22274 -1894 22894 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 32514 -1894 33134 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 42754 -1894 43374 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 52994 -1894 53614 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 63234 -1894 63854 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73474 -1894 74094 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 83714 -1894 84334 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 93954 -1894 94574 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 104194 -1894 104814 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 114434 -1894 115054 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 124674 -1894 125294 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 134914 -1894 135534 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145154 -1894 145774 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 155394 -1894 156014 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 165634 -1894 166254 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 175874 -1894 176494 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 186114 -1894 186734 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 196354 -1894 196974 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 206594 -1894 207214 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 216834 -1894 217454 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 227074 -1894 227694 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 237314 -1894 237934 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 247554 -1894 248174 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 257794 -1894 258414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 268034 -1894 268654 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 278274 -1894 278894 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 288514 -1894 289134 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 298754 -1894 299374 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 308994 -1894 309614 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 319234 -1894 319854 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 329474 -1894 330094 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 339714 -1894 340334 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 349954 -1894 350574 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 360194 -1894 360814 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 370434 -1894 371054 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 380674 -1894 381294 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 390914 -1894 391534 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 401154 -1894 401774 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 411394 -1894 412014 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 421634 -1894 422254 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 431874 -1894 432494 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 442114 -1894 442734 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 452354 -1894 452974 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 462594 -1894 463214 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 472834 -1894 473454 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 483074 -1894 483694 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 493314 -1894 493934 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 503554 -1894 504174 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 513794 -1894 514414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 524034 -1894 524654 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 534274 -1894 534894 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 12034 -1894 12654 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 22274 657000 22894 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 32514 657000 33134 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 42754 657000 43374 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 52994 657000 53614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 63234 657000 63854 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73474 657000 74094 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 83714 657000 84334 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 93954 657000 94574 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 104194 657000 104814 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 114434 657000 115054 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 124674 657000 125294 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 134914 657000 135534 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145154 657000 145774 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 155394 657000 156014 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 165634 657000 166254 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 175874 657000 176494 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 186114 657000 186734 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 196354 657000 196974 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 206594 657000 207214 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 216834 657000 217454 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 227074 657000 227694 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 237314 657000 237934 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 247554 657000 248174 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 257794 657000 258414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 268034 657000 268654 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 278274 657000 278894 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 288514 657000 289134 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 298754 657000 299374 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 308994 657000 309614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 319234 657000 319854 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 329474 657000 330094 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 339714 657000 340334 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 349954 657000 350574 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 360194 657000 360814 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 370434 657000 371054 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 380674 657000 381294 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 390914 657000 391534 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 401154 657000 401774 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 411394 657000 412014 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 421634 657000 422254 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 431874 657000 432494 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 442114 657000 442734 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 452354 657000 452974 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 462594 657000 463214 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 472834 657000 473454 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 483074 657000 483694 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 493314 657000 493934 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 503554 657000 504174 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 513794 657000 514414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 524034 657000 524654 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 534274 657000 534894 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 544514 -1894 545134 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 554754 -1894 555374 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 564994 -1894 565614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 575234 -1894 575854 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 25994 -3814 26614 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 36234 -3814 36854 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 46474 -3814 47094 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 56714 -3814 57334 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 66954 -3814 67574 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77194 -3814 77814 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 87434 -3814 88054 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 97674 -3814 98294 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 107914 -3814 108534 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 118154 -3814 118774 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 128394 -3814 129014 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 138634 -3814 139254 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 148874 -3814 149494 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 159114 -3814 159734 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 169354 -3814 169974 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 179594 -3814 180214 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 189834 -3814 190454 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 200074 -3814 200694 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 210314 -3814 210934 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 220554 -3814 221174 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 230794 -3814 231414 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 241034 -3814 241654 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 251274 -3814 251894 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 261514 -3814 262134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 271754 -3814 272374 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 281994 -3814 282614 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 292234 -3814 292854 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 302474 -3814 303094 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 312714 -3814 313334 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 322954 -3814 323574 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 333194 -3814 333814 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 343434 -3814 344054 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 353674 -3814 354294 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 363914 -3814 364534 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 374154 -3814 374774 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 384394 -3814 385014 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 394634 -3814 395254 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 404874 -3814 405494 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 415114 -3814 415734 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 425354 -3814 425974 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 435594 -3814 436214 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 445834 -3814 446454 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 456074 -3814 456694 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 466314 -3814 466934 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 476554 -3814 477174 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 486794 -3814 487414 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 497034 -3814 497654 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 507274 -3814 507894 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 517514 -3814 518134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 527754 -3814 528374 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 537994 -3814 538614 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 15754 -3814 16374 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 25994 657000 26614 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 36234 657000 36854 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 46474 657000 47094 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 56714 657000 57334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 66954 657000 67574 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77194 657000 77814 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 87434 657000 88054 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 97674 657000 98294 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 107914 657000 108534 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 118154 657000 118774 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 128394 657000 129014 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 138634 657000 139254 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 148874 657000 149494 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 159114 657000 159734 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 169354 657000 169974 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 179594 657000 180214 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 189834 657000 190454 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 200074 657000 200694 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 210314 657000 210934 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 220554 657000 221174 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 230794 657000 231414 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 241034 657000 241654 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 251274 657000 251894 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 261514 657000 262134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 271754 657000 272374 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 281994 657000 282614 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 292234 657000 292854 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 302474 657000 303094 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 312714 657000 313334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 322954 657000 323574 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 333194 657000 333814 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 343434 657000 344054 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 353674 657000 354294 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 363914 657000 364534 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 374154 657000 374774 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 384394 657000 385014 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 394634 657000 395254 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 404874 657000 405494 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 415114 657000 415734 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 425354 657000 425974 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 435594 657000 436214 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 445834 657000 446454 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 456074 657000 456694 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 466314 657000 466934 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 476554 657000 477174 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 486794 657000 487414 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 497034 657000 497654 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 507274 657000 507894 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 517514 657000 518134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 527754 657000 528374 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 537994 657000 538614 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 548234 -3814 548854 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 558474 -3814 559094 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 568714 -3814 569334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 578954 -3814 579574 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 19474 -5734 20094 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 29714 -5734 30334 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 39954 -5734 40574 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 50194 -5734 50814 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 60434 -5734 61054 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 70674 -5734 71294 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 80914 -5734 81534 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 91154 -5734 91774 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 101394 -5734 102014 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 111634 -5734 112254 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 121874 -5734 122494 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 132114 -5734 132734 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 142354 -5734 142974 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 152594 -5734 153214 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 162834 -5734 163454 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 173074 -5734 173694 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 183314 -5734 183934 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 193554 -5734 194174 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 203794 -5734 204414 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 214034 -5734 214654 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 224274 -5734 224894 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 234514 -5734 235134 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 244754 -5734 245374 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 254994 -5734 255614 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 265234 -5734 265854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 275474 -5734 276094 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 285714 -5734 286334 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 295954 -5734 296574 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 306194 -5734 306814 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 316434 -5734 317054 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 326674 -5734 327294 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 336914 -5734 337534 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 347154 -5734 347774 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 357394 -5734 358014 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 367634 -5734 368254 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 377874 -5734 378494 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 388114 -5734 388734 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 398354 -5734 398974 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 408594 -5734 409214 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 418834 -5734 419454 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 429074 -5734 429694 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 439314 -5734 439934 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 449554 -5734 450174 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 459794 -5734 460414 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 470034 -5734 470654 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 480274 -5734 480894 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 490514 -5734 491134 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 500754 -5734 501374 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 510994 -5734 511614 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 521234 -5734 521854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 531474 -5734 532094 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 19474 657000 20094 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 29714 657000 30334 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 39954 657000 40574 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 50194 657000 50814 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 60434 657000 61054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 70674 657000 71294 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 80914 657000 81534 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 91154 657000 91774 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 101394 657000 102014 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 111634 657000 112254 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 121874 657000 122494 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 132114 657000 132734 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 142354 657000 142974 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 152594 657000 153214 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 162834 657000 163454 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 173074 657000 173694 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 183314 657000 183934 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 193554 657000 194174 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 203794 657000 204414 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 214034 657000 214654 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 224274 657000 224894 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 234514 657000 235134 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 244754 657000 245374 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 254994 657000 255614 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 265234 657000 265854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 275474 657000 276094 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 285714 657000 286334 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 295954 657000 296574 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 306194 657000 306814 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 316434 657000 317054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 326674 657000 327294 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 336914 657000 337534 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 347154 657000 347774 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 357394 657000 358014 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 367634 657000 368254 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 377874 657000 378494 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 388114 657000 388734 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 398354 657000 398974 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 408594 657000 409214 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 418834 657000 419454 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 429074 657000 429694 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 439314 657000 439934 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 449554 657000 450174 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 459794 657000 460414 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 470034 657000 470654 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 480274 657000 480894 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 490514 657000 491134 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 500754 657000 501374 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 510994 657000 511614 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 521234 657000 521854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 531474 657000 532094 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 541714 -5734 542334 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 551954 -5734 552574 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 562194 -5734 562814 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 572434 -5734 573054 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 23194 -7654 23814 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 33434 -7654 34054 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 43674 -7654 44294 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 53914 -7654 54534 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 64154 -7654 64774 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 74394 -7654 75014 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84634 -7654 85254 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 94874 -7654 95494 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 105114 -7654 105734 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 115354 -7654 115974 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 125594 -7654 126214 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 135834 -7654 136454 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 146074 -7654 146694 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156314 -7654 156934 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 166554 -7654 167174 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 176794 -7654 177414 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 187034 -7654 187654 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 197274 -7654 197894 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 207514 -7654 208134 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 217754 -7654 218374 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 227994 -7654 228614 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 238234 -7654 238854 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 248474 -7654 249094 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 258714 -7654 259334 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 268954 -7654 269574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 279194 -7654 279814 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 289434 -7654 290054 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 299674 -7654 300294 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 309914 -7654 310534 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 320154 -7654 320774 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 330394 -7654 331014 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 340634 -7654 341254 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 350874 -7654 351494 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 361114 -7654 361734 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 371354 -7654 371974 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 381594 -7654 382214 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 391834 -7654 392454 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 402074 -7654 402694 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 412314 -7654 412934 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 422554 -7654 423174 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 432794 -7654 433414 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 443034 -7654 443654 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 453274 -7654 453894 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 463514 -7654 464134 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 473754 -7654 474374 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 483994 -7654 484614 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 494234 -7654 494854 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 504474 -7654 505094 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 514714 -7654 515334 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 524954 -7654 525574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 535194 -7654 535814 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 23194 657000 23814 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 33434 657000 34054 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 43674 657000 44294 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 53914 657000 54534 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 64154 657000 64774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 74394 657000 75014 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84634 657000 85254 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 94874 657000 95494 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 105114 657000 105734 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 115354 657000 115974 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 125594 657000 126214 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 135834 657000 136454 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 146074 657000 146694 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156314 657000 156934 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 166554 657000 167174 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 176794 657000 177414 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 187034 657000 187654 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 197274 657000 197894 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 207514 657000 208134 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 217754 657000 218374 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 227994 657000 228614 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 238234 657000 238854 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 248474 657000 249094 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 258714 657000 259334 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 268954 657000 269574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 279194 657000 279814 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 289434 657000 290054 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 299674 657000 300294 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 309914 657000 310534 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 320154 657000 320774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 330394 657000 331014 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 340634 657000 341254 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 350874 657000 351494 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 361114 657000 361734 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 371354 657000 371974 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 381594 657000 382214 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 391834 657000 392454 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 402074 657000 402694 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 412314 657000 412934 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 422554 657000 423174 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 432794 657000 433414 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 443034 657000 443654 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 453274 657000 453894 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 463514 657000 464134 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 473754 657000 474374 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 483994 657000 484614 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 494234 657000 494854 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 504474 657000 505094 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 514714 657000 515334 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 524954 657000 525574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 535194 657000 535814 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 545434 -7654 546054 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 555674 -7654 556294 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 565914 -7654 566534 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 576154 -7654 576774 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 24594 -5734 25214 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 34834 -5734 35454 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 45074 -5734 45694 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 55314 -5734 55934 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 65554 -5734 66174 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 75794 -5734 76414 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 86034 -5734 86654 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 96274 -5734 96894 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 106514 -5734 107134 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 116754 -5734 117374 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 126994 -5734 127614 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 137234 -5734 137854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 147474 -5734 148094 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 157714 -5734 158334 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 167954 -5734 168574 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 178194 -5734 178814 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 188434 -5734 189054 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 198674 -5734 199294 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 208914 -5734 209534 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 219154 -5734 219774 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 229394 -5734 230014 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 239634 -5734 240254 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 249874 -5734 250494 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 260114 -5734 260734 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 270354 -5734 270974 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 280594 -5734 281214 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 290834 -5734 291454 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 301074 -5734 301694 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 311314 -5734 311934 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 321554 -5734 322174 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 331794 -5734 332414 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 342034 -5734 342654 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 352274 -5734 352894 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 362514 -5734 363134 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 372754 -5734 373374 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 382994 -5734 383614 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 393234 -5734 393854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 403474 -5734 404094 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 413714 -5734 414334 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423954 -5734 424574 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 434194 -5734 434814 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 444434 -5734 445054 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 454674 -5734 455294 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 464914 -5734 465534 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 475154 -5734 475774 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 485394 -5734 486014 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495634 -5734 496254 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 505874 -5734 506494 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 516114 -5734 516734 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 526354 -5734 526974 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 536594 -5734 537214 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 14354 -5734 14974 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 24594 657000 25214 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 34834 657000 35454 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 45074 657000 45694 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 55314 657000 55934 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 65554 657000 66174 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 75794 657000 76414 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 86034 657000 86654 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 96274 657000 96894 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 106514 657000 107134 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 116754 657000 117374 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 126994 657000 127614 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 137234 657000 137854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 147474 657000 148094 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 157714 657000 158334 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 167954 657000 168574 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 178194 657000 178814 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 188434 657000 189054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 198674 657000 199294 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 208914 657000 209534 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 219154 657000 219774 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 229394 657000 230014 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 239634 657000 240254 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 249874 657000 250494 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 260114 657000 260734 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 270354 657000 270974 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 280594 657000 281214 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 290834 657000 291454 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 301074 657000 301694 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 311314 657000 311934 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 321554 657000 322174 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 331794 657000 332414 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 342034 657000 342654 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 352274 657000 352894 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 362514 657000 363134 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 372754 657000 373374 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 382994 657000 383614 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 393234 657000 393854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 403474 657000 404094 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 413714 657000 414334 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423954 657000 424574 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 434194 657000 434814 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 444434 657000 445054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 454674 657000 455294 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 464914 657000 465534 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 475154 657000 475774 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 485394 657000 486014 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495634 657000 496254 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 505874 657000 506494 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 516114 657000 516734 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 526354 657000 526974 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 536594 657000 537214 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 546834 -5734 547454 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 557074 -5734 557694 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567314 -5734 567934 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 577554 -5734 578174 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 18074 -7654 18694 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 28314 -7654 28934 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 38554 -7654 39174 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 48794 -7654 49414 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 59034 -7654 59654 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 69274 -7654 69894 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 79514 -7654 80134 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 89754 -7654 90374 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 99994 -7654 100614 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 110234 -7654 110854 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 120474 -7654 121094 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 130714 -7654 131334 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 140954 -7654 141574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 151194 -7654 151814 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 161434 -7654 162054 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 171674 -7654 172294 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 181914 -7654 182534 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 192154 -7654 192774 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 202394 -7654 203014 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 212634 -7654 213254 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 222874 -7654 223494 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 233114 -7654 233734 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 243354 -7654 243974 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 253594 -7654 254214 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 263834 -7654 264454 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 274074 -7654 274694 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 284314 -7654 284934 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 294554 -7654 295174 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 304794 -7654 305414 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 315034 -7654 315654 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 325274 -7654 325894 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 335514 -7654 336134 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 345754 -7654 346374 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 355994 -7654 356614 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 366234 -7654 366854 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 376474 -7654 377094 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 386714 -7654 387334 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 396954 -7654 397574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 407194 -7654 407814 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 417434 -7654 418054 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 427674 -7654 428294 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 437914 -7654 438534 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 448154 -7654 448774 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 458394 -7654 459014 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 468634 -7654 469254 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 478874 -7654 479494 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 489114 -7654 489734 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 499354 -7654 499974 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 509594 -7654 510214 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 519834 -7654 520454 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 530074 -7654 530694 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 540314 -7654 540934 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 18074 657000 18694 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 28314 657000 28934 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 38554 657000 39174 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 48794 657000 49414 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 59034 657000 59654 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 69274 657000 69894 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 79514 657000 80134 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 89754 657000 90374 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 99994 657000 100614 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 110234 657000 110854 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 120474 657000 121094 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 130714 657000 131334 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 140954 657000 141574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 151194 657000 151814 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 161434 657000 162054 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 171674 657000 172294 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 181914 657000 182534 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 192154 657000 192774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 202394 657000 203014 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 212634 657000 213254 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 222874 657000 223494 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 233114 657000 233734 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 243354 657000 243974 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 253594 657000 254214 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 263834 657000 264454 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 274074 657000 274694 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 284314 657000 284934 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 294554 657000 295174 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 304794 657000 305414 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 315034 657000 315654 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 325274 657000 325894 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 335514 657000 336134 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 345754 657000 346374 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 355994 657000 356614 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 366234 657000 366854 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 376474 657000 377094 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 386714 657000 387334 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 396954 657000 397574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 407194 657000 407814 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 417434 657000 418054 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 427674 657000 428294 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 437914 657000 438534 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 448154 657000 448774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 458394 657000 459014 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 468634 657000 469254 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 478874 657000 479494 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 489114 657000 489734 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 499354 657000 499974 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 509594 657000 510214 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 519834 657000 520454 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 530074 657000 530694 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 540314 657000 540934 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 550554 -7654 551174 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 560794 -7654 561414 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 571034 -7654 571654 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 581274 -7654 581894 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 17154 -1894 17774 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 27394 -1894 28014 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 37634 -1894 38254 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 47874 -1894 48494 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 58114 -1894 58734 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 68354 -1894 68974 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 78594 -1894 79214 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 88834 -1894 89454 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 99074 -1894 99694 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 109314 -1894 109934 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 119554 -1894 120174 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 129794 -1894 130414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 140034 -1894 140654 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 150274 -1894 150894 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 160514 -1894 161134 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 170754 -1894 171374 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 180994 -1894 181614 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 191234 -1894 191854 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 201474 -1894 202094 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 211714 -1894 212334 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 221954 -1894 222574 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 232194 -1894 232814 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 242434 -1894 243054 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 252674 -1894 253294 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 262914 -1894 263534 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 273154 -1894 273774 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 283394 -1894 284014 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 293634 -1894 294254 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 303874 -1894 304494 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 314114 -1894 314734 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 324354 -1894 324974 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 334594 -1894 335214 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 344834 -1894 345454 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 355074 -1894 355694 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 365314 -1894 365934 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 375554 -1894 376174 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 385794 -1894 386414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 396034 -1894 396654 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 406274 -1894 406894 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 416514 -1894 417134 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 426754 -1894 427374 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 436994 -1894 437614 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 447234 -1894 447854 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 457474 -1894 458094 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 467714 -1894 468334 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 477954 -1894 478574 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 488194 -1894 488814 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 498434 -1894 499054 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 508674 -1894 509294 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 518914 -1894 519534 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 529154 -1894 529774 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 539394 -1894 540014 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 6914 -1894 7534 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 17154 657000 17774 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 27394 657000 28014 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 37634 657000 38254 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 47874 657000 48494 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 58114 657000 58734 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 68354 657000 68974 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 78594 657000 79214 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 88834 657000 89454 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 99074 657000 99694 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 109314 657000 109934 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 119554 657000 120174 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 129794 657000 130414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 140034 657000 140654 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 150274 657000 150894 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 160514 657000 161134 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 170754 657000 171374 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 180994 657000 181614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 191234 657000 191854 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 201474 657000 202094 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 211714 657000 212334 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 221954 657000 222574 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 232194 657000 232814 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 242434 657000 243054 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 252674 657000 253294 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 262914 657000 263534 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 273154 657000 273774 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 283394 657000 284014 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 293634 657000 294254 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 303874 657000 304494 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 314114 657000 314734 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 324354 657000 324974 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 334594 657000 335214 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 344834 657000 345454 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 355074 657000 355694 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 365314 657000 365934 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 375554 657000 376174 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 385794 657000 386414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 396034 657000 396654 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 406274 657000 406894 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 416514 657000 417134 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 426754 657000 427374 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 436994 657000 437614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 447234 657000 447854 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 457474 657000 458094 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 467714 657000 468334 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 477954 657000 478574 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 488194 657000 488814 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 498434 657000 499054 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 508674 657000 509294 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 518914 657000 519534 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 529154 657000 529774 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 539394 657000 540014 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 549634 -1894 550254 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559874 -1894 560494 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 570114 -1894 570734 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 580354 -1894 580974 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 20874 -3814 21494 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 31114 -3814 31734 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 41354 -3814 41974 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 51594 -3814 52214 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 61834 -3814 62454 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 72074 -3814 72694 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 82314 -3814 82934 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 92554 -3814 93174 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 102794 -3814 103414 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 113034 -3814 113654 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 123274 -3814 123894 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 133514 -3814 134134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 143754 -3814 144374 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 153994 -3814 154614 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 164234 -3814 164854 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 174474 -3814 175094 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 184714 -3814 185334 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 194954 -3814 195574 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 205194 -3814 205814 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 215434 -3814 216054 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 225674 -3814 226294 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 235914 -3814 236534 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 246154 -3814 246774 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 256394 -3814 257014 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 266634 -3814 267254 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 276874 -3814 277494 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 287114 -3814 287734 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 297354 -3814 297974 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 307594 -3814 308214 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 317834 -3814 318454 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 328074 -3814 328694 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 338314 -3814 338934 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 348554 -3814 349174 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 358794 -3814 359414 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 369034 -3814 369654 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 379274 -3814 379894 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 389514 -3814 390134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 399754 -3814 400374 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 409994 -3814 410614 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 420234 -3814 420854 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 430474 -3814 431094 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 440714 -3814 441334 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 450954 -3814 451574 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 461194 -3814 461814 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 471434 -3814 472054 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 481674 -3814 482294 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491914 -3814 492534 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 502154 -3814 502774 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 512394 -3814 513014 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 522634 -3814 523254 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 532874 -3814 533494 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 10634 -3814 11254 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 20874 657000 21494 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 31114 657000 31734 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 41354 657000 41974 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 51594 657000 52214 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 61834 657000 62454 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 72074 657000 72694 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 82314 657000 82934 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 92554 657000 93174 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 102794 657000 103414 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 113034 657000 113654 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 123274 657000 123894 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 133514 657000 134134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 143754 657000 144374 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 153994 657000 154614 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 164234 657000 164854 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 174474 657000 175094 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 184714 657000 185334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 194954 657000 195574 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 205194 657000 205814 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 215434 657000 216054 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 225674 657000 226294 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 235914 657000 236534 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 246154 657000 246774 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 256394 657000 257014 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 266634 657000 267254 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 276874 657000 277494 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 287114 657000 287734 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 297354 657000 297974 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 307594 657000 308214 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 317834 657000 318454 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 328074 657000 328694 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 338314 657000 338934 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 348554 657000 349174 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 358794 657000 359414 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 369034 657000 369654 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 379274 657000 379894 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 389514 657000 390134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 399754 657000 400374 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 409994 657000 410614 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 420234 657000 420854 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 430474 657000 431094 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 440714 657000 441334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 450954 657000 451574 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 461194 657000 461814 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 471434 657000 472054 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 481674 657000 482294 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491914 657000 492534 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 502154 657000 502774 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 512394 657000 513014 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 522634 657000 523254 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 532874 657000 533494 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 543114 -3814 543734 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 553354 -3814 553974 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563594 -3814 564214 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 573834 -3814 574454 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
