* NGSPICE file created from tile_clb.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_4 abstract view
.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_8 abstract view
.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

.subckt tile_clb bi_u1y0n_L1[0] bi_u1y0n_L1[10] bi_u1y0n_L1[11] bi_u1y0n_L1[1] bi_u1y0n_L1[2]
+ bi_u1y0n_L1[3] bi_u1y0n_L1[4] bi_u1y0n_L1[5] bi_u1y0n_L1[6] bi_u1y0n_L1[7] bi_u1y0n_L1[8]
+ bi_u1y0n_L1[9] bi_u1y0s_L1[0] bi_u1y0s_L1[10] bi_u1y0s_L1[11] bi_u1y0s_L1[1] bi_u1y0s_L1[2]
+ bi_u1y0s_L1[3] bi_u1y0s_L1[4] bi_u1y0s_L1[5] bi_u1y0s_L1[6] bi_u1y0s_L1[7] bi_u1y0s_L1[8]
+ bi_u1y0s_L1[9] clk cu_x0y0n_L1[0] cu_x0y0n_L1[10] cu_x0y0n_L1[11] cu_x0y0n_L1[1]
+ cu_x0y0n_L1[2] cu_x0y0n_L1[3] cu_x0y0n_L1[4] cu_x0y0n_L1[5] cu_x0y0n_L1[6] cu_x0y0n_L1[7]
+ cu_x0y0n_L1[8] cu_x0y0n_L1[9] cu_x0y0s_L1[0] cu_x0y0s_L1[10] cu_x0y0s_L1[11] cu_x0y0s_L1[1]
+ cu_x0y0s_L1[2] cu_x0y0s_L1[3] cu_x0y0s_L1[4] cu_x0y0s_L1[5] cu_x0y0s_L1[6] cu_x0y0s_L1[7]
+ cu_x0y0s_L1[8] cu_x0y0s_L1[9] prog_clk prog_din prog_done prog_dout prog_rst prog_we
+ prog_we_o vccd1 vssd1
XFILLER_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2106_ _2749_/Q _2100_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _2106_/X sky130_fd_sc_hd__o21ba_1
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2037_ _2763_/Q _2037_/B _2037_/C vssd1 vssd1 vccd1 vccd1 _2038_/A sky130_fd_sc_hd__and3_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2939_ _2949_/CLK _2939_/D vssd1 vssd1 vccd1 vccd1 _2939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1606_ _1604_/X _1605_/X _1457_/A vssd1 vssd1 vccd1 vccd1 _1607_/S sky130_fd_sc_hd__o21a_1
X_2655_ _2668_/CLK _2655_/D vssd1 vssd1 vccd1 vccd1 _2655_/Q sky130_fd_sc_hd__dfxtp_1
X_2724_ _2766_/CLK _2724_/D vssd1 vssd1 vccd1 vccd1 _2724_/Q sky130_fd_sc_hd__dfxtp_1
X_1468_ _2909_/Q _2908_/Q _1664_/A _1466_/Y _1467_/Y vssd1 vssd1 vccd1 vccd1 _1468_/X
+ sky130_fd_sc_hd__a311o_2
X_1537_ _2902_/Q _1753_/B _1536_/Y _1661_/X _1598_/B vssd1 vssd1 vccd1 vccd1 _1538_/B
+ sky130_fd_sc_hd__o221a_1
X_2586_ _2931_/Q _2574_/X _2585_/X vssd1 vssd1 vccd1 vccd1 _2928_/D sky130_fd_sc_hd__o21a_1
X_1399_ _2794_/Q _1389_/Y _1396_/X _2791_/Q vssd1 vssd1 vccd1 vccd1 _1399_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2440_ _2872_/Q _2430_/X _2436_/X vssd1 vssd1 vccd1 vccd1 _2440_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1322_ input21/X input3/X _1322_/S vssd1 vssd1 vccd1 vccd1 _1322_/X sky130_fd_sc_hd__mux2_1
X_2371_ _1366_/S _2353_/X _2359_/X vssd1 vssd1 vccd1 vccd1 _2371_/X sky130_fd_sc_hd__o21ba_1
XFILLER_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2707_ _2881_/CLK _2707_/D vssd1 vssd1 vccd1 vccd1 _2707_/Q sky130_fd_sc_hd__dfxtp_1
X_2638_ _1561_/Y _1588_/X _1596_/X _1598_/X _2658_/Q vssd1 vssd1 vccd1 vccd1 _2950_/D
+ sky130_fd_sc_hd__o2111a_1
X_2569_ _2925_/Q _2561_/X _2568_/X vssd1 vssd1 vccd1 vccd1 _2922_/D sky130_fd_sc_hd__o21a_1
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1940_ _2153_/A vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1871_ _2662_/Q _1850_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__o21ba_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2423_ _2866_/Q _2417_/X _2422_/X vssd1 vssd1 vccd1 vccd1 _2423_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2354_ _1322_/S _2353_/X _2345_/X vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__o21ba_1
X_2285_ _2301_/A vssd1 vssd1 vccd1 vccd1 _2285_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2946_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2070_ _2735_/Q _2068_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__o21ba_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1854_ _2657_/Q _1850_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _1854_/X sky130_fd_sc_hd__o21ba_1
X_1923_ _1486_/Y _1861_/X _2639_/A vssd1 vssd1 vccd1 vccd1 _1923_/Y sky130_fd_sc_hd__a21oi_1
X_1785_ _2819_/Q _1783_/Y _2954_/A _1784_/X vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__a31o_1
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2406_ _1377_/S _2397_/X _2405_/X vssd1 vssd1 vccd1 vccd1 _2859_/D sky130_fd_sc_hd__o21a_1
X_2337_ _1384_/S _2324_/X _2332_/X vssd1 vssd1 vccd1 vccd1 _2337_/X sky130_fd_sc_hd__o21ba_1
XFILLER_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2199_ _2783_/Q _2196_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _2199_/X sky130_fd_sc_hd__o21ba_1
X_2268_ _2268_/A vssd1 vssd1 vccd1 vccd1 _2460_/A sky130_fd_sc_hd__buf_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1570_ _1593_/C _1589_/D _1583_/B vssd1 vssd1 vccd1 vccd1 _1570_/Y sky130_fd_sc_hd__o21ai_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2053_ _2053_/A vssd1 vssd1 vccd1 vccd1 _2053_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2122_ _2754_/Q _2110_/X _2121_/X vssd1 vssd1 vccd1 vccd1 _2755_/D sky130_fd_sc_hd__o21a_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2955_ _2955_/A vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1906_ _2675_/Q _1899_/X _1901_/X vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__o21ba_1
X_1837_ _1899_/A vssd1 vssd1 vccd1 vccd1 _1837_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2886_ _2891_/CLK _2886_/D vssd1 vssd1 vccd1 vccd1 _2886_/Q sky130_fd_sc_hd__dfxtp_1
X_1768_ _2783_/Q _2037_/B _1768_/C vssd1 vssd1 vccd1 vccd1 _1769_/A sky130_fd_sc_hd__and3_1
XFILLER_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1699_ _1368_/X _1369_/X _2928_/Q vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput42 _2960_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[10] sky130_fd_sc_hd__clkbuf_1
Xoutput53 _2829_/Q vssd1 vssd1 vccd1 vccd1 prog_dout sky130_fd_sc_hd__clkbuf_1
Xoutput31 _2961_/A vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[11] sky130_fd_sc_hd__clkbuf_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2671_ _2677_/CLK _2671_/D vssd1 vssd1 vccd1 vccd1 _2671_/Q sky130_fd_sc_hd__dfxtp_1
X_2740_ _2755_/CLK _2740_/D vssd1 vssd1 vccd1 vccd1 _2740_/Q sky130_fd_sc_hd__dfxtp_1
X_1622_ _1502_/B input3/X _2873_/Q vssd1 vssd1 vccd1 vccd1 _1622_/X sky130_fd_sc_hd__mux2_1
X_1484_ _1778_/A _1484_/B vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__and2_1
X_1553_ _1502_/B input11/X _1553_/S vssd1 vssd1 vccd1 vccd1 _1553_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2036_ _2722_/Q _2026_/X _2035_/X vssd1 vssd1 vccd1 vccd1 _2723_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2105_ _2747_/Q _2097_/X _2104_/X vssd1 vssd1 vccd1 vccd1 _2748_/D sky130_fd_sc_hd__o21a_1
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2938_ _2943_/CLK _2938_/D vssd1 vssd1 vccd1 vccd1 _2938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2869_ _2872_/CLK _2869_/D vssd1 vssd1 vccd1 vccd1 _2869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xclkbuf_leaf_22_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2948_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2723_ _2881_/CLK _2723_/D vssd1 vssd1 vccd1 vccd1 _2723_/Q sky130_fd_sc_hd__dfxtp_1
X_2654_ _2668_/CLK _2654_/D vssd1 vssd1 vccd1 vccd1 _2654_/Q sky130_fd_sc_hd__dfxtp_1
X_1605_ _2901_/Q _2900_/Q _1605_/C vssd1 vssd1 vccd1 vccd1 _1605_/X sky130_fd_sc_hd__and3b_1
X_1536_ _2903_/Q _2902_/Q vssd1 vssd1 vccd1 vccd1 _1536_/Y sky130_fd_sc_hd__nand2_1
X_2585_ _2928_/Q _2583_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__o21ba_1
X_1467_ _2908_/Q _1467_/B vssd1 vssd1 vccd1 vccd1 _1467_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1398_ _2788_/Q _1391_/Y _1396_/X _2787_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1398_/X
+ sky130_fd_sc_hd__a221o_1
X_2019_ _2715_/Q _2013_/X _2018_/X vssd1 vssd1 vccd1 vccd1 _2716_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1321_ input18/X input9/X _2840_/Q vssd1 vssd1 vccd1 vccd1 _1321_/X sky130_fd_sc_hd__mux2_1
X_2370_ _2384_/A vssd1 vssd1 vccd1 vccd1 _2370_/X sky130_fd_sc_hd__clkbuf_2
X_2706_ _2881_/CLK _2706_/D vssd1 vssd1 vccd1 vccd1 _2706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1519_ _1520_/B _1522_/B vssd1 vssd1 vccd1 vccd1 _1519_/Y sky130_fd_sc_hd__nor2_1
X_2499_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__clkbuf_2
X_2568_ _2922_/Q _2550_/X _2551_/X vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__o21ba_1
X_2637_ _2637_/A vssd1 vssd1 vccd1 vccd1 _2949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1870_ _1927_/A vssd1 vssd1 vccd1 vccd1 _1870_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2353_ _2400_/S vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__clkbuf_2
X_2422_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2284_ _2817_/Q _2282_/X _2283_/X vssd1 vssd1 vccd1 vccd1 _2814_/D sky130_fd_sc_hd__o21a_1
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1999_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1999_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1922_ _2679_/Q _1910_/X _1921_/X vssd1 vssd1 vccd1 vccd1 _2680_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1853_ _2655_/Q _1849_/X _1852_/X vssd1 vssd1 vccd1 vccd1 _2656_/D sky130_fd_sc_hd__o21a_1
X_1784_ _2819_/Q _2818_/Q _2151_/B _1784_/D vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__and4b_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2336_ _2832_/Q _2321_/X _2335_/X vssd1 vssd1 vccd1 vccd1 _2833_/D sky130_fd_sc_hd__o21a_1
X_2405_ _2859_/Q _2404_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _2405_/X sky130_fd_sc_hd__o21ba_1
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2198_ _2254_/A vssd1 vssd1 vccd1 vccd1 _2198_/X sky130_fd_sc_hd__clkbuf_1
X_2267_ _2510_/A vssd1 vssd1 vccd1 vccd1 _2268_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2052_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2052_/X sky130_fd_sc_hd__clkbuf_2
X_2121_ _2755_/Q _2113_/X _2114_/X vssd1 vssd1 vccd1 vccd1 _2121_/X sky130_fd_sc_hd__o21ba_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1905_ _2673_/Q _1896_/X _1904_/X vssd1 vssd1 vccd1 vccd1 _2674_/D sky130_fd_sc_hd__o21a_1
X_2885_ _2943_/CLK _2885_/D vssd1 vssd1 vccd1 vccd1 _2885_/Q sky130_fd_sc_hd__dfxtp_1
X_2954_ _2954_/A vssd1 vssd1 vccd1 vccd1 _2954_/X sky130_fd_sc_hd__clkbuf_1
X_1836_ _2614_/A vssd1 vssd1 vccd1 vccd1 _1899_/A sky130_fd_sc_hd__buf_2
X_1698_ _2928_/Q _1698_/B vssd1 vssd1 vccd1 vccd1 _1698_/X sky130_fd_sc_hd__and2_1
X_1767_ _1756_/X _1761_/X _1767_/S vssd1 vssd1 vccd1 vccd1 _1768_/C sky130_fd_sc_hd__mux2_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2319_ _2464_/A _2830_/Q vssd1 vssd1 vccd1 vccd1 _2364_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput43 _2961_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[11] sky130_fd_sc_hd__clkbuf_1
Xoutput54 _2881_/Q vssd1 vssd1 vccd1 vccd1 prog_we_o sky130_fd_sc_hd__clkbuf_1
Xoutput32 _2954_/A vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[1] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2670_ _2677_/CLK _2670_/D vssd1 vssd1 vccd1 vccd1 _2670_/Q sky130_fd_sc_hd__dfxtp_1
X_1552_ _1548_/Y _1549_/X _1551_/X vssd1 vssd1 vccd1 vccd1 _1552_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1621_ _2874_/Q vssd1 vssd1 vccd1 vccd1 _1621_/Y sky130_fd_sc_hd__inv_2
X_1483_ _2723_/Q _1424_/Y _2682_/Q _1482_/X vssd1 vssd1 vccd1 vccd1 _1484_/B sky130_fd_sc_hd__a31o_1
X_2104_ _2748_/Q _2100_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _2104_/X sky130_fd_sc_hd__o21ba_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2035_ _2723_/Q _2022_/X _2023_/X vssd1 vssd1 vccd1 vccd1 _2035_/X sky130_fd_sc_hd__o21ba_1
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2868_ _2872_/CLK _2868_/D vssd1 vssd1 vccd1 vccd1 _2868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2937_ _2937_/CLK _2937_/D vssd1 vssd1 vccd1 vccd1 _2937_/Q sky130_fd_sc_hd__dfxtp_1
X_1819_ _1849_/A vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2799_ _2872_/CLK _2799_/D vssd1 vssd1 vccd1 vccd1 _2799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2722_ _2914_/CLK _2722_/D vssd1 vssd1 vccd1 vccd1 _2722_/Q sky130_fd_sc_hd__dfxtp_2
X_2653_ _2668_/CLK _2653_/D vssd1 vssd1 vccd1 vccd1 _2653_/Q sky130_fd_sc_hd__dfxtp_1
X_1604_ _1547_/Y _1617_/A _1617_/B _1603_/X _2901_/Q vssd1 vssd1 vccd1 vccd1 _1604_/X
+ sky130_fd_sc_hd__o311a_1
X_1535_ _1531_/X _1534_/X _2839_/Q vssd1 vssd1 vccd1 vccd1 _1753_/B sky130_fd_sc_hd__mux2_4
X_2584_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1466_ _2908_/Q _1380_/B _2909_/Q vssd1 vssd1 vccd1 vccd1 _1466_/Y sky130_fd_sc_hd__a21oi_1
X_1397_ _2790_/Q _1389_/Y _1390_/Y _2789_/Q vssd1 vssd1 vccd1 vccd1 _1397_/X sky130_fd_sc_hd__a22o_1
X_2018_ _2716_/Q _2008_/X _2009_/X vssd1 vssd1 vccd1 vccd1 _2018_/X sky130_fd_sc_hd__o21ba_1
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1320_ _1322_/S input6/X vssd1 vssd1 vccd1 vccd1 _1320_/X sky130_fd_sc_hd__and2_1
X_2705_ _2881_/CLK _2705_/D vssd1 vssd1 vccd1 vccd1 _2705_/Q sky130_fd_sc_hd__dfxtp_1
X_2636_ _2268_/A _2827_/Q vssd1 vssd1 vccd1 vccd1 _2637_/A sky130_fd_sc_hd__and2b_1
X_1518_ _1598_/B _1520_/B _1522_/B vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__and3_1
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2567_ _2920_/Q _2561_/X _2566_/Y vssd1 vssd1 vccd1 vccd1 _2921_/D sky130_fd_sc_hd__o21a_1
X_2498_ _2894_/Q _2492_/X _2497_/X vssd1 vssd1 vccd1 vccd1 _2895_/D sky130_fd_sc_hd__o21a_1
X_1449_ _2856_/Q _1449_/B input5/X vssd1 vssd1 vccd1 vccd1 _1449_/X sky130_fd_sc_hd__and3b_1
XFILLER_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2352_ _2384_/A vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2421_ _1315_/S _2412_/X _2420_/X vssd1 vssd1 vccd1 vccd1 _2865_/D sky130_fd_sc_hd__o21a_1
X_2283_ _2814_/Q _2264_/X _2277_/X vssd1 vssd1 vccd1 vccd1 _2283_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1998_ _2707_/Q _1985_/X _1997_/X vssd1 vssd1 vccd1 vccd1 _2708_/D sky130_fd_sc_hd__o21a_1
XFILLER_69_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2619_ _2940_/Q _2611_/X _2618_/X vssd1 vssd1 vccd1 vccd1 _2941_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1921_ _2680_/Q _1915_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _1921_/X sky130_fd_sc_hd__o21ba_1
X_1852_ _2656_/Q _1850_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _1852_/X sky130_fd_sc_hd__o21ba_1
X_1783_ _2818_/Q vssd1 vssd1 vccd1 vccd1 _1783_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2335_ _2833_/Q _2324_/X _2332_/X vssd1 vssd1 vccd1 vccd1 _2335_/X sky130_fd_sc_hd__o21ba_1
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2404_ _2430_/A vssd1 vssd1 vccd1 vccd1 _2404_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2266_ _2811_/Q _2262_/X _2265_/X vssd1 vssd1 vccd1 vccd1 _2808_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2197_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2254_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_16_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2931_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2120_ _2753_/Q _2110_/X _2119_/X vssd1 vssd1 vccd1 vccd1 _2754_/D sky130_fd_sc_hd__o21a_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2051_ _2728_/Q _2039_/X _2050_/X vssd1 vssd1 vccd1 vccd1 _2729_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1904_ _2674_/Q _1899_/X _1901_/X vssd1 vssd1 vccd1 vccd1 _1904_/X sky130_fd_sc_hd__o21ba_1
X_2953_ _2960_/A vssd1 vssd1 vccd1 vccd1 _2953_/X sky130_fd_sc_hd__clkbuf_1
X_1835_ _2482_/A vssd1 vssd1 vccd1 vccd1 _2614_/A sky130_fd_sc_hd__clkbuf_2
X_2884_ _2943_/CLK _2884_/D vssd1 vssd1 vccd1 vccd1 _2884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1697_ _1697_/A vssd1 vssd1 vccd1 vccd1 _2037_/B sky130_fd_sc_hd__clkbuf_2
X_1766_ _2933_/Q _1763_/Y _1764_/X _1765_/X vssd1 vssd1 vccd1 vccd1 _1767_/S sky130_fd_sc_hd__a31o_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2249_ _2802_/Q _2240_/X _2241_/X vssd1 vssd1 vccd1 vccd1 _2249_/X sky130_fd_sc_hd__o21ba_1
X_2318_ _2318_/A vssd1 vssd1 vccd1 vccd1 _2827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput44 _2954_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[1] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput33 _1792_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_63_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1482_ _2723_/Q _2722_/Q _1925_/B vssd1 vssd1 vccd1 vccd1 _1482_/X sky130_fd_sc_hd__and3b_2
X_1620_ _1616_/Y _2892_/Q _1451_/X _1619_/X vssd1 vssd1 vccd1 vccd1 _1657_/S sky130_fd_sc_hd__a31oi_4
X_1551_ _1553_/S _1551_/B _2832_/Q vssd1 vssd1 vccd1 vccd1 _1551_/X sky130_fd_sc_hd__and3b_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2103_ _2746_/Q _2097_/X _2102_/X vssd1 vssd1 vccd1 vccd1 _2747_/D sky130_fd_sc_hd__o21a_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ _2721_/Q _2026_/X _2033_/Y vssd1 vssd1 vccd1 vccd1 _2722_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_prog_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_1818_ _2644_/Q _1802_/X _1817_/X vssd1 vssd1 vccd1 vccd1 _2645_/D sky130_fd_sc_hd__o21a_1
X_2798_ _2872_/CLK _2798_/D vssd1 vssd1 vccd1 vccd1 _2798_/Q sky130_fd_sc_hd__dfxtp_1
X_2867_ _2872_/CLK _2867_/D vssd1 vssd1 vccd1 vccd1 _2867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2936_ _2937_/CLK _2936_/D vssd1 vssd1 vccd1 vccd1 _2936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1749_ _2774_/Q _1747_/X _1748_/X _2772_/Q vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2721_ _2721_/CLK _2721_/D vssd1 vssd1 vccd1 vccd1 _2721_/Q sky130_fd_sc_hd__dfxtp_1
X_2652_ _2668_/CLK _2652_/D vssd1 vssd1 vccd1 vccd1 _2652_/Q sky130_fd_sc_hd__dfxtp_1
X_1603_ _2900_/Q _1764_/B vssd1 vssd1 vccd1 vccd1 _1603_/X sky130_fd_sc_hd__or2_1
X_1465_ _1661_/X vssd1 vssd1 vccd1 vccd1 _1664_/A sky130_fd_sc_hd__inv_2
X_1534_ _1532_/X _1533_/X _2838_/Q vssd1 vssd1 vccd1 vccd1 _1534_/X sky130_fd_sc_hd__mux2_1
X_2583_ _2614_/A vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__clkbuf_2
X_2017_ _2714_/Q _2013_/X _2016_/X vssd1 vssd1 vccd1 vccd1 _2715_/D sky130_fd_sc_hd__o21a_1
X_1396_ _1396_/A _1396_/B vssd1 vssd1 vccd1 vccd1 _1396_/X sky130_fd_sc_hd__and2_1
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2919_ _2931_/CLK _2919_/D vssd1 vssd1 vccd1 vccd1 _2919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2704_ _2881_/CLK _2704_/D vssd1 vssd1 vccd1 vccd1 _2704_/Q sky130_fd_sc_hd__dfxtp_1
X_2635_ _2635_/A vssd1 vssd1 vccd1 vccd1 _2948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2566_ _1673_/Y _2542_/X _2510_/X vssd1 vssd1 vccd1 vccd1 _2566_/Y sky130_fd_sc_hd__a21oi_1
X_1517_ _1581_/A _1517_/B _1516_/X vssd1 vssd1 vccd1 vccd1 _1522_/B sky130_fd_sc_hd__or3b_2
X_2497_ _2895_/Q _2483_/X _2484_/X vssd1 vssd1 vccd1 vccd1 _2497_/X sky130_fd_sc_hd__o21ba_1
X_1448_ input17/X input9/X _2855_/Q vssd1 vssd1 vccd1 vccd1 _1448_/X sky130_fd_sc_hd__mux2_1
X_1379_ _1375_/X _1376_/X _1377_/X _1378_/X _2859_/Q _2860_/Q vssd1 vssd1 vccd1 vccd1
+ _1380_/B sky130_fd_sc_hd__mux4_2
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2420_ _2865_/Q _2417_/X _2409_/X vssd1 vssd1 vccd1 vccd1 _2420_/X sky130_fd_sc_hd__o21ba_1
X_2351_ _2838_/Q _2339_/X _2350_/X vssd1 vssd1 vccd1 vccd1 _2839_/D sky130_fd_sc_hd__o21a_1
XFILLER_43_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2282_ _2296_/A vssd1 vssd1 vccd1 vccd1 _2282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1997_ _2708_/Q _1995_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__o21ba_1
XFILLER_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2549_ _2917_/Q _2545_/X _2548_/X vssd1 vssd1 vccd1 vccd1 _2914_/D sky130_fd_sc_hd__o21a_1
X_2618_ _2941_/Q _2614_/X _2615_/X vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__o21ba_1
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1920_ _2678_/Q _1910_/X _1919_/X vssd1 vssd1 vccd1 vccd1 _2679_/D sky130_fd_sc_hd__o21a_1
X_1851_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1851_/X sky130_fd_sc_hd__clkbuf_1
X_1782_ _1780_/Y _1781_/X _1420_/A vssd1 vssd1 vccd1 vccd1 _1782_/Y sky130_fd_sc_hd__a21oi_2
X_2403_ _2863_/Q _2397_/X _2402_/X vssd1 vssd1 vccd1 vccd1 _2858_/D sky130_fd_sc_hd__o21a_1
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2334_ _1553_/S _2321_/X _2333_/X vssd1 vssd1 vccd1 vccd1 _2832_/D sky130_fd_sc_hd__o21a_1
X_2196_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2196_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2265_ _2808_/Q _2264_/X _2254_/X vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__o21ba_1
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2050_ _2729_/Q _2040_/X _2041_/X vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__o21ba_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2952_ _2961_/A vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1903_ _2672_/Q _1896_/X _1902_/X vssd1 vssd1 vccd1 vccd1 _2673_/D sky130_fd_sc_hd__o21a_1
X_1834_ _1849_/A vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1765_ _2933_/Q _2932_/Q _1765_/C vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__and3b_1
X_2883_ _2937_/CLK _2883_/D vssd1 vssd1 vccd1 vccd1 _2883_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _1667_/X _1686_/X _1695_/X _2741_/Q _1778_/A vssd1 vssd1 vccd1 vccd1 _1983_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2179_ _2775_/Q _2167_/X _2178_/X vssd1 vssd1 vccd1 vccd1 _2776_/D sky130_fd_sc_hd__o21a_1
X_2248_ _2477_/A vssd1 vssd1 vccd1 vccd1 _2248_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2317_ _2313_/X _2317_/B vssd1 vssd1 vccd1 vccd1 _2318_/A sky130_fd_sc_hd__and2b_1
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput34 _2955_/A vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_56_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput45 _1779_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1481_ _2720_/Q _1731_/A _1481_/C vssd1 vssd1 vccd1 vccd1 _1925_/B sky130_fd_sc_hd__and3_1
X_1550_ _2831_/Q vssd1 vssd1 vccd1 vccd1 _1553_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_2033_ _1424_/Y _1861_/X _1972_/X vssd1 vssd1 vccd1 vccd1 _2033_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_1_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2947_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2102_ _2747_/Q _2100_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__o21ba_1
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2935_ _2951_/CLK _2935_/D vssd1 vssd1 vccd1 vccd1 _2935_/Q sky130_fd_sc_hd__dfxtp_1
X_1817_ _2645_/Q _1805_/X _1808_/X vssd1 vssd1 vccd1 vccd1 _1817_/X sky130_fd_sc_hd__o21ba_1
X_2866_ _2866_/CLK _2866_/D vssd1 vssd1 vccd1 vccd1 _2866_/Q sky130_fd_sc_hd__dfxtp_1
X_2797_ _2872_/CLK _2797_/D vssd1 vssd1 vccd1 vccd1 _2797_/Q sky130_fd_sc_hd__dfxtp_1
X_1748_ _1746_/B _1748_/B vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__and2b_1
X_1679_ _2729_/Q _2730_/Q _2731_/Q _2732_/Q _1672_/X _1692_/B vssd1 vssd1 vccd1 vccd1
+ _1679_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2720_ _2721_/CLK _2720_/D vssd1 vssd1 vccd1 vccd1 _2720_/Q sky130_fd_sc_hd__dfxtp_1
X_1602_ _2659_/Q _2950_/Q _2660_/Q vssd1 vssd1 vccd1 vccd1 _1617_/B sky130_fd_sc_hd__and3b_1
X_2651_ _2668_/CLK _2651_/D vssd1 vssd1 vccd1 vccd1 _2651_/Q sky130_fd_sc_hd__dfxtp_1
X_2582_ _2926_/Q _2574_/X _2581_/X vssd1 vssd1 vccd1 vccd1 _2927_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1464_ _2705_/Q _1455_/Y _1460_/X _1476_/A vssd1 vssd1 vccd1 vccd1 _1464_/X sky130_fd_sc_hd__a211o_1
X_1533_ _1530_/B _1533_/B vssd1 vssd1 vccd1 vccd1 _1533_/X sky130_fd_sc_hd__and2b_1
X_1395_ _1328_/Y _1373_/X _1388_/X _1394_/X vssd1 vssd1 vccd1 vccd1 _1395_/X sky130_fd_sc_hd__o211a_1
X_2016_ _2715_/Q _2008_/X _2009_/X vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__o21ba_1
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2918_ _2923_/CLK _2918_/D vssd1 vssd1 vccd1 vccd1 _2918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2849_ _2866_/CLK _2849_/D vssd1 vssd1 vccd1 vccd1 _2849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1516_ _2904_/Q _1514_/X _1515_/Y _2955_/A vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__o22a_1
X_2565_ _2923_/Q _2561_/X _2564_/X vssd1 vssd1 vccd1 vccd1 _2920_/D sky130_fd_sc_hd__o21a_1
X_2703_ _2766_/CLK _2703_/D vssd1 vssd1 vccd1 vccd1 _2703_/Q sky130_fd_sc_hd__dfxtp_1
X_2634_ _2268_/A _2634_/B vssd1 vssd1 vccd1 vccd1 _2635_/A sky130_fd_sc_hd__and2b_1
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2496_ _2897_/Q _2492_/X _2495_/Y vssd1 vssd1 vccd1 vccd1 _2894_/D sky130_fd_sc_hd__o21a_1
X_1447_ _1442_/Y _1444_/X _1445_/X _1446_/Y vssd1 vssd1 vccd1 vccd1 _1451_/A sky130_fd_sc_hd__a211o_1
X_1378_ _1377_/S _1624_/B vssd1 vssd1 vccd1 vccd1 _1378_/X sky130_fd_sc_hd__and2b_1
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2350_ _2839_/Q _2340_/X _2345_/X vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__o21ba_1
X_2281_ _2812_/Q _2262_/X _2280_/X vssd1 vssd1 vccd1 vccd1 _2813_/D sky130_fd_sc_hd__o21a_1
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1996_ _2041_/A vssd1 vssd1 vccd1 vccd1 _1996_/X sky130_fd_sc_hd__clkbuf_1
X_2548_ _2914_/Q _2532_/X _2533_/X vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__o21ba_1
X_2617_ _2943_/Q _2611_/X _2616_/X vssd1 vssd1 vccd1 vccd1 _2940_/D sky130_fd_sc_hd__o21a_1
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2479_ _2891_/Q _2477_/X _2478_/X vssd1 vssd1 vccd1 vccd1 _2888_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1850_ _1899_/A vssd1 vssd1 vccd1 vccd1 _1850_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1781_ _2816_/Q _1794_/B _2817_/Q vssd1 vssd1 vccd1 vccd1 _1781_/X sky130_fd_sc_hd__or3b_1
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2333_ _2832_/Q _2324_/X _2332_/X vssd1 vssd1 vccd1 vccd1 _2333_/X sky130_fd_sc_hd__o21ba_1
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2402_ _1377_/S _2387_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _2402_/X sky130_fd_sc_hd__o21ba_1
X_2195_ _2781_/Q _2193_/X _2194_/X vssd1 vssd1 vccd1 vccd1 _2782_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2264_ _2301_/A vssd1 vssd1 vccd1 vccd1 _2264_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1979_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xclkbuf_leaf_25_prog_clk clkbuf_2_0_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2943_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1902_ _2673_/Q _1899_/X _1901_/X vssd1 vssd1 vccd1 vccd1 _1902_/X sky130_fd_sc_hd__o21ba_1
X_2951_ _2951_/CLK _2951_/D vssd1 vssd1 vccd1 vccd1 _2951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1833_ _2649_/Q _1819_/X _1832_/X vssd1 vssd1 vccd1 vccd1 _2650_/D sky130_fd_sc_hd__o21a_1
X_1764_ _2932_/Q _1764_/B vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__or2_1
X_2882_ _2943_/CLK _2882_/D vssd1 vssd1 vccd1 vccd1 _2882_/Q sky130_fd_sc_hd__dfxtp_1
X_1695_ _1686_/S _1687_/X _1688_/Y _1694_/X _2269_/A vssd1 vssd1 vccd1 vccd1 _1695_/X
+ sky130_fd_sc_hd__a2111o_1
X_2316_ _2316_/A vssd1 vssd1 vccd1 vccd1 _2826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2178_ _2776_/Q _2170_/X _2171_/X vssd1 vssd1 vccd1 vccd1 _2178_/X sky130_fd_sc_hd__o21ba_1
X_2247_ _2800_/Q _2235_/X _2246_/X vssd1 vssd1 vccd1 vccd1 _2801_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput46 _2955_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[3] sky130_fd_sc_hd__clkbuf_1
Xoutput35 _2952_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[4] sky130_fd_sc_hd__clkbuf_1
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1480_ _1464_/X _1468_/X _1473_/X _1476_/X _1479_/X vssd1 vssd1 vccd1 vccd1 _1481_/C
+ sky130_fd_sc_hd__a32o_1
X_2032_ _2720_/Q _2026_/X _2031_/X vssd1 vssd1 vccd1 vccd1 _2721_/D sky130_fd_sc_hd__o21a_1
X_2101_ _2114_/A vssd1 vssd1 vccd1 vccd1 _2101_/X sky130_fd_sc_hd__clkbuf_1
X_2934_ _2951_/CLK _2934_/D vssd1 vssd1 vccd1 vccd1 _2934_/Q sky130_fd_sc_hd__dfxtp_1
X_2865_ _2866_/CLK _2865_/D vssd1 vssd1 vccd1 vccd1 _2865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1678_ _1689_/A vssd1 vssd1 vccd1 vccd1 _1692_/B sky130_fd_sc_hd__clkbuf_2
X_1816_ _2643_/Q _1802_/X _1815_/X vssd1 vssd1 vccd1 vccd1 _2644_/D sky130_fd_sc_hd__o21a_1
X_2796_ _2872_/CLK _2796_/D vssd1 vssd1 vccd1 vccd1 _2796_/Q sky130_fd_sc_hd__dfxtp_1
X_1747_ _1747_/A _1747_/B _1747_/C vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__and3_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1601_ _1561_/Y _1588_/X _1596_/X _1598_/X _1600_/X vssd1 vssd1 vccd1 vccd1 _1617_/A
+ sky130_fd_sc_hd__o2111a_2
X_2650_ _2839_/CLK _2650_/D vssd1 vssd1 vccd1 vccd1 _2650_/Q sky130_fd_sc_hd__dfxtp_1
X_1532_ input21/X input12/X _2837_/Q vssd1 vssd1 vccd1 vccd1 _1532_/X sky130_fd_sc_hd__mux2_1
X_2581_ _2927_/Q _2570_/X _2571_/X vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__o21ba_1
XFILLER_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1463_ _1461_/X _1462_/X _2911_/Q vssd1 vssd1 vccd1 vccd1 _1476_/A sky130_fd_sc_hd__mux2_2
X_1394_ _2798_/Q _1389_/Y _1392_/X _1393_/X vssd1 vssd1 vccd1 vccd1 _1394_/X sky130_fd_sc_hd__a211o_1
X_2015_ _2713_/Q _2013_/X _2014_/X vssd1 vssd1 vccd1 vccd1 _2714_/D sky130_fd_sc_hd__o21a_1
X_2917_ _2923_/CLK _2917_/D vssd1 vssd1 vccd1 vccd1 _2917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2848_ _2858_/CLK _2848_/D vssd1 vssd1 vccd1 vccd1 _2848_/Q sky130_fd_sc_hd__dfxtp_1
X_2779_ _2781_/CLK _2779_/D vssd1 vssd1 vccd1 vccd1 _2779_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2702_ _2881_/CLK _2702_/D vssd1 vssd1 vccd1 vccd1 _2702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1515_ _2905_/Q _2904_/Q vssd1 vssd1 vccd1 vccd1 _1515_/Y sky130_fd_sc_hd__nand2_1
X_2495_ _1487_/Y _2090_/X _2293_/X vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__a21oi_1
X_2564_ _2920_/Q _2550_/X _2551_/X vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__o21ba_1
X_2633_ _2948_/Q input25/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2634_/B sky130_fd_sc_hd__mux2_1
X_1446_ _2857_/Q vssd1 vssd1 vccd1 vccd1 _1446_/Y sky130_fd_sc_hd__inv_2
X_1377_ _1337_/B input3/X _1377_/S vssd1 vssd1 vccd1 vccd1 _1377_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2280_ _2813_/Q _2264_/X _2277_/X vssd1 vssd1 vccd1 vccd1 _2280_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1995_ _2053_/A vssd1 vssd1 vccd1 vccd1 _1995_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2616_ _2940_/Q _2614_/X _2615_/X vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__o21ba_1
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2547_ _2912_/Q _2545_/X _2546_/Y vssd1 vssd1 vccd1 vccd1 _2913_/D sky130_fd_sc_hd__o21a_1
X_1429_ _2744_/Q _1427_/Y _2703_/Q _1428_/X vssd1 vssd1 vccd1 vccd1 _1430_/B sky130_fd_sc_hd__a31o_2
X_2478_ _2888_/Q _2469_/X _2470_/X vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__o21ba_1
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1780_ _2817_/Q _2816_/Q _1793_/C vssd1 vssd1 vccd1 vccd1 _1780_/Y sky130_fd_sc_hd__nand3b_1
X_2332_ _2345_/A vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__clkbuf_1
X_2401_ _2460_/A _2401_/B vssd1 vssd1 vccd1 vccd1 _2857_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2194_ _2782_/Q _2183_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _2194_/X sky130_fd_sc_hd__o21ba_1
X_2263_ _2464_/A _2809_/Q vssd1 vssd1 vccd1 vccd1 _2301_/A sky130_fd_sc_hd__and2_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1978_ _2807_/Q vssd1 vssd1 vccd1 vccd1 _2276_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2881_ _2881_/CLK _2881_/D vssd1 vssd1 vccd1 vccd1 _2881_/Q sky130_fd_sc_hd__dfxtp_1
X_1901_ _1960_/A vssd1 vssd1 vccd1 vccd1 _1901_/X sky130_fd_sc_hd__clkbuf_1
X_2950_ _2950_/CLK _2950_/D vssd1 vssd1 vccd1 vccd1 _2950_/Q sky130_fd_sc_hd__dfxtp_1
X_1832_ _2650_/Q _1820_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1832_/X sky130_fd_sc_hd__o21ba_1
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1694_ _1683_/X _1684_/X _1691_/X _1693_/X _1697_/A vssd1 vssd1 vccd1 vccd1 _1694_/X
+ sky130_fd_sc_hd__o221a_1
X_1763_ _2932_/Q _1794_/B vssd1 vssd1 vccd1 vccd1 _1763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2315_ _2313_/X _2315_/B vssd1 vssd1 vccd1 vccd1 _2316_/A sky130_fd_sc_hd__and2b_1
X_2246_ _2801_/Q _2240_/X _2241_/X vssd1 vssd1 vccd1 vccd1 _2246_/X sky130_fd_sc_hd__o21ba_1
XFILLER_65_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2177_ _2774_/Q _2167_/X _2176_/X vssd1 vssd1 vccd1 vccd1 _2775_/D sky130_fd_sc_hd__o21a_1
XFILLER_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput47 _2956_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[4] sky130_fd_sc_hd__clkbuf_1
Xoutput36 _2953_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2100_ _2126_/A vssd1 vssd1 vccd1 vccd1 _2100_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2031_ _2721_/Q _2022_/X _2023_/X vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__o21ba_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1815_ _2644_/Q _1805_/X _1808_/X vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__o21ba_1
X_2933_ _2933_/CLK _2933_/D vssd1 vssd1 vccd1 vccd1 _2933_/Q sky130_fd_sc_hd__dfxtp_1
X_2795_ _2872_/CLK _2795_/D vssd1 vssd1 vccd1 vccd1 _2795_/Q sky130_fd_sc_hd__dfxtp_1
X_2864_ _2875_/CLK _2864_/D vssd1 vssd1 vccd1 vccd1 _2864_/Q sky130_fd_sc_hd__dfxtp_1
X_1677_ _1743_/A _1677_/B vssd1 vssd1 vccd1 vccd1 _1689_/A sky130_fd_sc_hd__and2_1
X_1746_ _1748_/B _1746_/B vssd1 vssd1 vccd1 vccd1 _1746_/Y sky130_fd_sc_hd__nor2_1
X_2229_ _2794_/Q _2227_/X _2228_/X vssd1 vssd1 vccd1 vccd1 _2229_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1462_ _1613_/B _2955_/A _2910_/Q vssd1 vssd1 vccd1 vccd1 _1462_/X sky130_fd_sc_hd__mux2_1
X_1600_ _1600_/A _2659_/Q vssd1 vssd1 vccd1 vccd1 _1600_/X sky130_fd_sc_hd__and2_2
X_1531_ _2838_/Q _1529_/X _1530_/X vssd1 vssd1 vccd1 vccd1 _1531_/X sky130_fd_sc_hd__a21o_1
X_2580_ _2929_/Q _2574_/X _2579_/X vssd1 vssd1 vccd1 vccd1 _2926_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1393_ _2795_/Q _1396_/A _1396_/B _1328_/A vssd1 vssd1 vccd1 vccd1 _1393_/X sky130_fd_sc_hd__a31o_1
X_2014_ _2714_/Q _2008_/X _2009_/X vssd1 vssd1 vccd1 vccd1 _2014_/X sky130_fd_sc_hd__o21ba_1
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2916_ _2931_/CLK _2916_/D vssd1 vssd1 vccd1 vccd1 _2916_/Q sky130_fd_sc_hd__dfxtp_1
X_2847_ _2858_/CLK _2847_/D vssd1 vssd1 vccd1 vccd1 _2847_/Q sky130_fd_sc_hd__dfxtp_1
X_2778_ _2781_/CLK _2778_/D vssd1 vssd1 vccd1 vccd1 _2778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1729_ _2925_/Q _2924_/Q vssd1 vssd1 vccd1 vccd1 _1729_/Y sky130_fd_sc_hd__nand2_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_prog_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2701_ _2881_/CLK _2701_/D vssd1 vssd1 vccd1 vccd1 _2701_/Q sky130_fd_sc_hd__dfxtp_2
X_2632_ _2946_/Q _2639_/B _2631_/X vssd1 vssd1 vccd1 vccd1 _2947_/D sky130_fd_sc_hd__o21a_1
X_2563_ _2918_/Q _2561_/X _2562_/X vssd1 vssd1 vccd1 vccd1 _2919_/D sky130_fd_sc_hd__o21a_1
X_2494_ _2892_/Q _2492_/X _2493_/X vssd1 vssd1 vccd1 vccd1 _2893_/D sky130_fd_sc_hd__o21a_1
X_1514_ _1514_/A _1514_/B vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__and2_2
X_1445_ _1449_/B _1551_/B _2856_/Q vssd1 vssd1 vccd1 vccd1 _1445_/X sky130_fd_sc_hd__and3b_1
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1376_ input20/X input11/X _2858_/Q vssd1 vssd1 vccd1 vccd1 _1376_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_19_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2765_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _2212_/A vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2615_ _2615_/A vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__clkbuf_1
X_2546_ _1425_/Y _2542_/X _2510_/X vssd1 vssd1 vccd1 vccd1 _2546_/Y sky130_fd_sc_hd__a21oi_1
X_1428_ _2744_/Q _2743_/Q _1983_/C vssd1 vssd1 vccd1 vccd1 _1428_/X sky130_fd_sc_hd__and3b_2
X_2477_ _2477_/A vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1359_ _1356_/B _1551_/B vssd1 vssd1 vccd1 vccd1 _1359_/X sky130_fd_sc_hd__and2b_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2400_ _1446_/Y _1442_/Y _2400_/S vssd1 vssd1 vccd1 vccd1 _2401_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2331_ _2836_/Q _2321_/X _2330_/X vssd1 vssd1 vccd1 vccd1 _2831_/D sky130_fd_sc_hd__o21a_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2262_ _2296_/A vssd1 vssd1 vccd1 vccd1 _2262_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2193_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2193_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1977_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2529_ _2907_/Q _2518_/X _2520_/X vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__o21ba_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1900_ _2615_/A vssd1 vssd1 vccd1 vccd1 _1960_/A sky130_fd_sc_hd__clkbuf_2
X_1831_ _2648_/Q _1819_/X _1830_/X vssd1 vssd1 vccd1 vccd1 _2649_/D sky130_fd_sc_hd__o21a_1
X_2880_ _2949_/CLK _2880_/D vssd1 vssd1 vccd1 vccd1 _2880_/Q sky130_fd_sc_hd__dfxtp_1
X_1693_ _2740_/Q _1672_/X _1692_/B _1692_/X vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__a31o_1
X_1762_ _1762_/A vssd1 vssd1 vccd1 vccd1 _1794_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2314_ _2882_/Q _2826_/Q _2314_/S vssd1 vssd1 vccd1 vccd1 _2315_/B sky130_fd_sc_hd__mux2_1
X_2176_ _2775_/Q _2170_/X _2171_/X vssd1 vssd1 vccd1 vccd1 _2176_/X sky130_fd_sc_hd__o21ba_1
X_2245_ _2799_/Q _2235_/X _2244_/X vssd1 vssd1 vccd1 vccd1 _2800_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput48 _2957_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[5] sky130_fd_sc_hd__clkbuf_1
Xoutput37 _2958_/A vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2030_ _2719_/Q _2026_/X _2029_/X vssd1 vssd1 vccd1 vccd1 _2720_/D sky130_fd_sc_hd__o21a_1
XFILLER_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2932_ _2933_/CLK _2932_/D vssd1 vssd1 vccd1 vccd1 _2932_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1814_ _2642_/Q _1802_/X _1813_/X vssd1 vssd1 vccd1 vccd1 _2643_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ _2875_/CLK _2863_/D vssd1 vssd1 vccd1 vccd1 _2863_/Q sky130_fd_sc_hd__dfxtp_1
X_2794_ _2872_/CLK _2794_/D vssd1 vssd1 vccd1 vccd1 _2794_/Q sky130_fd_sc_hd__dfxtp_1
X_1745_ _1748_/B _1746_/B vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__and2b_1
X_1676_ _1673_/Y _2920_/Q _1741_/C _1675_/X vssd1 vssd1 vccd1 vccd1 _1677_/B sky130_fd_sc_hd__a31o_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2228_ _2254_/A vssd1 vssd1 vccd1 vccd1 _2228_/X sky130_fd_sc_hd__clkbuf_1
X_2159_ _2768_/Q _2157_/X _2158_/X vssd1 vssd1 vccd1 vccd1 _2159_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1461_ _2910_/Q _1572_/B vssd1 vssd1 vccd1 vccd1 _1461_/X sky130_fd_sc_hd__and2_1
X_1530_ _2838_/Q _1530_/B input4/X vssd1 vssd1 vccd1 vccd1 _1530_/X sky130_fd_sc_hd__and3b_1
X_1392_ _2797_/Q _1390_/Y _1391_/Y _2796_/Q vssd1 vssd1 vccd1 vccd1 _1392_/X sky130_fd_sc_hd__a22o_1
X_2013_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2915_ _2931_/CLK _2915_/D vssd1 vssd1 vccd1 vccd1 _2915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1728_ _2924_/Q _1380_/B _2925_/Q vssd1 vssd1 vccd1 vccd1 _1731_/B sky130_fd_sc_hd__a21o_1
X_2777_ _2781_/CLK _2777_/D vssd1 vssd1 vccd1 vccd1 _2777_/Q sky130_fd_sc_hd__dfxtp_1
X_2846_ _2866_/CLK _2846_/D vssd1 vssd1 vccd1 vccd1 _2846_/Q sky130_fd_sc_hd__dfxtp_1
X_1659_ _2678_/Q _1697_/A _1659_/C _1659_/D vssd1 vssd1 vccd1 vccd1 _1796_/B sky130_fd_sc_hd__and4_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2700_ _2914_/CLK _2700_/D vssd1 vssd1 vccd1 vccd1 _2700_/Q sky130_fd_sc_hd__dfxtp_1
X_2562_ _2919_/Q _2550_/X _2551_/X vssd1 vssd1 vccd1 vccd1 _2562_/X sky130_fd_sc_hd__o21ba_1
X_2631_ _2947_/Q _1820_/A _1972_/A vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__o21ba_1
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2493_ _2893_/Q _2483_/X _2484_/X vssd1 vssd1 vccd1 vccd1 _2493_/X sky130_fd_sc_hd__o21ba_1
X_1513_ _2844_/Q _1511_/X _1512_/X _2845_/Q vssd1 vssd1 vccd1 vccd1 _1514_/B sky130_fd_sc_hd__a211o_1
X_1444_ input21/X input2/X _1449_/B vssd1 vssd1 vccd1 vccd1 _1444_/X sky130_fd_sc_hd__mux2_1
X_1375_ _1377_/S input8/X vssd1 vssd1 vccd1 vccd1 _1375_/X sky130_fd_sc_hd__and2_1
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2829_ _2839_/CLK _2829_/D vssd1 vssd1 vccd1 vccd1 _2829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _2706_/Q _1985_/X _1992_/X vssd1 vssd1 vccd1 vccd1 _2707_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2545_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2545_/X sky130_fd_sc_hd__clkbuf_2
X_2614_ _2614_/A vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1427_ _2743_/Q vssd1 vssd1 vccd1 vccd1 _1427_/Y sky130_fd_sc_hd__inv_2
X_2476_ _1572_/A _2461_/X _2475_/X vssd1 vssd1 vccd1 vccd1 _2887_/D sky130_fd_sc_hd__o21a_1
X_1358_ input21/X input2/X _2870_/Q vssd1 vssd1 vccd1 vccd1 _1358_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2330_ _1553_/S _2324_/X _2306_/X vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__o21ba_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2261_ _2269_/A _2809_/Q vssd1 vssd1 vccd1 vccd1 _2296_/A sky130_fd_sc_hd__nand2_1
X_2192_ _2780_/Q _2180_/X _2191_/X vssd1 vssd1 vccd1 vccd1 _2781_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_4_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2668_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1976_ _2700_/Q _1967_/X _1975_/X vssd1 vssd1 vccd1 vccd1 _2701_/D sky130_fd_sc_hd__o21a_1
X_2528_ _2909_/Q _2517_/X _2527_/X vssd1 vssd1 vccd1 vccd1 _2906_/D sky130_fd_sc_hd__o21a_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2459_ _2460_/A _2459_/B vssd1 vssd1 vccd1 vccd1 _2880_/D sky130_fd_sc_hd__nor2_1
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1830_ _2649_/Q _1820_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1830_/X sky130_fd_sc_hd__o21ba_1
X_1761_ _1758_/X _1760_/X _1761_/S vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__mux2_1
X_1692_ _1672_/A _1692_/B _2739_/Q vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__and3b_1
X_2313_ _2510_/A vssd1 vssd1 vccd1 vccd1 _2313_/X sky130_fd_sc_hd__clkbuf_2
X_2175_ _2773_/Q _2167_/X _2174_/X vssd1 vssd1 vccd1 vccd1 _2774_/D sky130_fd_sc_hd__o21a_1
X_2244_ _2800_/Q _2240_/X _2241_/X vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1959_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1959_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput38 _1788_/Y vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[7] sky130_fd_sc_hd__clkbuf_1
Xoutput49 _2958_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2931_ _2931_/CLK _2931_/D vssd1 vssd1 vccd1 vccd1 _2931_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_clk repeater2/X vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1813_ _2643_/Q _1805_/X _1808_/X vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__o21ba_1
X_2793_ _2872_/CLK _2793_/D vssd1 vssd1 vccd1 vccd1 _2793_/Q sky130_fd_sc_hd__dfxtp_1
X_2862_ _2875_/CLK _2862_/D vssd1 vssd1 vccd1 vccd1 _2862_/Q sky130_fd_sc_hd__dfxtp_1
X_1744_ _2767_/Q _2768_/Q _2769_/Q _2770_/Q _1748_/B _1746_/B vssd1 vssd1 vccd1 vccd1
+ _1744_/X sky130_fd_sc_hd__mux4_1
X_1675_ _2920_/Q _1514_/X _1674_/Y _2921_/Q vssd1 vssd1 vccd1 vccd1 _1675_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2089_ _2741_/Q _2081_/X _2088_/X vssd1 vssd1 vccd1 vccd1 _2742_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2227_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2227_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2158_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2158_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1460_ _2707_/Q _1456_/X _1458_/Y _2706_/Q _1459_/X vssd1 vssd1 vccd1 vccd1 _1460_/X
+ sky130_fd_sc_hd__a221o_1
X_1391_ _1391_/A _1396_/B vssd1 vssd1 vccd1 vccd1 _1391_/Y sky130_fd_sc_hd__nor2_1
X_2012_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2066_/A sky130_fd_sc_hd__clkbuf_2
X_2914_ _2914_/CLK _2914_/D vssd1 vssd1 vccd1 vccd1 _2914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2845_ _2891_/CLK _2845_/D vssd1 vssd1 vccd1 vccd1 _2845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1658_ _1658_/A _1658_/B _1658_/C vssd1 vssd1 vccd1 vccd1 _1659_/D sky130_fd_sc_hd__or3_1
X_1727_ _1723_/X _1726_/X _1727_/S vssd1 vssd1 vccd1 vccd1 _1727_/X sky130_fd_sc_hd__mux2_1
X_2776_ _2781_/CLK _2776_/D vssd1 vssd1 vccd1 vccd1 _2776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _2648_/Q _1593_/B _1593_/C _1589_/D vssd1 vssd1 vccd1 vccd1 _1589_/X sky130_fd_sc_hd__and4_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2492_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__clkbuf_2
X_2630_ _2660_/Q _2639_/B _2629_/X vssd1 vssd1 vccd1 vccd1 _2946_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2561_ _2611_/A vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__clkbuf_2
X_1512_ _2844_/Q _1512_/B input8/X vssd1 vssd1 vccd1 vccd1 _1512_/X sky130_fd_sc_hd__and3b_1
X_1443_ _2855_/Q vssd1 vssd1 vccd1 vccd1 _1449_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1374_ _2858_/Q vssd1 vssd1 vccd1 vccd1 _1377_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2828_ _2872_/CLK _2828_/D vssd1 vssd1 vccd1 vccd1 _2828_/Q sky130_fd_sc_hd__dfxtp_1
X_2759_ _2765_/CLK _2759_/D vssd1 vssd1 vccd1 vccd1 _2759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_prog_clk clkbuf_2_0_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2875_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1992_ _2707_/Q _1977_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _1992_/X sky130_fd_sc_hd__o21ba_1
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2544_ _2915_/Q _2531_/X _2543_/Y vssd1 vssd1 vccd1 vccd1 _2912_/D sky130_fd_sc_hd__o21a_1
X_2475_ _2887_/Q _2469_/X _2470_/X vssd1 vssd1 vccd1 vccd1 _2475_/X sky130_fd_sc_hd__o21ba_1
X_2613_ _2938_/Q _2611_/X _2612_/Y vssd1 vssd1 vccd1 vccd1 _2939_/D sky130_fd_sc_hd__o21a_1
X_1426_ _2912_/Q vssd1 vssd1 vccd1 vccd1 _1426_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1357_ _2871_/Q _1355_/X _1356_/X vssd1 vssd1 vccd1 vccd1 _1357_/X sky130_fd_sc_hd__a21o_1
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2191_ _2781_/Q _2183_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _2191_/X sky130_fd_sc_hd__o21ba_1
X_2260_ _2805_/Q _2248_/X _2259_/X vssd1 vssd1 vccd1 vccd1 _2806_/D sky130_fd_sc_hd__o21a_1
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1975_ _2701_/Q _1959_/X _1960_/X vssd1 vssd1 vccd1 vccd1 _1975_/X sky130_fd_sc_hd__o21ba_1
X_1409_ _1731_/A vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__buf_2
X_2527_ _2906_/Q _2518_/X _2520_/X vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__o21ba_1
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2458_ _2458_/A vssd1 vssd1 vccd1 vccd1 _2879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2389_ _2857_/Q _2384_/X _2388_/X vssd1 vssd1 vccd1 vccd1 _2852_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1691_ _2738_/Q _1672_/X _1690_/B _1690_/X vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__a31o_1
X_1760_ _2780_/Q _1748_/X _1745_/X _2781_/Q _1759_/X vssd1 vssd1 vccd1 vccd1 _1760_/X
+ sky130_fd_sc_hd__a221o_1
X_2312_ _2824_/Q _2459_/B _2311_/X vssd1 vssd1 vccd1 vccd1 _2825_/D sky130_fd_sc_hd__o21a_1
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2174_ _2774_/Q _2170_/X _2171_/X vssd1 vssd1 vccd1 vccd1 _2174_/X sky130_fd_sc_hd__o21ba_1
X_2243_ _2798_/Q _2235_/X _2242_/X vssd1 vssd1 vccd1 vccd1 _2799_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1958_ _2693_/Q _1954_/X _1957_/X vssd1 vssd1 vccd1 vccd1 _2694_/D sky130_fd_sc_hd__o21a_1
X_1889_ _2667_/Q _1883_/X _1888_/X vssd1 vssd1 vccd1 vccd1 _2668_/D sky130_fd_sc_hd__o21a_1
Xoutput39 _1785_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2930_ _2933_/CLK _2930_/D vssd1 vssd1 vccd1 vccd1 _2930_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2861_ _2875_/CLK _2861_/D vssd1 vssd1 vccd1 vccd1 _2861_/Q sky130_fd_sc_hd__dfxtp_1
X_1812_ _2641_/Q _1802_/X _1811_/X vssd1 vssd1 vccd1 vccd1 _2642_/D sky130_fd_sc_hd__o21a_1
X_1674_ _2920_/Q _1736_/B vssd1 vssd1 vccd1 vccd1 _1674_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2792_ _2937_/CLK _2792_/D vssd1 vssd1 vccd1 vccd1 _2792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1743_ _1743_/A _1747_/C vssd1 vssd1 vccd1 vccd1 _1746_/B sky130_fd_sc_hd__and2_1
X_2226_ _2792_/Q _2222_/X _2225_/X vssd1 vssd1 vccd1 vccd1 _2793_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2088_ _2742_/Q _2082_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__o21ba_1
X_2157_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ _1390_/A _1396_/A vssd1 vssd1 vccd1 vccd1 _1390_/Y sky130_fd_sc_hd__nor2_1
X_2011_ _2712_/Q _1999_/X _2010_/X vssd1 vssd1 vccd1 vccd1 _2713_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2913_ _2914_/CLK _2913_/D vssd1 vssd1 vccd1 vccd1 _2913_/Q sky130_fd_sc_hd__dfxtp_1
X_2844_ _2891_/CLK _2844_/D vssd1 vssd1 vccd1 vccd1 _2844_/Q sky130_fd_sc_hd__dfxtp_1
X_1657_ _1654_/X _1656_/X _1657_/S vssd1 vssd1 vccd1 vccd1 _1658_/C sky130_fd_sc_hd__mux2_1
X_1588_ _1576_/X _1582_/X _1583_/X _1585_/X _1587_/X vssd1 vssd1 vccd1 vccd1 _1588_/X
+ sky130_fd_sc_hd__o32a_1
X_1726_ _2759_/Q _1709_/Y _1724_/X _1725_/X vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__a211o_1
X_2775_ _2781_/CLK _2775_/D vssd1 vssd1 vccd1 vccd1 _2775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2209_ _2948_/Q _2207_/X _2208_/X vssd1 vssd1 vccd1 vccd1 _2787_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2491_ _2560_/A vssd1 vssd1 vccd1 vccd1 _2545_/A sky130_fd_sc_hd__clkbuf_2
X_1511_ input20/X input11/X _2843_/Q vssd1 vssd1 vccd1 vccd1 _1511_/X sky130_fd_sc_hd__mux2_1
X_2560_ _2560_/A vssd1 vssd1 vccd1 vccd1 _2611_/A sky130_fd_sc_hd__clkbuf_2
X_1442_ _2856_/Q vssd1 vssd1 vccd1 vccd1 _1442_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1373_ _2802_/Q _2801_/Q _2800_/Q _2799_/Q _1396_/B _1396_/A vssd1 vssd1 vccd1 vccd1
+ _1373_/X sky130_fd_sc_hd__mux4_1
X_2758_ _2765_/CLK _2758_/D vssd1 vssd1 vccd1 vccd1 _2758_/Q sky130_fd_sc_hd__dfxtp_1
X_2827_ _2949_/CLK _2827_/D vssd1 vssd1 vccd1 vccd1 _2827_/Q sky130_fd_sc_hd__dfxtp_1
X_2689_ _2907_/CLK _2689_/D vssd1 vssd1 vccd1 vccd1 _2689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1709_ _1724_/B _1724_/C vssd1 vssd1 vccd1 vccd1 _1709_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1991_ _2705_/Q _1985_/X _1990_/X vssd1 vssd1 vccd1 vccd1 _2706_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2612_ _1735_/Y _1849_/A _2313_/X vssd1 vssd1 vccd1 vccd1 _2612_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1425_ _2913_/Q vssd1 vssd1 vccd1 vccd1 _1425_/Y sky130_fd_sc_hd__inv_2
X_2543_ _1426_/Y _2542_/X _2510_/X vssd1 vssd1 vccd1 vccd1 _2543_/Y sky130_fd_sc_hd__a21oi_1
X_2474_ _2889_/Q _2461_/X _2473_/X vssd1 vssd1 vccd1 vccd1 _2886_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1356_ _2871_/Q _1356_/B input5/X vssd1 vssd1 vccd1 vccd1 _1356_/X sky130_fd_sc_hd__and3b_1
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2190_ _2779_/Q _2180_/X _2189_/X vssd1 vssd1 vccd1 vccd1 _2780_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ _2699_/Q _1967_/X _1973_/Y vssd1 vssd1 vccd1 vccd1 _2700_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2526_ _2904_/Q _2517_/X _2525_/X vssd1 vssd1 vccd1 vccd1 _2905_/D sky130_fd_sc_hd__o21a_1
X_1408_ _1747_/A vssd1 vssd1 vccd1 vccd1 _1731_/A sky130_fd_sc_hd__buf_2
X_2388_ _1345_/S _2387_/X _2379_/X vssd1 vssd1 vccd1 vccd1 _2388_/X sky130_fd_sc_hd__o21ba_1
X_2457_ _2268_/A _2457_/B vssd1 vssd1 vccd1 vccd1 _2458_/A sky130_fd_sc_hd__and2b_1
XFILLER_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1339_ _2946_/Q _1703_/C vssd1 vssd1 vccd1 vccd1 _1339_/X sky130_fd_sc_hd__and2_1
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2721_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1690_ _1672_/A _1690_/B _2737_/Q vssd1 vssd1 vccd1 vccd1 _1690_/X sky130_fd_sc_hd__and3b_1
X_2311_ _2825_/Q _2301_/X _2306_/X vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__o21ba_1
X_2242_ _2799_/Q _2240_/X _2241_/X vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__o21ba_1
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2173_ _2772_/Q _2167_/X _2172_/X vssd1 vssd1 vccd1 vccd1 _2773_/D sky130_fd_sc_hd__o21a_1
X_1957_ _2694_/Q _1946_/X _1947_/X vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__o21ba_1
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1888_ _2668_/Q _1886_/X _1887_/X vssd1 vssd1 vccd1 vccd1 _1888_/X sky130_fd_sc_hd__o21ba_1
X_2509_ _2898_/Q _2505_/X _2508_/Y vssd1 vssd1 vccd1 vccd1 _2899_/D sky130_fd_sc_hd__o21a_1
Xoutput29 _1795_/Y vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1811_ _2642_/Q _1805_/X _1808_/X vssd1 vssd1 vccd1 vccd1 _1811_/X sky130_fd_sc_hd__o21ba_1
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2791_ _2937_/CLK _2791_/D vssd1 vssd1 vccd1 vccd1 _2791_/Q sky130_fd_sc_hd__dfxtp_1
X_2860_ _2866_/CLK _2860_/D vssd1 vssd1 vccd1 vccd1 _2860_/Q sky130_fd_sc_hd__dfxtp_1
X_1673_ _2921_/Q vssd1 vssd1 vccd1 vccd1 _1673_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1742_ _2937_/Q _1740_/X _1741_/X vssd1 vssd1 vccd1 vccd1 _1747_/C sky130_fd_sc_hd__a21o_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2225_ _2793_/Q _2213_/X _2214_/X vssd1 vssd1 vccd1 vccd1 _2225_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2087_ _2740_/Q _2081_/X _2086_/X vssd1 vssd1 vccd1 vccd1 _2741_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2156_ _2806_/Q _2154_/X _2155_/X vssd1 vssd1 vccd1 vccd1 _2767_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2010_ _2713_/Q _2008_/X _2009_/X vssd1 vssd1 vccd1 vccd1 _2010_/X sky130_fd_sc_hd__o21ba_1
X_2912_ _2923_/CLK _2912_/D vssd1 vssd1 vccd1 vccd1 _2912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1725_ _2758_/Q _1708_/Y _1716_/X _2761_/Q vssd1 vssd1 vccd1 vccd1 _1725_/X sky130_fd_sc_hd__a22o_1
X_2843_ _2858_/CLK _2843_/D vssd1 vssd1 vccd1 vccd1 _2843_/Q sky130_fd_sc_hd__dfxtp_1
X_2774_ _2781_/CLK _2774_/D vssd1 vssd1 vccd1 vccd1 _2774_/Q sky130_fd_sc_hd__dfxtp_1
X_1656_ _2664_/Q _1639_/Y _1641_/Y _2665_/Q _1655_/X vssd1 vssd1 vccd1 vccd1 _1656_/X
+ sky130_fd_sc_hd__a221o_1
X_1587_ _2652_/Q _1578_/X _1597_/C vssd1 vssd1 vccd1 vccd1 _1587_/X sky130_fd_sc_hd__a21o_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _2760_/Q _2137_/X _2138_/X vssd1 vssd1 vccd1 vccd1 _2761_/D sky130_fd_sc_hd__o21a_1
X_2208_ _2787_/Q _2196_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _2208_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1441_ _2914_/Q _1703_/C vssd1 vssd1 vccd1 vccd1 _1441_/X sky130_fd_sc_hd__and2_1
X_2490_ _2895_/Q _2477_/X _2489_/X vssd1 vssd1 vccd1 vccd1 _2892_/D sky130_fd_sc_hd__o21a_1
X_1510_ _1505_/Y _1507_/X _1508_/X _1509_/Y vssd1 vssd1 vccd1 vccd1 _1514_/A sky130_fd_sc_hd__a211o_1
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1372_ _1739_/A _1391_/A vssd1 vssd1 vccd1 vccd1 _1396_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2688_ _2907_/CLK _2688_/D vssd1 vssd1 vccd1 vccd1 _2688_/Q sky130_fd_sc_hd__dfxtp_1
X_1708_ _1716_/B _1716_/C _1747_/A vssd1 vssd1 vccd1 vccd1 _1708_/Y sky130_fd_sc_hd__o21ai_2
X_2757_ _2765_/CLK _2757_/D vssd1 vssd1 vccd1 vccd1 _2757_/Q sky130_fd_sc_hd__dfxtp_1
X_2826_ _2951_/CLK _2826_/D vssd1 vssd1 vccd1 vccd1 _2826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1639_ _1641_/A _1645_/B vssd1 vssd1 vccd1 vccd1 _1639_/Y sky130_fd_sc_hd__nor2_2
XFILLER_58_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1990_ _2706_/Q _1977_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _1990_/X sky130_fd_sc_hd__o21ba_1
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2542_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2542_/X sky130_fd_sc_hd__buf_2
X_2611_ _2611_/A vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1424_ _2722_/Q vssd1 vssd1 vccd1 vccd1 _1424_/Y sky130_fd_sc_hd__inv_2
X_2473_ _1572_/A _2469_/X _2470_/X vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__o21ba_1
X_1355_ input17/X input9/X _1356_/B vssd1 vssd1 vccd1 vccd1 _1355_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2809_ _2951_/CLK _2809_/D vssd1 vssd1 vccd1 vccd1 _2809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ _1867_/A _1861_/X _1972_/X vssd1 vssd1 vccd1 vccd1 _1973_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2525_ _2905_/Q _2518_/X _2520_/X vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__o21ba_1
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1338_ _1334_/X _1335_/X _1336_/X _1337_/X _2877_/Q _2878_/Q vssd1 vssd1 vccd1 vccd1
+ _1703_/C sky130_fd_sc_hd__mux4_2
X_2387_ _2430_/A vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__clkbuf_2
X_1407_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1747_/A sky130_fd_sc_hd__clkbuf_2
X_2456_ _2879_/Q _2808_/Q _2456_/S vssd1 vssd1 vccd1 vccd1 _2457_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2172_ _2773_/Q _2170_/X _2171_/X vssd1 vssd1 vccd1 vccd1 _2172_/X sky130_fd_sc_hd__o21ba_1
X_2241_ _2254_/A vssd1 vssd1 vccd1 vccd1 _2241_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2310_ _2826_/Q _2459_/B _2309_/X vssd1 vssd1 vccd1 vccd1 _2824_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1956_ _2692_/Q _1954_/X _1955_/X vssd1 vssd1 vccd1 vccd1 _2693_/D sky130_fd_sc_hd__o21a_1
X_1887_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1887_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2508_ _1634_/Y _2090_/X _2293_/X vssd1 vssd1 vccd1 vccd1 _2508_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2439_ _2439_/A vssd1 vssd1 vccd1 vccd1 _2439_/X sky130_fd_sc_hd__clkbuf_2
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1810_ _2681_/Q _1802_/X _1809_/X vssd1 vssd1 vccd1 vccd1 _2641_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2790_ _2948_/CLK _2790_/D vssd1 vssd1 vccd1 vccd1 _2790_/Q sky130_fd_sc_hd__dfxtp_1
X_1741_ _2937_/Q _2936_/Q _1741_/C vssd1 vssd1 vccd1 vccd1 _1741_/X sky130_fd_sc_hd__and3b_1
X_1672_ _1672_/A vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2224_ _2791_/Q _2222_/X _2223_/X vssd1 vssd1 vccd1 vccd1 _2792_/D sky130_fd_sc_hd__o21a_1
X_2155_ _2767_/Q _2141_/X _2142_/X vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2086_ _2741_/Q _2082_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1939_ _2686_/Q _1927_/X _1938_/X vssd1 vssd1 vccd1 vccd1 _2687_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2911_ _2914_/CLK _2911_/D vssd1 vssd1 vccd1 vccd1 _2911_/Q sky130_fd_sc_hd__dfxtp_1
X_2842_ _2858_/CLK _2842_/D vssd1 vssd1 vccd1 vccd1 _2842_/Q sky130_fd_sc_hd__dfxtp_1
X_1724_ _2760_/Q _1724_/B _1724_/C vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__and3_1
X_2773_ _2781_/CLK _2773_/D vssd1 vssd1 vccd1 vccd1 _2773_/Q sky130_fd_sc_hd__dfxtp_1
X_1655_ _2663_/Q _1644_/Y _1645_/Y _2662_/Q vssd1 vssd1 vccd1 vccd1 _1655_/X sky130_fd_sc_hd__a22o_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ _2887_/Q _1572_/X _1753_/B _1572_/A _1574_/X vssd1 vssd1 vccd1 vccd1 _1597_/C
+ sky130_fd_sc_hd__o221a_2
X_2069_ _2114_/A vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__clkbuf_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2138_ _2761_/Q _2126_/X _2128_/X vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__o21ba_1
X_2207_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2207_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1440_ _1425_/Y _2912_/Q _1698_/B _1439_/X vssd1 vssd1 vccd1 vccd1 _1457_/B sky130_fd_sc_hd__a31o_1
X_1371_ _1362_/X _1370_/X _2945_/Q vssd1 vssd1 vccd1 vccd1 _1391_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_7_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2907_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2825_ _2933_/CLK _2825_/D vssd1 vssd1 vccd1 vccd1 _2825_/Q sky130_fd_sc_hd__dfxtp_1
X_2687_ _2687_/CLK _2687_/D vssd1 vssd1 vccd1 vccd1 _2687_/Q sky130_fd_sc_hd__dfxtp_1
X_1638_ _1643_/A _1640_/B vssd1 vssd1 vccd1 vccd1 _1645_/B sky130_fd_sc_hd__and2_1
X_2756_ _2765_/CLK _2756_/D vssd1 vssd1 vccd1 vccd1 _2756_/Q sky130_fd_sc_hd__dfxtp_1
X_1707_ _1724_/C _1707_/B vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__and2_1
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1569_ _2891_/Q _1566_/X _1567_/X _1568_/X vssd1 vssd1 vccd1 vccd1 _1589_/D sky130_fd_sc_hd__a31o_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2541_ _2910_/Q _2531_/X _2540_/X vssd1 vssd1 vccd1 vccd1 _2911_/D sky130_fd_sc_hd__o21a_1
X_2472_ _2884_/Q _2461_/X _2471_/X vssd1 vssd1 vccd1 vccd1 _2885_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2610_ _2941_/Q _2600_/X _2609_/X vssd1 vssd1 vccd1 vccd1 _2938_/D sky130_fd_sc_hd__o21a_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1423_ _1421_/X _1422_/X _1778_/A vssd1 vssd1 vccd1 vccd1 _2959_/A sky130_fd_sc_hd__o21a_4
X_1354_ _2870_/Q vssd1 vssd1 vccd1 vccd1 _1356_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2808_ _2951_/CLK _2808_/D vssd1 vssd1 vccd1 vccd1 _2808_/Q sky130_fd_sc_hd__dfxtp_1
X_2739_ _2739_/CLK _2739_/D vssd1 vssd1 vccd1 vccd1 _2739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1972_ _1972_/A vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__clkbuf_4
X_2524_ _2907_/Q _2517_/X _2523_/X vssd1 vssd1 vccd1 vccd1 _2904_/D sky130_fd_sc_hd__o21a_1
X_2455_ _2877_/Q _2460_/B _2454_/X vssd1 vssd1 vccd1 vccd1 _2878_/D sky130_fd_sc_hd__o21a_1
X_1406_ _1643_/A vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__buf_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1337_ _1336_/S _1337_/B vssd1 vssd1 vccd1 vccd1 _1337_/X sky130_fd_sc_hd__and2b_1
X_2386_ _2850_/Q _2384_/X _2385_/X vssd1 vssd1 vccd1 vccd1 _2851_/D sky130_fd_sc_hd__o21a_1
XFILLER_3_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_21_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2781_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2171_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2171_/X sky130_fd_sc_hd__clkbuf_1
X_2240_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2240_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1955_ _2693_/Q _1946_/X _1947_/X vssd1 vssd1 vccd1 vccd1 _1955_/X sky130_fd_sc_hd__o21ba_1
X_1886_ _1899_/A vssd1 vssd1 vccd1 vccd1 _1886_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2507_ _2901_/Q _2505_/X _2506_/X vssd1 vssd1 vccd1 vccd1 _2898_/D sky130_fd_sc_hd__o21a_1
X_2438_ _1356_/B _2425_/X _2437_/X vssd1 vssd1 vccd1 vccd1 _2871_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2369_ _2460_/A _2369_/B vssd1 vssd1 vccd1 vccd1 _2845_/D sky130_fd_sc_hd__nor2_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1671_ _1731_/A _1671_/B _1671_/C vssd1 vssd1 vccd1 vccd1 _1672_/A sky130_fd_sc_hd__and3_1
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1740_ _1514_/X _1784_/D _2936_/Q vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2085_ _2739_/Q _2081_/X _2084_/X vssd1 vssd1 vccd1 vccd1 _2740_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2223_ _2792_/Q _2213_/X _2214_/X vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__o21ba_1
X_2154_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2154_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1938_ _2687_/Q _1932_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _1938_/X sky130_fd_sc_hd__o21ba_1
X_1869_ _2153_/A vssd1 vssd1 vccd1 vccd1 _1927_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2910_ _2923_/CLK _2910_/D vssd1 vssd1 vccd1 vccd1 _2910_/Q sky130_fd_sc_hd__dfxtp_1
X_2841_ _2858_/CLK _2841_/D vssd1 vssd1 vccd1 vccd1 _2841_/Q sky130_fd_sc_hd__dfxtp_1
X_1654_ _2671_/Q _1644_/Y _1645_/Y _2670_/Q _1653_/X vssd1 vssd1 vccd1 vccd1 _1654_/X
+ sky130_fd_sc_hd__a221o_1
X_1723_ _2754_/Q _1708_/Y _1709_/Y _2755_/Q _1722_/X vssd1 vssd1 vccd1 vccd1 _1723_/X
+ sky130_fd_sc_hd__a221o_1
X_2772_ _2815_/CLK _2772_/D vssd1 vssd1 vccd1 vccd1 _2772_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _2649_/Q _1570_/Y _1581_/Y _2651_/Q _1584_/X vssd1 vssd1 vccd1 vccd1 _1585_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2785_/Q _2193_/X _2205_/X vssd1 vssd1 vccd1 vccd1 _2786_/D sky130_fd_sc_hd__o21a_1
X_2068_ _2126_/A vssd1 vssd1 vccd1 vccd1 _2068_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2137_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1370_ _1368_/X _1369_/X _2944_/Q vssd1 vssd1 vccd1 vccd1 _1370_/X sky130_fd_sc_hd__mux2_1
X_2824_ _2951_/CLK _2824_/D vssd1 vssd1 vccd1 vccd1 _2824_/Q sky130_fd_sc_hd__dfxtp_1
X_2686_ _2687_/CLK _2686_/D vssd1 vssd1 vccd1 vccd1 _2686_/Q sky130_fd_sc_hd__dfxtp_1
X_1637_ _1634_/Y _2898_/Q _1703_/C _1636_/X vssd1 vssd1 vccd1 vccd1 _1640_/B sky130_fd_sc_hd__a31o_1
X_2755_ _2755_/CLK _2755_/D vssd1 vssd1 vccd1 vccd1 _2755_/Q sky130_fd_sc_hd__dfxtp_1
X_1706_ _2749_/Q _2748_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1707_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1568_ _2891_/Q _2890_/Q _1703_/C vssd1 vssd1 vccd1 vccd1 _1568_/X sky130_fd_sc_hd__and3b_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1501_/S input1/X vssd1 vssd1 vccd1 vccd1 _1499_/X sky130_fd_sc_hd__and2_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2540_ _2911_/Q _2532_/X _2533_/X vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__o21ba_1
X_2471_ _2885_/Q _2469_/X _2470_/X vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__o21ba_1
XFILLER_9_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1422_ _2765_/Q _2764_/Q _2037_/C vssd1 vssd1 vccd1 vccd1 _1422_/X sky130_fd_sc_hd__and3b_2
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1353_ _1739_/A _1390_/A vssd1 vssd1 vccd1 vccd1 _1396_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2738_ _2931_/CLK _2738_/D vssd1 vssd1 vccd1 vccd1 _2738_/Q sky130_fd_sc_hd__dfxtp_1
X_2807_ _2872_/CLK _2828_/Q vssd1 vssd1 vccd1 vccd1 _2807_/Q sky130_fd_sc_hd__dfxtp_1
X_2669_ _2677_/CLK _2669_/D vssd1 vssd1 vccd1 vccd1 _2669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1971_ _2698_/Q _1967_/X _1970_/Y vssd1 vssd1 vccd1 vccd1 _2699_/D sky130_fd_sc_hd__o21a_1
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1405_ _1457_/A vssd1 vssd1 vccd1 vccd1 _1643_/A sky130_fd_sc_hd__clkbuf_2
X_2523_ _2904_/Q _2518_/X _2520_/X vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__o21ba_1
X_2454_ _2878_/Q _2444_/X _2449_/X vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__o21ba_1
X_2385_ _2851_/Q _2374_/X _2379_/X vssd1 vssd1 vccd1 vccd1 _2385_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1336_ _1385_/B input11/X _1336_/S vssd1 vssd1 vccd1 vccd1 _1336_/X sky130_fd_sc_hd__mux2_1
Xinput1 bi_u1y0n_L1[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0_prog_clk repeater3/X vssd1 vssd1 vccd1 vccd1 clkbuf_0_prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2170_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2170_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1954_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1954_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1885_ _2666_/Q _1883_/X _1884_/X vssd1 vssd1 vccd1 vccd1 _2667_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2506_ _2898_/Q _2499_/X _2500_/X vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__o21ba_1
X_2368_ _1509_/Y _1505_/Y _2400_/S vssd1 vssd1 vccd1 vccd1 _2369_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2437_ _2871_/Q _2430_/X _2436_/X vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__o21ba_1
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _2840_/Q vssd1 vssd1 vccd1 vccd1 _1322_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_2299_ _2820_/Q _2285_/X _2290_/X vssd1 vssd1 vccd1 vccd1 _2299_/X sky130_fd_sc_hd__o21ba_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1670_ _2922_/Q _1438_/B _1669_/Y _1793_/C vssd1 vssd1 vccd1 vccd1 _1671_/C sky130_fd_sc_hd__o22a_1
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2222_ _2477_/A vssd1 vssd1 vccd1 vccd1 _2222_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2084_ _2740_/Q _2082_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _2084_/X sky130_fd_sc_hd__o21ba_1
XFILLER_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2153_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2207_/A sky130_fd_sc_hd__clkbuf_2
X_1937_ _2685_/Q _1927_/X _1936_/X vssd1 vssd1 vccd1 vccd1 _2686_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1868_ _1868_/A vssd1 vssd1 vccd1 vccd1 _2153_/A sky130_fd_sc_hd__buf_4
X_1799_ _2464_/A _2883_/Q vssd1 vssd1 vccd1 vccd1 _1868_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2840_ _2858_/CLK _2840_/D vssd1 vssd1 vccd1 vccd1 _2840_/Q sky130_fd_sc_hd__dfxtp_1
X_2771_ _2815_/CLK _2771_/D vssd1 vssd1 vccd1 vccd1 _2771_/Q sky130_fd_sc_hd__dfxtp_1
X_1653_ _2672_/Q _1639_/Y _1641_/Y _2673_/Q vssd1 vssd1 vccd1 vccd1 _1653_/X sky130_fd_sc_hd__a22o_1
X_1584_ _2650_/Q _1593_/B _1584_/C _1589_/D vssd1 vssd1 vccd1 vccd1 _1584_/X sky130_fd_sc_hd__and4_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _2757_/Q _1716_/X _1721_/X vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__a21o_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2786_/Q _2196_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__o21ba_1
X_2067_ _2212_/A vssd1 vssd1 vccd1 vccd1 _2126_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2136_ _2759_/Q _2123_/X _2135_/X vssd1 vssd1 vccd1 vccd1 _2760_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2754_ _2755_/CLK _2754_/D vssd1 vssd1 vccd1 vccd1 _2754_/Q sky130_fd_sc_hd__dfxtp_1
X_1705_ _1743_/A _1716_/B vssd1 vssd1 vccd1 vccd1 _1724_/B sky130_fd_sc_hd__nand2_2
X_2823_ _2951_/CLK _2823_/D vssd1 vssd1 vccd1 vccd1 _2823_/Q sky130_fd_sc_hd__dfxtp_1
X_2685_ _2687_/CLK _2685_/D vssd1 vssd1 vccd1 vccd1 _2685_/Q sky130_fd_sc_hd__dfxtp_1
X_1636_ _2898_/Q _1765_/C _1635_/Y _2899_/Q vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__o211a_1
X_1567_ _2958_/A _2890_/Q vssd1 vssd1 vccd1 vccd1 _1567_/X sky130_fd_sc_hd__or2b_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2119_ _2754_/Q _2113_/X _2114_/X vssd1 vssd1 vccd1 vccd1 _2119_/X sky130_fd_sc_hd__o21ba_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _2861_/Q vssd1 vssd1 vccd1 vccd1 _1501_/S sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_15_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2755_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2470_ _2500_/A vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__clkbuf_1
X_1421_ _2764_/Q _2724_/Q _2765_/Q vssd1 vssd1 vccd1 vccd1 _1421_/X sky130_fd_sc_hd__and3b_1
X_1352_ _1339_/X _1351_/X _2947_/Q vssd1 vssd1 vccd1 vccd1 _1390_/A sky130_fd_sc_hd__mux2_2
X_2668_ _2668_/CLK _2668_/D vssd1 vssd1 vccd1 vccd1 _2668_/Q sky130_fd_sc_hd__dfxtp_1
X_2737_ _2739_/CLK _2737_/D vssd1 vssd1 vccd1 vccd1 _2737_/Q sky130_fd_sc_hd__dfxtp_1
X_2806_ _2937_/CLK _2806_/D vssd1 vssd1 vccd1 vccd1 _2806_/Q sky130_fd_sc_hd__dfxtp_1
X_1619_ _2892_/Q _1467_/B _1618_/Y _2893_/Q vssd1 vssd1 vccd1 vccd1 _1619_/X sky130_fd_sc_hd__o211a_1
X_2599_ _2932_/Q _2587_/X _2598_/X vssd1 vssd1 vccd1 vccd1 _2933_/D sky130_fd_sc_hd__o21a_1
XFILLER_75_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1970_ _1867_/B _1861_/X _2639_/A vssd1 vssd1 vccd1 vccd1 _1970_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2522_ _2902_/Q _2517_/X _2521_/X vssd1 vssd1 vccd1 vccd1 _2903_/D sky130_fd_sc_hd__o21a_1
X_2453_ _1336_/S _2460_/B _2452_/X vssd1 vssd1 vccd1 vccd1 _2877_/D sky130_fd_sc_hd__o21a_1
X_1404_ _2806_/Q _2805_/Q _2151_/C vssd1 vssd1 vccd1 vccd1 _1404_/X sky130_fd_sc_hd__and3b_2
X_2384_ _2384_/A vssd1 vssd1 vccd1 vccd1 _2384_/X sky130_fd_sc_hd__clkbuf_2
X_1335_ input13/X input7/X _2876_/Q vssd1 vssd1 vccd1 vccd1 _1335_/X sky130_fd_sc_hd__mux2_1
Xinput2 bi_u1y0n_L1[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_prog_clk clkbuf_2_0_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2858_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1953_ _2691_/Q _1941_/X _1952_/X vssd1 vssd1 vccd1 vccd1 _2692_/D sky130_fd_sc_hd__o21a_1
X_1884_ _2667_/Q _1873_/X _1874_/X vssd1 vssd1 vccd1 vccd1 _1884_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2505_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2367_ _1512_/B _2352_/X _2366_/Y vssd1 vssd1 vccd1 vccd1 _2844_/D sky130_fd_sc_hd__o21a_1
X_2298_ _2818_/Q _2296_/X _2297_/X vssd1 vssd1 vccd1 vccd1 _2819_/D sky130_fd_sc_hd__o21a_1
X_1318_ _2942_/Q _1572_/B vssd1 vssd1 vccd1 vccd1 _1318_/X sky130_fd_sc_hd__and2_1
X_2436_ _2500_/A vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__clkbuf_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2221_ _2560_/A vssd1 vssd1 vccd1 vccd1 _2477_/A sky130_fd_sc_hd__clkbuf_2
X_2152_ _2152_/A vssd1 vssd1 vccd1 vccd1 _2766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2083_ _2114_/A vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1936_ _2686_/Q _1932_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__o21ba_1
X_1867_ _1867_/A _1867_/B _2269_/A _1867_/D vssd1 vssd1 vccd1 vccd1 _2661_/D sky130_fd_sc_hd__nor4_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1798_ _2322_/A vssd1 vssd1 vccd1 vccd1 _2464_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2419_ _2869_/Q _2412_/X _2418_/X vssd1 vssd1 vccd1 vccd1 _2864_/D sky130_fd_sc_hd__o21a_1
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1721_ _2756_/Q _1724_/B _1724_/C vssd1 vssd1 vccd1 vccd1 _1721_/X sky130_fd_sc_hd__and3_1
X_2770_ _2815_/CLK _2770_/D vssd1 vssd1 vccd1 vccd1 _2770_/Q sky130_fd_sc_hd__dfxtp_1
X_1652_ _1658_/A _1658_/B _1647_/X _1651_/X vssd1 vssd1 vccd1 vccd1 _1659_/C sky130_fd_sc_hd__a2bb2o_1
X_1583_ _2654_/Q _1583_/B _1584_/C _1593_/D vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__and4_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _2760_/Q _2126_/X _2128_/X vssd1 vssd1 vccd1 vccd1 _2135_/X sky130_fd_sc_hd__o21ba_1
X_2204_ _2784_/Q _2193_/X _2203_/Y vssd1 vssd1 vccd1 vccd1 _2785_/D sky130_fd_sc_hd__o21a_1
X_2066_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2066_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1919_ _2679_/Q _1915_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__o21ba_1
X_2899_ _2947_/CLK _2899_/D vssd1 vssd1 vccd1 vccd1 _2899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2684_ _2687_/CLK _2684_/D vssd1 vssd1 vccd1 vccd1 _2684_/Q sky130_fd_sc_hd__dfxtp_1
X_2753_ _2755_/CLK _2753_/D vssd1 vssd1 vccd1 vccd1 _2753_/Q sky130_fd_sc_hd__dfxtp_1
X_1704_ _2931_/Q _1702_/X _1703_/X vssd1 vssd1 vccd1 vccd1 _1716_/B sky130_fd_sc_hd__a21o_1
X_2822_ _2822_/CLK _2822_/D vssd1 vssd1 vccd1 vccd1 _2822_/Q sky130_fd_sc_hd__dfxtp_1
X_1497_ _1495_/X _1496_/X _2907_/Q vssd1 vssd1 vccd1 vccd1 _1520_/B sky130_fd_sc_hd__mux2_1
X_1635_ _2898_/Q _1736_/B vssd1 vssd1 vccd1 vccd1 _1635_/Y sky130_fd_sc_hd__nand2_1
X_1566_ _1451_/A _1451_/B _2890_/Q vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__a21o_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ _2727_/Q _2039_/X _2048_/X vssd1 vssd1 vccd1 vccd1 _2728_/D sky130_fd_sc_hd__o21a_1
X_2118_ _2752_/Q _2110_/X _2117_/X vssd1 vssd1 vccd1 vccd1 _2753_/D sky130_fd_sc_hd__o21a_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1351_ _1765_/C _1793_/C _2946_/Q vssd1 vssd1 vccd1 vccd1 _1351_/X sky130_fd_sc_hd__mux2_1
X_1420_ _1420_/A _1736_/B vssd1 vssd1 vccd1 vccd1 _2961_/A sky130_fd_sc_hd__nor2_4
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2805_ _2937_/CLK _2805_/D vssd1 vssd1 vccd1 vccd1 _2805_/Q sky130_fd_sc_hd__dfxtp_2
X_2667_ _2668_/CLK _2667_/D vssd1 vssd1 vccd1 vccd1 _2667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2736_ _2739_/CLK _2736_/D vssd1 vssd1 vccd1 vccd1 _2736_/Q sky130_fd_sc_hd__dfxtp_1
X_1618_ _2892_/Q _1762_/A vssd1 vssd1 vccd1 vccd1 _1618_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1549_ _1337_/B input2/X _2831_/Q vssd1 vssd1 vccd1 vccd1 _1549_/X sky130_fd_sc_hd__mux2_1
X_2598_ _2933_/Q _2596_/X _2597_/X vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__o21ba_1
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2521_ _2903_/Q _2518_/X _2520_/X vssd1 vssd1 vccd1 vccd1 _2521_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2452_ _2877_/Q _2444_/X _2449_/X vssd1 vssd1 vccd1 vccd1 _2452_/X sky130_fd_sc_hd__o21ba_1
X_2383_ _1435_/S _2370_/X _2382_/X vssd1 vssd1 vccd1 vccd1 _2850_/D sky130_fd_sc_hd__o21a_1
X_1403_ _1395_/X _1402_/X _2803_/Q vssd1 vssd1 vccd1 vccd1 _2151_/C sky130_fd_sc_hd__o21a_1
X_1334_ _1336_/S input1/X vssd1 vssd1 vccd1 vccd1 _1334_/X sky130_fd_sc_hd__and2_1
Xinput3 bi_u1y0n_L1[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2719_ _2721_/CLK _2719_/D vssd1 vssd1 vccd1 vccd1 _2719_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_0_prog_clk clkbuf_2_0_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2891_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1952_ _2692_/Q _1946_/X _1947_/X vssd1 vssd1 vccd1 vccd1 _1952_/X sky130_fd_sc_hd__o21ba_1
X_1883_ _1927_/A vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__clkbuf_2
X_2504_ _2896_/Q _2492_/X _2503_/X vssd1 vssd1 vccd1 vccd1 _2897_/D sky130_fd_sc_hd__o21a_1
X_2435_ _2519_/A vssd1 vssd1 vccd1 vccd1 _2500_/A sky130_fd_sc_hd__clkbuf_2
X_2366_ _1505_/Y _2460_/B _2293_/X vssd1 vssd1 vccd1 vccd1 _2366_/Y sky130_fd_sc_hd__a21oi_1
X_2297_ _2819_/Q _2285_/X _2290_/X vssd1 vssd1 vccd1 vccd1 _2297_/X sky130_fd_sc_hd__o21ba_1
X_1317_ _1313_/X _1314_/X _1315_/X _1316_/X _2865_/Q _2866_/Q vssd1 vssd1 vccd1 vccd1
+ _1572_/B sky130_fd_sc_hd__mux4_2
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2082_ _2126_/A vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2220_ _2790_/Q _2207_/X _2219_/X vssd1 vssd1 vccd1 vccd1 _2791_/D sky130_fd_sc_hd__o21a_1
X_2151_ _2804_/Q _2151_/B _2151_/C vssd1 vssd1 vccd1 vccd1 _2152_/A sky130_fd_sc_hd__and3_1
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1935_ _2684_/Q _1927_/X _1934_/X vssd1 vssd1 vccd1 vccd1 _2685_/D sky130_fd_sc_hd__o21a_1
X_1797_ _1797_/A vssd1 vssd1 vccd1 vccd1 _2640_/D sky130_fd_sc_hd__clkbuf_1
X_1866_ _2700_/Q vssd1 vssd1 vccd1 vccd1 _1867_/A sky130_fd_sc_hd__inv_2
X_2418_ _1315_/S _2417_/X _2409_/X vssd1 vssd1 vccd1 vccd1 _2418_/X sky130_fd_sc_hd__o21ba_1
X_2349_ _1530_/B _2339_/X _2348_/X vssd1 vssd1 vccd1 vccd1 _2838_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1651_ _1651_/A _1651_/B _1651_/C vssd1 vssd1 vccd1 vccd1 _1651_/X sky130_fd_sc_hd__or3_1
X_1720_ _1707_/X _1715_/X _1719_/X vssd1 vssd1 vccd1 vccd1 _1720_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1582_ _2656_/Q _1578_/X _1581_/Y _2655_/Q vssd1 vssd1 vccd1 vccd1 _1582_/X sky130_fd_sc_hd__a22o_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2065_ _2733_/Q _2052_/X _2064_/X vssd1 vssd1 vccd1 vccd1 _2734_/D sky130_fd_sc_hd__o21a_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _2758_/Q _2123_/X _2133_/X vssd1 vssd1 vccd1 vccd1 _2759_/D sky130_fd_sc_hd__o21a_1
X_2203_ _1417_/Y _2090_/X _1972_/X vssd1 vssd1 vccd1 vccd1 _2203_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1918_ _2677_/Q _1910_/X _1917_/X vssd1 vssd1 vccd1 vccd1 _2678_/D sky130_fd_sc_hd__o21a_1
X_1849_ _1849_/A vssd1 vssd1 vccd1 vccd1 _1849_/X sky130_fd_sc_hd__clkbuf_2
X_2898_ _2947_/CLK _2898_/D vssd1 vssd1 vccd1 vccd1 _2898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2821_ _2822_/CLK _2821_/D vssd1 vssd1 vccd1 vccd1 _2821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2683_ _2907_/CLK _2683_/D vssd1 vssd1 vccd1 vccd1 _2683_/Q sky130_fd_sc_hd__dfxtp_1
X_2752_ _2755_/CLK _2752_/D vssd1 vssd1 vccd1 vccd1 _2752_/Q sky130_fd_sc_hd__dfxtp_1
X_1634_ _2899_/Q vssd1 vssd1 vccd1 vccd1 _1634_/Y sky130_fd_sc_hd__inv_2
X_1703_ _2931_/Q _2930_/Q _1703_/C vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__and3b_1
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1496_ _1368_/X _2959_/A _2906_/Q vssd1 vssd1 vccd1 vccd1 _1496_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1565_ _2889_/Q _1562_/X _1563_/Y _1564_/X _1698_/B vssd1 vssd1 vccd1 vccd1 _1593_/C
+ sky130_fd_sc_hd__a32o_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2048_ _2728_/Q _2040_/X _2041_/X vssd1 vssd1 vccd1 vccd1 _2048_/X sky130_fd_sc_hd__o21ba_1
X_2117_ _2753_/Q _2113_/X _2114_/X vssd1 vssd1 vccd1 vccd1 _2117_/X sky130_fd_sc_hd__o21ba_1
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1350_ _2958_/A vssd1 vssd1 vccd1 vccd1 _1793_/C sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_24_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2951_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2804_ _2937_/CLK _2804_/D vssd1 vssd1 vccd1 vccd1 _2804_/Q sky130_fd_sc_hd__dfxtp_1
X_2666_ _2668_/CLK _2666_/D vssd1 vssd1 vccd1 vccd1 _2666_/Q sky130_fd_sc_hd__dfxtp_1
X_2735_ _2735_/CLK _2735_/D vssd1 vssd1 vccd1 vccd1 _2735_/Q sky130_fd_sc_hd__dfxtp_1
X_1617_ _1617_/A _1617_/B vssd1 vssd1 vccd1 vccd1 _1762_/A sky130_fd_sc_hd__nor2_2
X_2597_ _2615_/A vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1479_ _1469_/Y _1478_/X _1468_/X vssd1 vssd1 vccd1 vccd1 _1479_/X sky130_fd_sc_hd__o21ba_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1548_ _2832_/Q vssd1 vssd1 vccd1 vccd1 _1548_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2520_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__clkbuf_1
X_1402_ _1328_/A _1398_/X _1401_/X vssd1 vssd1 vccd1 vccd1 _1402_/X sky130_fd_sc_hd__o21a_1
X_2451_ _2879_/Q _2439_/X _2450_/X vssd1 vssd1 vccd1 vccd1 _2876_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2382_ _2850_/Q _2374_/X _2379_/X vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__o21ba_1
Xinput4 bi_u1y0n_L1[1] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
X_1333_ _2876_/Q vssd1 vssd1 vccd1 vccd1 _1336_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2718_ _2735_/CLK _2718_/D vssd1 vssd1 vccd1 vccd1 _2718_/Q sky130_fd_sc_hd__dfxtp_1
X_2649_ _2839_/CLK _2649_/D vssd1 vssd1 vccd1 vccd1 _2649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1951_ _2690_/Q _1941_/X _1950_/X vssd1 vssd1 vccd1 vccd1 _2691_/D sky130_fd_sc_hd__o21a_1
X_1882_ _2665_/Q _1870_/X _1881_/X vssd1 vssd1 vccd1 vccd1 _2666_/D sky130_fd_sc_hd__o21a_1
X_2503_ _2897_/Q _2499_/X _2500_/X vssd1 vssd1 vccd1 vccd1 _2503_/X sky130_fd_sc_hd__o21ba_1
X_2365_ _2439_/A vssd1 vssd1 vccd1 vccd1 _2460_/B sky130_fd_sc_hd__clkbuf_2
X_2434_ _2875_/Q _2425_/X _2433_/X vssd1 vssd1 vccd1 vccd1 _2870_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1316_ _1315_/S _1533_/B vssd1 vssd1 vccd1 vccd1 _1316_/X sky130_fd_sc_hd__and2b_1
X_2296_ _2296_/A vssd1 vssd1 vccd1 vccd1 _2296_/X sky130_fd_sc_hd__clkbuf_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2081_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__clkbuf_2
X_2150_ _2764_/Q _2137_/X _2149_/X vssd1 vssd1 vccd1 vccd1 _2765_/D sky130_fd_sc_hd__o21a_1
X_1934_ _2685_/Q _1932_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__o21ba_1
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1796_ _2679_/Q _1796_/B vssd1 vssd1 vccd1 vccd1 _1797_/A sky130_fd_sc_hd__and2_1
X_1865_ _2659_/Q _1849_/X _1864_/Y vssd1 vssd1 vccd1 vccd1 _2660_/D sky130_fd_sc_hd__o21a_1
X_2348_ _2838_/Q _2340_/X _2345_/X vssd1 vssd1 vccd1 vccd1 _2348_/X sky130_fd_sc_hd__o21ba_1
X_2417_ _2430_/A vssd1 vssd1 vccd1 vccd1 _2417_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2279_ _2815_/Q _2262_/X _2278_/X vssd1 vssd1 vccd1 vccd1 _2812_/D sky130_fd_sc_hd__o21a_1
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1650_ _2667_/Q _1644_/Y _1645_/Y _2666_/Q vssd1 vssd1 vccd1 vccd1 _1651_/C sky130_fd_sc_hd__a22o_1
X_1581_ _1581_/A _1584_/C _1593_/D vssd1 vssd1 vccd1 vccd1 _1581_/Y sky130_fd_sc_hd__nor3_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2783_/Q _2193_/X _2201_/X vssd1 vssd1 vccd1 vccd1 _2784_/D sky130_fd_sc_hd__o21a_1
X_2064_ _2734_/Q _2053_/X _2055_/X vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__o21ba_1
X_2133_ _2759_/Q _2126_/X _2128_/X vssd1 vssd1 vccd1 vccd1 _2133_/X sky130_fd_sc_hd__o21ba_1
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1917_ _2678_/Q _1915_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__o21ba_1
X_2897_ _2947_/CLK _2897_/D vssd1 vssd1 vccd1 vccd1 _2897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1848_ _2654_/Q _1834_/X _1847_/X vssd1 vssd1 vccd1 vccd1 _2655_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1779_ _1779_/A vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2751_ _2755_/CLK _2751_/D vssd1 vssd1 vccd1 vccd1 _2751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2820_ _2822_/CLK _2820_/D vssd1 vssd1 vccd1 vccd1 _2820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1633_ _1739_/A _1643_/B vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__nand2_1
X_2682_ _2950_/CLK _2682_/D vssd1 vssd1 vccd1 vccd1 _2682_/Q sky130_fd_sc_hd__dfxtp_1
X_1702_ _1451_/X _1793_/C _2930_/Q vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__mux2_1
X_1564_ _2889_/Q _2888_/Q vssd1 vssd1 vccd1 vccd1 _1564_/X sky130_fd_sc_hd__and2b_1
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1495_ _2906_/Q _1741_/C vssd1 vssd1 vccd1 vccd1 _1495_/X sky130_fd_sc_hd__and2_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ _2726_/Q _2039_/X _2046_/X vssd1 vssd1 vccd1 vccd1 _2727_/D sky130_fd_sc_hd__o21a_1
X_2116_ _2751_/Q _2110_/X _2115_/X vssd1 vssd1 vccd1 vccd1 _2752_/D sky130_fd_sc_hd__o21a_1
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2949_ _2949_/CLK _2949_/D vssd1 vssd1 vccd1 vccd1 _2949_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2734_ _2735_/CLK _2734_/D vssd1 vssd1 vccd1 vccd1 _2734_/Q sky130_fd_sc_hd__dfxtp_1
X_2803_ _2937_/CLK _2803_/D vssd1 vssd1 vccd1 vccd1 _2803_/Q sky130_fd_sc_hd__dfxtp_1
X_2665_ _2668_/CLK _2665_/D vssd1 vssd1 vccd1 vccd1 _2665_/Q sky130_fd_sc_hd__dfxtp_1
X_1547_ _2900_/Q vssd1 vssd1 vccd1 vccd1 _1547_/Y sky130_fd_sc_hd__inv_2
X_1616_ _2893_/Q vssd1 vssd1 vccd1 vccd1 _1616_/Y sky130_fd_sc_hd__inv_2
X_2596_ _2614_/A vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__clkbuf_2
X_1478_ _2719_/Q _1456_/X _1458_/Y _2718_/Q _1477_/X vssd1 vssd1 vccd1 vccd1 _1478_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2381_ _2854_/Q _2370_/X _2380_/X vssd1 vssd1 vccd1 vccd1 _2849_/D sky130_fd_sc_hd__o21a_1
X_1401_ _1328_/Y _1400_/X _1388_/X vssd1 vssd1 vccd1 vccd1 _1401_/X sky130_fd_sc_hd__o21ba_1
X_2450_ _1336_/S _2444_/X _2449_/X vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__o21ba_1
X_1332_ _1457_/A vssd1 vssd1 vccd1 vccd1 _1739_/A sky130_fd_sc_hd__buf_4
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput5 bi_u1y0n_L1[2] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2717_ _2735_/CLK _2717_/D vssd1 vssd1 vccd1 vccd1 _2717_/Q sky130_fd_sc_hd__dfxtp_1
X_2648_ _2839_/CLK _2648_/D vssd1 vssd1 vccd1 vccd1 _2648_/Q sky130_fd_sc_hd__dfxtp_1
X_2579_ _2926_/Q _2570_/X _2571_/X vssd1 vssd1 vccd1 vccd1 _2579_/X sky130_fd_sc_hd__o21ba_1
XFILLER_10_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1950_ _2691_/Q _1946_/X _1947_/X vssd1 vssd1 vccd1 vccd1 _1950_/X sky130_fd_sc_hd__o21ba_1
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1881_ _2666_/Q _1873_/X _1874_/X vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__o21ba_1
X_2502_ _2899_/Q _2492_/X _2501_/X vssd1 vssd1 vccd1 vccd1 _2896_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1315_ _1385_/B input12/X _1315_/S vssd1 vssd1 vccd1 vccd1 _1315_/X sky130_fd_sc_hd__mux2_1
X_2433_ _1356_/B _2430_/X _2422_/X vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__o21ba_1
X_2364_ _2364_/A vssd1 vssd1 vccd1 vccd1 _2439_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2295_ _2821_/Q _2282_/X _2294_/Y vssd1 vssd1 vccd1 vccd1 _2818_/D sky130_fd_sc_hd__o21a_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2080_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2137_/A sky130_fd_sc_hd__clkbuf_2
X_1933_ _1960_/A vssd1 vssd1 vccd1 vccd1 _1933_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1864_ _1600_/A _1861_/X _2639_/A vssd1 vssd1 vccd1 vccd1 _1864_/Y sky130_fd_sc_hd__a21oi_1
X_1795_ _1793_/Y _1794_/X _1420_/A vssd1 vssd1 vccd1 vccd1 _1795_/Y sky130_fd_sc_hd__a21oi_2
X_2347_ _2842_/Q _2339_/X _2346_/X vssd1 vssd1 vccd1 vccd1 _2837_/D sky130_fd_sc_hd__o21a_1
X_2416_ _2862_/Q _2412_/X _2415_/X vssd1 vssd1 vccd1 vccd1 _2863_/D sky130_fd_sc_hd__o21a_1
X_2278_ _2812_/Q _2264_/X _2277_/X vssd1 vssd1 vccd1 vccd1 _2278_/X sky130_fd_sc_hd__o21ba_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_18_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2822_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1580_ _1589_/D vssd1 vssd1 vccd1 vccd1 _1593_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _2757_/Q _2123_/X _2131_/X vssd1 vssd1 vccd1 vccd1 _2758_/D sky130_fd_sc_hd__o21a_1
X_2201_ _2784_/Q _2196_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _2201_/X sky130_fd_sc_hd__o21ba_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2063_ _2732_/Q _2052_/X _2062_/X vssd1 vssd1 vccd1 vccd1 _2733_/D sky130_fd_sc_hd__o21a_1
X_1916_ _1960_/A vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__clkbuf_1
X_1847_ _2655_/Q _1837_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _1847_/X sky130_fd_sc_hd__o21ba_1
X_2896_ _2947_/CLK _2896_/D vssd1 vssd1 vccd1 vccd1 _2896_/Q sky130_fd_sc_hd__dfxtp_1
X_1778_ _1778_/A _1778_/B _1778_/C vssd1 vssd1 vccd1 vccd1 _1779_/A sky130_fd_sc_hd__and3_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2681_ _2687_/CLK _2681_/D vssd1 vssd1 vccd1 vccd1 _2681_/Q sky130_fd_sc_hd__dfxtp_1
X_2750_ _2755_/CLK _2750_/D vssd1 vssd1 vccd1 vccd1 _2750_/Q sky130_fd_sc_hd__dfxtp_1
X_1701_ _1743_/A _1716_/C vssd1 vssd1 vccd1 vccd1 _1724_/C sky130_fd_sc_hd__and2_1
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1632_ _1630_/X _1631_/X _2897_/Q vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__mux2_1
X_1563_ _1581_/A _1736_/B _2888_/Q vssd1 vssd1 vccd1 vccd1 _1563_/Y sky130_fd_sc_hd__o21ai_2
X_1494_ _1490_/X _1491_/X _1492_/X _1493_/X _2868_/Q _2869_/Q vssd1 vssd1 vccd1 vccd1
+ _1741_/C sky130_fd_sc_hd__mux4_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2115_ _2752_/Q _2113_/X _2114_/X vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__o21ba_1
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2046_ _2727_/Q _2040_/X _2041_/X vssd1 vssd1 vccd1 vccd1 _2046_/X sky130_fd_sc_hd__o21ba_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2948_ _2948_/CLK _2948_/D vssd1 vssd1 vccd1 vccd1 _2948_/Q sky130_fd_sc_hd__dfxtp_1
X_2879_ _2949_/CLK _2879_/D vssd1 vssd1 vccd1 vccd1 _2879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2733_ _2735_/CLK _2733_/D vssd1 vssd1 vccd1 vccd1 _2733_/Q sky130_fd_sc_hd__dfxtp_1
X_2664_ _2668_/CLK _2664_/D vssd1 vssd1 vccd1 vccd1 _2664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2802_ _2949_/CLK _2802_/D vssd1 vssd1 vccd1 vccd1 _2802_/Q sky130_fd_sc_hd__dfxtp_1
X_1477_ _2717_/Q _1455_/Y _1471_/Y _2716_/Q vssd1 vssd1 vccd1 vccd1 _1477_/X sky130_fd_sc_hd__a22o_1
X_1546_ _1539_/S _1542_/Y _1545_/Y vssd1 vssd1 vccd1 vccd1 _1546_/X sky130_fd_sc_hd__a21o_1
X_1615_ _2895_/Q _2894_/Q _1754_/C vssd1 vssd1 vccd1 vccd1 _1658_/B sky130_fd_sc_hd__and3b_1
X_2595_ _2935_/Q _2587_/X _2594_/X vssd1 vssd1 vccd1 vccd1 _2932_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2029_ _2720_/Q _2022_/X _2023_/X vssd1 vssd1 vccd1 vccd1 _2029_/X sky130_fd_sc_hd__o21ba_1
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1331_ _1598_/B vssd1 vssd1 vccd1 vccd1 _1457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1400_ _2793_/Q _1390_/Y _1391_/Y _2792_/Q _1399_/X vssd1 vssd1 vccd1 vccd1 _1400_/X
+ sky130_fd_sc_hd__a221o_1
X_2380_ _1435_/S _2374_/X _2379_/X vssd1 vssd1 vccd1 vccd1 _2380_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput6 bi_u1y0n_L1[3] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_2716_ _2735_/CLK _2716_/D vssd1 vssd1 vccd1 vccd1 _2716_/Q sky130_fd_sc_hd__dfxtp_1
X_2647_ _2839_/CLK _2647_/D vssd1 vssd1 vccd1 vccd1 _2647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1529_ input16/X input9/X _1530_/B vssd1 vssd1 vccd1 vccd1 _1529_/X sky130_fd_sc_hd__mux2_1
X_2578_ _2924_/Q _2574_/X _2577_/X vssd1 vssd1 vccd1 vccd1 _2925_/D sky130_fd_sc_hd__o21a_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1880_ _2664_/Q _1870_/X _1879_/X vssd1 vssd1 vccd1 vccd1 _2665_/D sky130_fd_sc_hd__o21a_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2501_ _2896_/Q _2499_/X _2500_/X vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__o21ba_1
X_2294_ _1783_/Y _2459_/B _2293_/X vssd1 vssd1 vccd1 vccd1 _2294_/Y sky130_fd_sc_hd__a21oi_1
X_2363_ _2848_/Q _2352_/X _2362_/X vssd1 vssd1 vccd1 vccd1 _2843_/D sky130_fd_sc_hd__o21a_1
X_2432_ _2868_/Q _2425_/X _2431_/X vssd1 vssd1 vccd1 vccd1 _2869_/D sky130_fd_sc_hd__o21a_1
X_1314_ input16/X input7/X _2864_/Q vssd1 vssd1 vccd1 vccd1 _1314_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1932_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1932_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1863_ _1972_/A vssd1 vssd1 vccd1 vccd1 _2639_/A sky130_fd_sc_hd__buf_2
Xinput20 bi_u1y0s_L1[5] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
X_1794_ _2824_/Q _1794_/B _2825_/Q vssd1 vssd1 vccd1 vccd1 _1794_/X sky130_fd_sc_hd__or3b_1
X_2415_ _2863_/Q _2404_/X _2409_/X vssd1 vssd1 vccd1 vccd1 _2415_/X sky130_fd_sc_hd__o21ba_1
X_2346_ _1530_/B _2340_/X _2345_/X vssd1 vssd1 vccd1 vccd1 _2346_/X sky130_fd_sc_hd__o21ba_1
X_2277_ _2345_/A vssd1 vssd1 vccd1 vccd1 _2277_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2062_ _2733_/Q _2053_/X _2055_/X vssd1 vssd1 vccd1 vccd1 _2062_/X sky130_fd_sc_hd__o21ba_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _2758_/Q _2126_/X _2128_/X vssd1 vssd1 vccd1 vccd1 _2131_/X sky130_fd_sc_hd__o21ba_1
X_2200_ _2782_/Q _2193_/X _2199_/X vssd1 vssd1 vccd1 vccd1 _2783_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1915_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1915_/X sky130_fd_sc_hd__clkbuf_2
X_1846_ _2653_/Q _1834_/X _1845_/X vssd1 vssd1 vccd1 vccd1 _2654_/D sky130_fd_sc_hd__o21a_1
X_2895_ _2947_/CLK _2895_/D vssd1 vssd1 vccd1 vccd1 _2895_/Q sky130_fd_sc_hd__dfxtp_1
X_1777_ _2814_/Q _1369_/X _2815_/Q vssd1 vssd1 vccd1 vccd1 _1778_/C sky130_fd_sc_hd__a21o_1
XFILLER_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2329_ _2329_/A vssd1 vssd1 vccd1 vccd1 _2830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2680_ _2687_/CLK _2680_/D vssd1 vssd1 vccd1 vccd1 _2680_/Q sky130_fd_sc_hd__dfxtp_2
X_1631_ _1368_/X _2955_/A _2896_/Q vssd1 vssd1 vccd1 vccd1 _1631_/X sky130_fd_sc_hd__mux2_1
X_1700_ _1698_/X _1699_/X _2929_/Q vssd1 vssd1 vccd1 vccd1 _1716_/C sky130_fd_sc_hd__mux2_1
X_1562_ _1514_/A _1514_/B _2888_/Q vssd1 vssd1 vccd1 vccd1 _1562_/X sky130_fd_sc_hd__a21o_1
X_1493_ _1492_/S _1533_/B vssd1 vssd1 vccd1 vccd1 _1493_/X sky130_fd_sc_hd__and2b_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2045_ _2725_/Q _2039_/X _2044_/X vssd1 vssd1 vccd1 vccd1 _2726_/D sky130_fd_sc_hd__o21a_1
X_2114_ _2114_/A vssd1 vssd1 vccd1 vccd1 _2114_/X sky130_fd_sc_hd__clkbuf_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2947_ _2947_/CLK _2947_/D vssd1 vssd1 vccd1 vccd1 _2947_/Q sky130_fd_sc_hd__dfxtp_1
X_1829_ _2647_/Q _1819_/X _1828_/X vssd1 vssd1 vccd1 vccd1 _2648_/D sky130_fd_sc_hd__o21a_1
X_2878_ _2891_/CLK _2878_/D vssd1 vssd1 vccd1 vccd1 _2878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_3_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2839_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2801_ _2949_/CLK _2801_/D vssd1 vssd1 vccd1 vccd1 _2801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2732_ _2735_/CLK _2732_/D vssd1 vssd1 vccd1 vccd1 _2732_/Q sky130_fd_sc_hd__dfxtp_1
X_2663_ _2668_/CLK _2663_/D vssd1 vssd1 vccd1 vccd1 _2663_/Q sky130_fd_sc_hd__dfxtp_1
X_1614_ _1487_/Y _2954_/A _1613_/X _2895_/Q vssd1 vssd1 vccd1 vccd1 _1658_/A sky130_fd_sc_hd__o211a_1
X_2594_ _2932_/Q _2583_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__o21ba_1
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1476_ _1476_/A _1476_/B _1476_/C vssd1 vssd1 vccd1 vccd1 _1476_/X sky130_fd_sc_hd__or3_1
X_1545_ _2695_/Q _1521_/X _1544_/X vssd1 vssd1 vccd1 vccd1 _1545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2028_ _2718_/Q _2026_/X _2027_/X vssd1 vssd1 vccd1 vccd1 _2719_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1330_ _1583_/B vssd1 vssd1 vccd1 vccd1 _1598_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput7 bi_u1y0n_L1[4] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2715_ _2735_/CLK _2715_/D vssd1 vssd1 vccd1 vccd1 _2715_/Q sky130_fd_sc_hd__dfxtp_1
X_2646_ _2839_/CLK _2646_/D vssd1 vssd1 vccd1 vccd1 _2646_/Q sky130_fd_sc_hd__dfxtp_1
X_2577_ _2925_/Q _2570_/X _2571_/X vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__o21ba_1
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1459_ _2704_/Q _1459_/B _1459_/C vssd1 vssd1 vccd1 vccd1 _1459_/X sky130_fd_sc_hd__and3_1
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1528_ _2837_/Q vssd1 vssd1 vccd1 vccd1 _1530_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2500_ _2500_/A vssd1 vssd1 vccd1 vccd1 _2500_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2431_ _2869_/Q _2430_/X _2422_/X vssd1 vssd1 vccd1 vccd1 _2431_/X sky130_fd_sc_hd__o21ba_1
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2293_ _2510_/A vssd1 vssd1 vccd1 vccd1 _2293_/X sky130_fd_sc_hd__buf_2
X_2362_ _1512_/B _2353_/X _2359_/X vssd1 vssd1 vccd1 vccd1 _2362_/X sky130_fd_sc_hd__o21ba_1
X_1313_ _1315_/S input4/X vssd1 vssd1 vccd1 vccd1 _1313_/X sky130_fd_sc_hd__and2_1
XFILLER_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2629_ _2946_/Q _1820_/A _1972_/A vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__o21ba_1
XFILLER_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_45 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1931_ _2683_/Q _1927_/X _1930_/X vssd1 vssd1 vccd1 vccd1 _2684_/D sky130_fd_sc_hd__o21a_1
Xinput10 bi_u1y0n_L1[7] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_2
Xinput21 bi_u1y0s_L1[6] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
X_1862_ _2615_/A vssd1 vssd1 vccd1 vccd1 _1972_/A sky130_fd_sc_hd__clkbuf_1
X_1793_ _2825_/Q _2824_/Q _1793_/C vssd1 vssd1 vccd1 vccd1 _1793_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2414_ _1501_/S _2412_/X _2413_/X vssd1 vssd1 vccd1 vccd1 _2862_/D sky130_fd_sc_hd__o21a_1
X_2345_ _2345_/A vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2276_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2345_/A sky130_fd_sc_hd__buf_2
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clkbuf_2_0_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2872_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2061_ _2731_/Q _2052_/X _2060_/X vssd1 vssd1 vccd1 vccd1 _2732_/D sky130_fd_sc_hd__o21a_1
X_2130_ _2756_/Q _2123_/X _2129_/X vssd1 vssd1 vccd1 vccd1 _2757_/D sky130_fd_sc_hd__o21a_1
X_1914_ _2212_/A vssd1 vssd1 vccd1 vccd1 _1977_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1845_ _2654_/Q _1837_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _1845_/X sky130_fd_sc_hd__o21ba_1
X_2894_ _2947_/CLK _2894_/D vssd1 vssd1 vccd1 vccd1 _2894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1776_ _2814_/Q _1786_/A _2815_/Q vssd1 vssd1 vccd1 vccd1 _1778_/B sky130_fd_sc_hd__o21ai_1
X_2328_ _2313_/X _2456_/S vssd1 vssd1 vccd1 vccd1 _2329_/A sky130_fd_sc_hd__and2b_1
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2259_ _2806_/Q _2253_/X _2254_/X vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1630_ _2896_/Q _1630_/B vssd1 vssd1 vccd1 vccd1 _1630_/X sky130_fd_sc_hd__and2_1
X_1561_ _1597_/B vssd1 vssd1 vccd1 vccd1 _1561_/Y sky130_fd_sc_hd__inv_2
X_1492_ input20/X input12/X _1492_/S vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__mux2_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2044_ _2726_/Q _2040_/X _2041_/X vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__o21ba_1
X_2113_ _2126_/A vssd1 vssd1 vccd1 vccd1 _2113_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2946_ _2946_/CLK _2946_/D vssd1 vssd1 vccd1 vccd1 _2946_/Q sky130_fd_sc_hd__dfxtp_1
X_2877_ _2891_/CLK _2877_/D vssd1 vssd1 vccd1 vccd1 _2877_/Q sky130_fd_sc_hd__dfxtp_1
X_1828_ _2648_/Q _1820_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1828_/X sky130_fd_sc_hd__o21ba_1
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1759_ _2782_/Q _1747_/X _1746_/Y _2779_/Q vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2731_ _2735_/CLK _2731_/D vssd1 vssd1 vccd1 vccd1 _2731_/Q sky130_fd_sc_hd__dfxtp_1
X_2800_ _2872_/CLK _2800_/D vssd1 vssd1 vccd1 vccd1 _2800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1544_ _2696_/Q _1518_/X _1543_/X _1539_/S vssd1 vssd1 vccd1 vccd1 _1544_/X sky130_fd_sc_hd__a211o_1
X_2662_ _2677_/CLK _2662_/D vssd1 vssd1 vccd1 vccd1 _2662_/Q sky130_fd_sc_hd__dfxtp_1
X_1613_ _2894_/Q _1613_/B vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__or2_1
X_2593_ _2930_/Q _2587_/X _2592_/X vssd1 vssd1 vccd1 vccd1 _2931_/D sky130_fd_sc_hd__o21a_1
X_1475_ _2713_/Q _1455_/Y _1458_/Y _2714_/Q vssd1 vssd1 vccd1 vccd1 _1476_/C sky130_fd_sc_hd__a22o_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2027_ _2719_/Q _2022_/X _2023_/X vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__o21ba_1
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2929_ _2933_/CLK _2929_/D vssd1 vssd1 vccd1 vccd1 _2929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput8 bi_u1y0n_L1[5] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2714_ _2735_/CLK _2714_/D vssd1 vssd1 vccd1 vccd1 _2714_/Q sky130_fd_sc_hd__dfxtp_1
X_1527_ _2902_/Q _1380_/B _2903_/Q vssd1 vssd1 vccd1 vccd1 _1538_/A sky130_fd_sc_hd__a21o_1
X_2645_ _2893_/CLK _2645_/D vssd1 vssd1 vccd1 vccd1 _2645_/Q sky130_fd_sc_hd__dfxtp_1
X_2576_ _2927_/Q _2574_/X _2575_/X vssd1 vssd1 vccd1 vccd1 _2924_/D sky130_fd_sc_hd__o21a_1
X_1458_ _1458_/A _1459_/C vssd1 vssd1 vccd1 vccd1 _1458_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1389_ _1396_/A _1396_/B vssd1 vssd1 vccd1 vccd1 _1389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2361_ _2841_/Q _2352_/X _2360_/X vssd1 vssd1 vccd1 vccd1 _2842_/D sky130_fd_sc_hd__o21a_1
X_2430_ _2430_/A vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2292_ _2816_/Q _2282_/X _2291_/X vssd1 vssd1 vccd1 vccd1 _2817_/D sky130_fd_sc_hd__o21a_1
X_1312_ _2864_/Q vssd1 vssd1 vccd1 vccd1 _1315_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_2559_ _2639_/A _2559_/B vssd1 vssd1 vccd1 vccd1 _2918_/D sky130_fd_sc_hd__nor2_1
X_2628_ _2944_/Q _2639_/B _2627_/X vssd1 vssd1 vccd1 vccd1 _2945_/D sky130_fd_sc_hd__o21a_1
XFILLER_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1930_ _2684_/Q _1915_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__o21ba_1
X_1861_ _2624_/A vssd1 vssd1 vccd1 vccd1 _1861_/X sky130_fd_sc_hd__clkbuf_2
Xinput11 bi_u1y0n_L1[8] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
Xinput22 bi_u1y0s_L1[7] vssd1 vssd1 vccd1 vccd1 _1502_/B sky130_fd_sc_hd__buf_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1792_ _1792_/A vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2344_ _2835_/Q _2339_/X _2343_/X vssd1 vssd1 vccd1 vccd1 _2836_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _2766_/CLK sky130_fd_sc_hd__clkbuf_16
X_2413_ _2862_/Q _2404_/X _2409_/X vssd1 vssd1 vccd1 vccd1 _2413_/X sky130_fd_sc_hd__o21ba_1
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2275_ _2810_/Q _2262_/X _2274_/X vssd1 vssd1 vccd1 vccd1 _2811_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2060_ _2732_/Q _2053_/X _2055_/X vssd1 vssd1 vccd1 vccd1 _2060_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1913_ _2482_/A vssd1 vssd1 vccd1 vccd1 _2212_/A sky130_fd_sc_hd__buf_4
X_2893_ _2893_/CLK _2893_/D vssd1 vssd1 vccd1 vccd1 _2893_/Q sky130_fd_sc_hd__dfxtp_1
X_1844_ _2652_/Q _1834_/X _1843_/X vssd1 vssd1 vccd1 vccd1 _2653_/D sky130_fd_sc_hd__o21a_1
Xrepeater1 repeater1/A vssd1 vssd1 vccd1 vccd1 _2950_/CLK sky130_fd_sc_hd__buf_2
X_1775_ _1773_/X _1774_/X _1420_/A vssd1 vssd1 vccd1 vccd1 _1775_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2258_ _2804_/Q _2248_/X _2257_/X vssd1 vssd1 vccd1 vccd1 _2805_/D sky130_fd_sc_hd__o21a_1
X_2327_ _2464_/A _2880_/Q vssd1 vssd1 vccd1 vccd1 _2456_/S sky130_fd_sc_hd__and2_1
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2189_ _2780_/Q _2183_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _2189_/X sky130_fd_sc_hd__o21ba_1
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1560_ _2884_/Q _1764_/B _1558_/X _1559_/X vssd1 vssd1 vccd1 vccd1 _1597_/B sky130_fd_sc_hd__o211a_2
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2112_ _2750_/Q _2110_/X _2111_/X vssd1 vssd1 vccd1 vccd1 _2751_/D sky130_fd_sc_hd__o21a_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1491_ input16/X input8/X _2867_/Q vssd1 vssd1 vccd1 vccd1 _1491_/X sky130_fd_sc_hd__mux2_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2043_ _2765_/Q _2039_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _2725_/D sky130_fd_sc_hd__o21a_1
X_1827_ _2646_/Q _1819_/X _1826_/X vssd1 vssd1 vccd1 vccd1 _2647_/D sky130_fd_sc_hd__o21a_1
X_2945_ _2947_/CLK _2945_/D vssd1 vssd1 vccd1 vccd1 _2945_/Q sky130_fd_sc_hd__dfxtp_1
X_2876_ _2943_/CLK _2876_/D vssd1 vssd1 vccd1 vccd1 _2876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1689_ _1689_/A vssd1 vssd1 vccd1 vccd1 _1690_/B sky130_fd_sc_hd__inv_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1758_ _2776_/Q _1748_/X _1745_/X _2777_/Q _1757_/X vssd1 vssd1 vccd1 vccd1 _1758_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2661_ _2950_/CLK _2661_/D vssd1 vssd1 vccd1 vccd1 _2661_/Q sky130_fd_sc_hd__dfxtp_1
X_2730_ _2735_/CLK _2730_/D vssd1 vssd1 vccd1 vccd1 _2730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1474_ _2715_/Q _1456_/X _1471_/Y _2712_/Q vssd1 vssd1 vccd1 vccd1 _1476_/B sky130_fd_sc_hd__a22o_1
X_1543_ _2698_/Q _1522_/Y _1519_/Y _2697_/Q vssd1 vssd1 vccd1 vccd1 _1543_/X sky130_fd_sc_hd__a22o_1
X_2592_ _2931_/Q _2583_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _2592_/X sky130_fd_sc_hd__o21ba_1
X_1612_ _1612_/A vssd1 vssd1 vccd1 vccd1 _2954_/A sky130_fd_sc_hd__buf_4
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_11_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2881_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2026_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2026_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2928_ _2931_/CLK _2928_/D vssd1 vssd1 vccd1 vccd1 _2928_/Q sky130_fd_sc_hd__dfxtp_1
X_2859_ _2866_/CLK _2859_/D vssd1 vssd1 vccd1 vccd1 _2859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput9 bi_u1y0n_L1[6] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2713_ _2735_/CLK _2713_/D vssd1 vssd1 vccd1 vccd1 _2713_/Q sky130_fd_sc_hd__dfxtp_1
X_2644_ _2893_/CLK _2644_/D vssd1 vssd1 vccd1 vccd1 _2644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1526_ _2684_/Q _1518_/X _1519_/Y _2685_/Q _1525_/X vssd1 vssd1 vccd1 vccd1 _1526_/X
+ sky130_fd_sc_hd__a221o_1
X_1457_ _1457_/A _1457_/B vssd1 vssd1 vccd1 vccd1 _1459_/C sky130_fd_sc_hd__nand2_1
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2575_ _2924_/Q _2570_/X _2571_/X vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__o21ba_1
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1388_ _1380_/X _1387_/X _2941_/Q vssd1 vssd1 vccd1 vccd1 _1388_/X sky130_fd_sc_hd__mux2_1
X_2009_ _2041_/A vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2360_ _2842_/Q _2353_/X _2359_/X vssd1 vssd1 vccd1 vccd1 _2360_/X sky130_fd_sc_hd__o21ba_1
X_2291_ _2817_/Q _2285_/X _2290_/X vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__o21ba_1
X_1311_ _2805_/Q _2766_/Q _2806_/Q vssd1 vssd1 vccd1 vccd1 _1311_/X sky130_fd_sc_hd__and3b_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2627_ _2945_/Q _1820_/A _1972_/A vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2558_ _1673_/Y _1681_/Y _2624_/A vssd1 vssd1 vccd1 vccd1 _2559_/B sky130_fd_sc_hd__mux2_1
X_2489_ _2892_/Q _2483_/X _2484_/X vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__o21ba_1
X_1509_ _2845_/Q vssd1 vssd1 vccd1 vccd1 _1509_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ _2560_/A vssd1 vssd1 vccd1 vccd1 _2624_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput12 bi_u1y0n_L1[9] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
Xinput23 bi_u1y0s_L1[8] vssd1 vssd1 vccd1 vccd1 _1337_/B sky130_fd_sc_hd__clkbuf_2
X_1791_ _2037_/B _1791_/B _1791_/C vssd1 vssd1 vccd1 vccd1 _1792_/A sky130_fd_sc_hd__and3_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2343_ _2836_/Q _2340_/X _2332_/X vssd1 vssd1 vccd1 vccd1 _2343_/X sky130_fd_sc_hd__o21ba_1
X_2412_ _2439_/A vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__clkbuf_2
X_2274_ _2811_/Q _2264_/X _2254_/X vssd1 vssd1 vccd1 vccd1 _2274_/X sky130_fd_sc_hd__o21ba_1
XFILLER_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1989_ _2704_/Q _1985_/X _1988_/X vssd1 vssd1 vccd1 vccd1 _2705_/D sky130_fd_sc_hd__o21a_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2961_ _2961_/A vssd1 vssd1 vccd1 vccd1 _2961_/X sky130_fd_sc_hd__clkbuf_1
X_1912_ _2676_/Q _1910_/X _1911_/X vssd1 vssd1 vccd1 vccd1 _2677_/D sky130_fd_sc_hd__o21a_1
X_1843_ _2653_/Q _1837_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _1843_/X sky130_fd_sc_hd__o21ba_1
X_2892_ _2893_/CLK _2892_/D vssd1 vssd1 vccd1 vccd1 _2892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1774_ _2812_/Q _1794_/B _2813_/Q vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__or3b_1
Xrepeater2 clk vssd1 vssd1 vccd1 vccd1 repeater2/X sky130_fd_sc_hd__buf_2
X_2326_ _2833_/Q _2321_/X _2325_/X vssd1 vssd1 vccd1 vccd1 _2829_/D sky130_fd_sc_hd__o21a_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2257_ _2805_/Q _2253_/X _2254_/X vssd1 vssd1 vccd1 vccd1 _2257_/X sky130_fd_sc_hd__o21ba_1
XFILLER_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2188_ _2778_/Q _2180_/X _2187_/X vssd1 vssd1 vccd1 vccd1 _2779_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1490_ _1492_/S input4/X vssd1 vssd1 vccd1 vccd1 _1490_/X sky130_fd_sc_hd__and2_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2042_ _2725_/Q _2040_/X _2041_/X vssd1 vssd1 vccd1 vccd1 _2042_/X sky130_fd_sc_hd__o21ba_1
X_2111_ _2751_/Q _2100_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _2111_/X sky130_fd_sc_hd__o21ba_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1826_ _2647_/Q _1820_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1826_/X sky130_fd_sc_hd__o21ba_1
X_2944_ _2947_/CLK _2944_/D vssd1 vssd1 vccd1 vccd1 _2944_/Q sky130_fd_sc_hd__dfxtp_1
X_2875_ _2875_/CLK _2875_/D vssd1 vssd1 vccd1 vccd1 _2875_/Q sky130_fd_sc_hd__dfxtp_2
X_1688_ _1662_/Y _1663_/X _1765_/C _1666_/X vssd1 vssd1 vccd1 vccd1 _1688_/Y sky130_fd_sc_hd__a31oi_1
X_1757_ _2778_/Q _1747_/X _1746_/Y _2775_/Q vssd1 vssd1 vccd1 vccd1 _1757_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2309_ _2824_/Q _2301_/X _2306_/X vssd1 vssd1 vccd1 vccd1 _2309_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2660_ _2946_/CLK _2660_/D vssd1 vssd1 vccd1 vccd1 _2660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1611_ _1747_/A _1611_/B vssd1 vssd1 vccd1 vccd1 _1612_/A sky130_fd_sc_hd__and2_1
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1542_ _2692_/Q _1518_/X _1519_/Y _2693_/Q _1541_/X vssd1 vssd1 vccd1 vccd1 _1542_/Y
+ sky130_fd_sc_hd__a221oi_1
X_1473_ _2711_/Q _1456_/X _1470_/X _1472_/X vssd1 vssd1 vccd1 vccd1 _1473_/X sky130_fd_sc_hd__a211o_1
X_2591_ _2933_/Q _2587_/X _2590_/X vssd1 vssd1 vccd1 vccd1 _2930_/D sky130_fd_sc_hd__o21a_1
X_2025_ _2717_/Q _2013_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _2718_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2927_ _2933_/CLK _2927_/D vssd1 vssd1 vccd1 vccd1 _2927_/Q sky130_fd_sc_hd__dfxtp_1
X_1809_ _2641_/Q _1805_/X _1808_/X vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__o21ba_1
X_2789_ _2937_/CLK _2789_/D vssd1 vssd1 vccd1 vccd1 _2789_/Q sky130_fd_sc_hd__dfxtp_1
X_2858_ _2858_/CLK _2858_/D vssd1 vssd1 vccd1 vccd1 _2858_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2712_ _2735_/CLK _2712_/D vssd1 vssd1 vccd1 vccd1 _2712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2643_ _2947_/CLK _2643_/D vssd1 vssd1 vccd1 vccd1 _2643_/Q sky130_fd_sc_hd__dfxtp_1
X_2574_ _2611_/A vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__clkbuf_2
X_1456_ _1643_/A _1457_/B _1458_/A vssd1 vssd1 vccd1 vccd1 _1456_/X sky130_fd_sc_hd__and3_1
X_1525_ _2683_/Q _1521_/X _1522_/Y _2686_/Q vssd1 vssd1 vccd1 vccd1 _1525_/X sky130_fd_sc_hd__a22o_1
X_1387_ _1467_/B _1661_/X _2940_/Q vssd1 vssd1 vccd1 vccd1 _1387_/X sky130_fd_sc_hd__mux2_1
X_2008_ _2053_/A vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2290_ _2345_/A vssd1 vssd1 vccd1 vccd1 _2290_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2557_ _1663_/X _2545_/X _2556_/Y vssd1 vssd1 vccd1 vccd1 _2917_/D sky130_fd_sc_hd__o21a_1
X_2626_ _2947_/Q _2639_/B _2625_/X vssd1 vssd1 vccd1 vccd1 _2944_/D sky130_fd_sc_hd__o21a_1
X_1439_ _1426_/Y _2960_/A _1438_/X _2913_/Q vssd1 vssd1 vccd1 vccd1 _1439_/X sky130_fd_sc_hd__o211a_1
X_2488_ _2890_/Q _2477_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _2891_/D sky130_fd_sc_hd__o21a_1
X_1508_ _1512_/B _1624_/B _2844_/Q vssd1 vssd1 vccd1 vccd1 _1508_/X sky130_fd_sc_hd__and3b_1
XFILLER_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 bi_u1y0s_L1[0] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1790_ _2822_/Q _1369_/X _2823_/Q vssd1 vssd1 vccd1 vccd1 _1791_/C sky130_fd_sc_hd__a21o_1
Xinput24 bi_u1y0s_L1[9] vssd1 vssd1 vccd1 vccd1 _1533_/B sky130_fd_sc_hd__buf_2
X_2411_ _2866_/Q _2397_/X _2410_/X vssd1 vssd1 vccd1 vccd1 _2861_/D sky130_fd_sc_hd__o21a_1
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2342_ _1384_/S _2339_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _2835_/D sky130_fd_sc_hd__o21a_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2273_ _2813_/Q _2262_/X _2272_/Y vssd1 vssd1 vccd1 vccd1 _2810_/D sky130_fd_sc_hd__o21a_1
XFILLER_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1988_ _2705_/Q _1977_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__o21ba_1
XFILLER_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xclkbuf_leaf_6_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2687_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2609_ _2938_/Q _2596_/X _2597_/X vssd1 vssd1 vccd1 vccd1 _2609_/X sky130_fd_sc_hd__o21ba_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2960_ _2960_/A vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1911_ _2677_/Q _1899_/X _1901_/X vssd1 vssd1 vccd1 vccd1 _1911_/X sky130_fd_sc_hd__o21ba_1
X_1842_ _2651_/Q _1834_/X _1841_/X vssd1 vssd1 vccd1 vccd1 _2652_/D sky130_fd_sc_hd__o21a_1
X_2891_ _2891_/CLK _2891_/D vssd1 vssd1 vccd1 vccd1 _2891_/Q sky130_fd_sc_hd__dfxtp_1
X_1773_ _1786_/A _2813_/Q _2812_/Q vssd1 vssd1 vccd1 vccd1 _1773_/X sky130_fd_sc_hd__or3b_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xrepeater3 prog_clk vssd1 vssd1 vccd1 vccd1 repeater3/X sky130_fd_sc_hd__buf_2
X_2325_ _2829_/Q _2324_/X _2306_/X vssd1 vssd1 vccd1 vccd1 _2325_/X sky130_fd_sc_hd__o21ba_1
X_2187_ _2779_/Q _2183_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _2187_/X sky130_fd_sc_hd__o21ba_1
X_2256_ _2803_/Q _2248_/X _2255_/X vssd1 vssd1 vccd1 vccd1 _2804_/D sky130_fd_sc_hd__o21a_1
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2041_ _2041_/A vssd1 vssd1 vccd1 vccd1 _2041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2110_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2110_/X sky130_fd_sc_hd__clkbuf_2
X_2943_ _2943_/CLK _2943_/D vssd1 vssd1 vccd1 vccd1 _2943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1825_ _2645_/Q _1819_/X _1824_/X vssd1 vssd1 vccd1 vccd1 _2646_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1756_ _1744_/X _1750_/X _1761_/S vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__mux2_1
X_2874_ _2949_/CLK _2874_/D vssd1 vssd1 vccd1 vccd1 _2874_/Q sky130_fd_sc_hd__dfxtp_1
X_1687_ _2733_/Q _2734_/Q _2735_/Q _2736_/Q _1672_/X _1692_/B vssd1 vssd1 vccd1 vccd1
+ _1687_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2308_ _2822_/Q _2296_/X _2307_/X vssd1 vssd1 vccd1 vccd1 _2823_/D sky130_fd_sc_hd__o21a_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2239_ _2797_/Q _2235_/X _2238_/X vssd1 vssd1 vccd1 vccd1 _2798_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1610_ _1867_/B _1867_/D _1608_/X _1609_/Y vssd1 vssd1 vccd1 vccd1 _1611_/B sky130_fd_sc_hd__o31ai_4
X_2590_ _2930_/Q _2583_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__o21ba_1
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1472_ _2710_/Q _1458_/Y _1471_/Y _2708_/Q vssd1 vssd1 vccd1 vccd1 _1472_/X sky130_fd_sc_hd__a22o_1
X_1541_ _2691_/Q _1521_/X _1522_/Y _2694_/Q vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2024_ _2718_/Q _2022_/X _2023_/X vssd1 vssd1 vccd1 vccd1 _2024_/X sky130_fd_sc_hd__o21ba_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2926_ _2933_/CLK _2926_/D vssd1 vssd1 vccd1 vccd1 _2926_/Q sky130_fd_sc_hd__dfxtp_1
X_2857_ _2891_/CLK _2857_/D vssd1 vssd1 vccd1 vccd1 _2857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xclkbuf_leaf_20_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2815_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1808_ _2510_/A vssd1 vssd1 vccd1 vccd1 _1808_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2788_ _2937_/CLK _2788_/D vssd1 vssd1 vccd1 vccd1 _2788_/Q sky130_fd_sc_hd__dfxtp_1
X_1739_ _1739_/A _1747_/B vssd1 vssd1 vccd1 vccd1 _1748_/B sky130_fd_sc_hd__and2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2711_ _2721_/CLK _2711_/D vssd1 vssd1 vccd1 vccd1 _2711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1524_ _2688_/Q _1518_/X _1519_/Y _2689_/Q _1523_/X vssd1 vssd1 vccd1 vccd1 _1524_/X
+ sky130_fd_sc_hd__a221o_1
X_2642_ _2893_/CLK _2642_/D vssd1 vssd1 vccd1 vccd1 _2642_/Q sky130_fd_sc_hd__dfxtp_1
X_2573_ _2922_/Q _2561_/X _2572_/X vssd1 vssd1 vccd1 vccd1 _2923_/D sky130_fd_sc_hd__o21a_1
X_1455_ _1457_/B _1459_/B vssd1 vssd1 vccd1 vccd1 _1455_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1386_ _1382_/X _1383_/X _1384_/X _1385_/X _2835_/Q _2836_/Q vssd1 vssd1 vccd1 vccd1
+ _1467_/B sky130_fd_sc_hd__mux4_2
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2007_ _2711_/Q _1999_/X _2006_/X vssd1 vssd1 vccd1 vccd1 _2712_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2909_ _2923_/CLK _2909_/D vssd1 vssd1 vccd1 vccd1 _2909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2556_ _1662_/Y _2542_/X _2510_/X vssd1 vssd1 vccd1 vccd1 _2556_/Y sky130_fd_sc_hd__a21oi_1
X_2487_ _2891_/Q _2483_/X _2484_/X vssd1 vssd1 vccd1 vccd1 _2487_/X sky130_fd_sc_hd__o21ba_1
X_1507_ _1337_/B input3/X _1512_/B vssd1 vssd1 vccd1 vccd1 _1507_/X sky130_fd_sc_hd__mux2_1
X_2625_ _2944_/Q _2614_/X _2615_/X vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__o21ba_1
X_1438_ _2912_/Q _1438_/B vssd1 vssd1 vccd1 vccd1 _1438_/X sky130_fd_sc_hd__or2_1
XFILLER_46_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1369_ _2959_/A vssd1 vssd1 vccd1 vccd1 _1369_/X sky130_fd_sc_hd__buf_2
XFILLER_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput14 bi_u1y0s_L1[10] vssd1 vssd1 vccd1 vccd1 _1551_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput25 prog_din vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2341_ _2835_/Q _2340_/X _2332_/X vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__o21ba_1
X_2410_ _1501_/S _2404_/X _2409_/X vssd1 vssd1 vccd1 vccd1 _2410_/X sky130_fd_sc_hd__o21ba_1
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2272_ _1770_/Y _2459_/B _1972_/X vssd1 vssd1 vccd1 vccd1 _2272_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1987_ _2744_/Q _1985_/X _1986_/X vssd1 vssd1 vccd1 vccd1 _2704_/D sky130_fd_sc_hd__o21a_1
XFILLER_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2539_ _2913_/Q _2531_/X _2538_/X vssd1 vssd1 vccd1 vccd1 _2910_/D sky130_fd_sc_hd__o21a_1
X_2608_ _2936_/Q _2600_/X _2607_/X vssd1 vssd1 vccd1 vccd1 _2937_/D sky130_fd_sc_hd__o21a_1
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1910_ _1927_/A vssd1 vssd1 vccd1 vccd1 _1910_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2890_ _2947_/CLK _2890_/D vssd1 vssd1 vccd1 vccd1 _2890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1841_ _2652_/Q _1837_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _1841_/X sky130_fd_sc_hd__o21ba_1
X_1772_ _2811_/Q _1770_/Y _2954_/A _1771_/X vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__a31o_2
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2324_ _2400_/S vssd1 vssd1 vccd1 vccd1 _2324_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2186_ _2777_/Q _2180_/X _2185_/X vssd1 vssd1 vccd1 vccd1 _2778_/D sky130_fd_sc_hd__o21a_1
X_2255_ _2804_/Q _2253_/X _2254_/X vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__o21ba_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2040_ _2053_/A vssd1 vssd1 vccd1 vccd1 _2040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2942_ _2943_/CLK _2942_/D vssd1 vssd1 vccd1 vccd1 _2942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2873_ _2891_/CLK _2873_/D vssd1 vssd1 vccd1 vccd1 _2873_/Q sky130_fd_sc_hd__dfxtp_1
X_1824_ _2646_/Q _1820_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1824_/X sky130_fd_sc_hd__o21ba_1
X_1686_ _1679_/X _1680_/X _1686_/S vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__mux2_1
X_1755_ _2935_/Q _1752_/X _1753_/X _1754_/X vssd1 vssd1 vccd1 vccd1 _1761_/S sky130_fd_sc_hd__a31o_1
X_2238_ _2798_/Q _2227_/X _2228_/X vssd1 vssd1 vccd1 vccd1 _2238_/X sky130_fd_sc_hd__o21ba_1
X_2307_ _2823_/Q _2301_/X _2306_/X vssd1 vssd1 vccd1 vccd1 _2307_/X sky130_fd_sc_hd__o21ba_1
XFILLER_72_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2169_ _2771_/Q _2167_/X _2168_/X vssd1 vssd1 vccd1 vccd1 _2772_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1540_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1540_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1471_ _1643_/A _1458_/A _1457_/B vssd1 vssd1 vccd1 vccd1 _1471_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2023_ _2041_/A vssd1 vssd1 vccd1 vccd1 _2023_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2856_ _2891_/CLK _2856_/D vssd1 vssd1 vccd1 vccd1 _2856_/Q sky130_fd_sc_hd__dfxtp_1
X_2925_ _2951_/CLK _2925_/D vssd1 vssd1 vccd1 vccd1 _2925_/Q sky130_fd_sc_hd__dfxtp_1
X_1807_ _2519_/A vssd1 vssd1 vccd1 vccd1 _2510_/A sky130_fd_sc_hd__clkbuf_2
X_1669_ _2923_/Q _2922_/Q vssd1 vssd1 vccd1 vccd1 _1669_/Y sky130_fd_sc_hd__nand2_1
X_2787_ _2948_/CLK _2787_/D vssd1 vssd1 vccd1 vccd1 _2787_/Q sky130_fd_sc_hd__dfxtp_1
X_1738_ _1735_/Y _2938_/Q _1630_/B _1737_/X vssd1 vssd1 vccd1 vccd1 _1747_/B sky130_fd_sc_hd__a31o_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2710_ _2721_/CLK _2710_/D vssd1 vssd1 vccd1 vccd1 _2710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1454_ _1457_/A _1458_/A vssd1 vssd1 vccd1 vccd1 _1459_/B sky130_fd_sc_hd__nand2_1
X_1523_ _2687_/Q _1521_/X _1522_/Y _2690_/Q vssd1 vssd1 vccd1 vccd1 _1523_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2641_ _2893_/CLK _2641_/D vssd1 vssd1 vccd1 vccd1 _2641_/Q sky130_fd_sc_hd__dfxtp_1
X_2572_ _2923_/Q _2570_/X _2571_/X vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__o21ba_1
X_1385_ _1384_/S _1385_/B vssd1 vssd1 vccd1 vccd1 _1385_/X sky130_fd_sc_hd__and2b_1
X_2006_ _2712_/Q _1995_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _2006_/X sky130_fd_sc_hd__o21ba_1
XFILLER_51_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2908_ _2923_/CLK _2908_/D vssd1 vssd1 vccd1 vccd1 _2908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2839_ _2839_/CLK _2839_/D vssd1 vssd1 vccd1 vccd1 _2839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2624_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2639_/B sky130_fd_sc_hd__clkbuf_2
X_2555_ _2919_/Q _2545_/X _2554_/X vssd1 vssd1 vccd1 vccd1 _2916_/D sky130_fd_sc_hd__o21a_1
X_2486_ _2893_/Q _2477_/X _2485_/X vssd1 vssd1 vccd1 vccd1 _2890_/D sky130_fd_sc_hd__o21a_1
X_1506_ _2843_/Q vssd1 vssd1 vccd1 vccd1 _1512_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1437_ _1433_/X _1434_/X _1435_/X _1436_/X _2850_/Q _2851_/Q vssd1 vssd1 vccd1 vccd1
+ _1438_/B sky130_fd_sc_hd__mux4_2
XFILLER_55_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1368_ _1364_/X _1365_/X _1366_/X _1367_/X _2847_/Q _2848_/Q vssd1 vssd1 vccd1 vccd1
+ _1368_/X sky130_fd_sc_hd__mux4_2
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 bi_u1y0s_L1[11] vssd1 vssd1 vccd1 vccd1 _1624_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput26 prog_done vssd1 vssd1 vccd1 vccd1 _2317_/B sky130_fd_sc_hd__clkbuf_1
X_2340_ _2400_/S vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__clkbuf_2
X_2271_ _2296_/A vssd1 vssd1 vccd1 vccd1 _2459_/B sky130_fd_sc_hd__clkbuf_2
X_1986_ _2704_/Q _1977_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__o21ba_1
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2607_ _2937_/Q _2596_/X _2597_/X vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__o21ba_1
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2538_ _2910_/Q _2532_/X _2533_/X vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__o21ba_1
X_2469_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1840_ _2650_/Q _1834_/X _1839_/X vssd1 vssd1 vccd1 vccd1 _2651_/D sky130_fd_sc_hd__o21a_1
X_1771_ _2811_/Q _2810_/Q _2151_/B _1784_/D vssd1 vssd1 vccd1 vccd1 _1771_/X sky130_fd_sc_hd__and4b_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_14_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2254_ _2254_/A vssd1 vssd1 vccd1 vccd1 _2254_/X sky130_fd_sc_hd__clkbuf_1
X_2323_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2400_/S sky130_fd_sc_hd__buf_2
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2185_ _2778_/Q _2183_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _2185_/X sky130_fd_sc_hd__o21ba_1
X_1969_ _2697_/Q _1967_/X _1968_/X vssd1 vssd1 vccd1 vccd1 _2698_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1823_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1823_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2872_ _2872_/CLK _2872_/D vssd1 vssd1 vccd1 vccd1 _2872_/Q sky130_fd_sc_hd__dfxtp_1
X_2941_ _2943_/CLK _2941_/D vssd1 vssd1 vccd1 vccd1 _2941_/Q sky130_fd_sc_hd__dfxtp_1
X_1685_ _1683_/X _1684_/X _1697_/A vssd1 vssd1 vccd1 vccd1 _1686_/S sky130_fd_sc_hd__o21ai_1
X_1754_ _2935_/Q _2934_/Q _1754_/C vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__and3b_1
X_2306_ _2345_/A vssd1 vssd1 vccd1 vccd1 _2306_/X sky130_fd_sc_hd__buf_2
X_2237_ _2796_/Q _2235_/X _2236_/X vssd1 vssd1 vccd1 vccd1 _2797_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2099_ _2786_/Q _2097_/X _2098_/X vssd1 vssd1 vccd1 vccd1 _2746_/D sky130_fd_sc_hd__o21a_1
X_2168_ _2772_/Q _2157_/X _2158_/X vssd1 vssd1 vccd1 vccd1 _2168_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1470_ _2709_/Q _1455_/Y _1469_/Y vssd1 vssd1 vccd1 vccd1 _1470_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2022_ _2053_/A vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2924_ _2943_/CLK _2924_/D vssd1 vssd1 vccd1 vccd1 _2924_/Q sky130_fd_sc_hd__dfxtp_1
X_2855_ _2858_/CLK _2855_/D vssd1 vssd1 vccd1 vccd1 _2855_/Q sky130_fd_sc_hd__dfxtp_1
X_2786_ _2948_/CLK _2786_/D vssd1 vssd1 vccd1 vccd1 _2786_/Q sky130_fd_sc_hd__dfxtp_2
X_1806_ _2807_/Q vssd1 vssd1 vccd1 vccd1 _2519_/A sky130_fd_sc_hd__clkbuf_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ _2660_/Q vssd1 vssd1 vccd1 vccd1 _1600_/A sky130_fd_sc_hd__inv_2
X_1668_ _2922_/Q _1630_/B _2923_/Q vssd1 vssd1 vccd1 vccd1 _1671_/B sky130_fd_sc_hd__a21o_1
X_1737_ _2938_/Q _1438_/B _1736_/Y _2939_/Q vssd1 vssd1 vccd1 vccd1 _1737_/X sky130_fd_sc_hd__o211a_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2640_ _2950_/CLK _2640_/D vssd1 vssd1 vccd1 vccd1 _2640_/Q sky130_fd_sc_hd__dfxtp_1
X_1522_ _1522_/A _1522_/B vssd1 vssd1 vccd1 vccd1 _1522_/Y sky130_fd_sc_hd__nor2_2
X_1453_ _1441_/X _1452_/X _2915_/Q vssd1 vssd1 vccd1 vccd1 _1458_/A sky130_fd_sc_hd__mux2_2
X_2571_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2571_/X sky130_fd_sc_hd__clkbuf_1
X_2005_ _2710_/Q _1999_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _2711_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1384_ input17/X input7/X _1384_/S vssd1 vssd1 vccd1 vccd1 _1384_/X sky130_fd_sc_hd__mux2_1
X_2907_ _2907_/CLK _2907_/D vssd1 vssd1 vccd1 vccd1 _2907_/Q sky130_fd_sc_hd__dfxtp_1
X_2838_ _2839_/CLK _2838_/D vssd1 vssd1 vccd1 vccd1 _2838_/Q sky130_fd_sc_hd__dfxtp_1
X_2769_ _2815_/CLK _2769_/D vssd1 vssd1 vccd1 vccd1 _2769_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2554_ _1663_/X _2550_/X _2551_/X vssd1 vssd1 vccd1 vccd1 _2554_/X sky130_fd_sc_hd__o21ba_1
X_2623_ _2942_/Q _2611_/X _2622_/X vssd1 vssd1 vccd1 vccd1 _2943_/D sky130_fd_sc_hd__o21a_1
X_2485_ _2890_/Q _2483_/X _2484_/X vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__o21ba_1
X_1505_ _2844_/Q vssd1 vssd1 vccd1 vccd1 _1505_/Y sky130_fd_sc_hd__inv_2
X_1367_ _1366_/S _1502_/B vssd1 vssd1 vccd1 vccd1 _1367_/X sky130_fd_sc_hd__and2b_1
X_1436_ _1435_/S _1533_/B vssd1 vssd1 vccd1 vccd1 _1436_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput16 bi_u1y0s_L1[1] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_2
Xinput27 prog_rst vssd1 vssd1 vccd1 vccd1 _2828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2270_ _2460_/A _2314_/S vssd1 vssd1 vccd1 vccd1 _2809_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1985_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2537_ _2908_/Q _2531_/X _2536_/X vssd1 vssd1 vccd1 vccd1 _2909_/D sky130_fd_sc_hd__o21a_1
X_2606_ _2939_/Q _2600_/X _2605_/X vssd1 vssd1 vccd1 vccd1 _2936_/D sky130_fd_sc_hd__o21a_1
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2399_ _1449_/B _2397_/X _2398_/Y vssd1 vssd1 vccd1 vccd1 _2856_/D sky130_fd_sc_hd__o21a_1
X_2468_ _2887_/Q _2461_/X _2467_/X vssd1 vssd1 vccd1 vccd1 _2884_/D sky130_fd_sc_hd__o21a_1
X_1419_ _2786_/Q _1417_/Y _2745_/Q _1418_/X vssd1 vssd1 vccd1 vccd1 _1736_/B sky130_fd_sc_hd__a31oi_4
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1770_ _2810_/Q vssd1 vssd1 vccd1 vccd1 _1770_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2184_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2184_/X sky130_fd_sc_hd__clkbuf_1
X_2253_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2253_/X sky130_fd_sc_hd__clkbuf_2
X_2322_ _2322_/A _2830_/Q vssd1 vssd1 vccd1 vccd1 _2444_/A sky130_fd_sc_hd__and2_1
X_1899_ _1899_/A vssd1 vssd1 vccd1 vccd1 _1899_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1968_ _2698_/Q _1959_/X _1960_/X vssd1 vssd1 vccd1 vccd1 _1968_/X sky130_fd_sc_hd__o21ba_1
XFILLER_33_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ _2943_/CLK _2940_/D vssd1 vssd1 vccd1 vccd1 _2940_/Q sky130_fd_sc_hd__dfxtp_1
X_1822_ _2615_/A vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__clkbuf_2
X_1753_ _2934_/Q _1753_/B vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__or2_1
X_2871_ _2872_/CLK _2871_/D vssd1 vssd1 vccd1 vccd1 _2871_/Q sky130_fd_sc_hd__dfxtp_1
X_1684_ _2919_/Q _2918_/Q _1754_/C vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__and3b_1
XFILLER_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2305_ _2825_/Q _2296_/X _2304_/X vssd1 vssd1 vccd1 vccd1 _2822_/D sky130_fd_sc_hd__o21a_1
X_2236_ _2797_/Q _2227_/X _2228_/X vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__o21ba_1
X_2167_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2098_ _2746_/Q _2082_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _2098_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2021_ _2716_/Q _2013_/X _2020_/X vssd1 vssd1 vccd1 vccd1 _2717_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2923_ _2923_/CLK _2923_/D vssd1 vssd1 vccd1 vccd1 _2923_/Q sky130_fd_sc_hd__dfxtp_1
X_1805_ _1820_/A vssd1 vssd1 vccd1 vccd1 _1805_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2854_ _2866_/CLK _2854_/D vssd1 vssd1 vccd1 vccd1 _2854_/Q sky130_fd_sc_hd__dfxtp_1
X_2785_ _2948_/CLK _2785_/D vssd1 vssd1 vccd1 vccd1 _2785_/Q sky130_fd_sc_hd__dfxtp_2
X_1736_ _2938_/Q _1736_/B vssd1 vssd1 vccd1 vccd1 _1736_/Y sky130_fd_sc_hd__nand2_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1598_ _2657_/Q _1598_/B _1598_/C vssd1 vssd1 vccd1 vccd1 _1598_/X sky130_fd_sc_hd__and3_1
X_1667_ _1662_/Y _1663_/X _1765_/C _1666_/X vssd1 vssd1 vccd1 vccd1 _1667_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2219_ _2791_/Q _2213_/X _2214_/X vssd1 vssd1 vccd1 vccd1 _2219_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2570_ _2614_/A vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1521_ _1522_/A _1522_/B vssd1 vssd1 vccd1 vccd1 _1521_/X sky130_fd_sc_hd__and2_1
XFILLER_58_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1452_ _1451_/X _1369_/X _2914_/Q vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__mux2_1
X_1383_ input13/X input5/X _2834_/Q vssd1 vssd1 vccd1 vccd1 _1383_/X sky130_fd_sc_hd__mux2_1
X_2004_ _2711_/Q _1995_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _2004_/X sky130_fd_sc_hd__o21ba_1
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2906_ _2946_/CLK _2906_/D vssd1 vssd1 vccd1 vccd1 _2906_/Q sky130_fd_sc_hd__dfxtp_1
X_2699_ _2914_/CLK _2699_/D vssd1 vssd1 vccd1 vccd1 _2699_/Q sky130_fd_sc_hd__dfxtp_1
X_2837_ _2839_/CLK _2837_/D vssd1 vssd1 vccd1 vccd1 _2837_/Q sky130_fd_sc_hd__dfxtp_1
X_1719_ _2751_/Q _1709_/Y _1717_/X _1718_/X vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__a211o_1
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2768_ _2815_/CLK _2768_/D vssd1 vssd1 vccd1 vccd1 _2768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_9_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2923_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1504_ _2904_/Q _1754_/C _2905_/Q vssd1 vssd1 vccd1 vccd1 _1517_/B sky130_fd_sc_hd__a21oi_1
X_2553_ _2914_/Q _2545_/X _2552_/X vssd1 vssd1 vccd1 vccd1 _2915_/D sky130_fd_sc_hd__o21a_1
X_2622_ _2943_/Q _2614_/X _2615_/X vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__o21ba_1
X_2484_ _2500_/A vssd1 vssd1 vccd1 vccd1 _2484_/X sky130_fd_sc_hd__clkbuf_1
X_1366_ input18/X input10/X _1366_/S vssd1 vssd1 vccd1 vccd1 _1366_/X sky130_fd_sc_hd__mux2_1
X_1435_ _1385_/B input12/X _1435_/S vssd1 vssd1 vccd1 vccd1 _1435_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 bi_u1y0s_L1[2] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
Xinput28 prog_we vssd1 vssd1 vccd1 vccd1 _2464_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ _1984_/A vssd1 vssd1 vccd1 vccd1 _2703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2536_ _2909_/Q _2532_/X _2533_/X vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__o21ba_1
X_2467_ _2884_/Q _2253_/X _2449_/X vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__o21ba_1
X_2605_ _2936_/Q _2596_/X _2597_/X vssd1 vssd1 vccd1 vccd1 _2605_/X sky130_fd_sc_hd__o21ba_1
XFILLER_57_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1349_ _1605_/C vssd1 vssd1 vccd1 vccd1 _1765_/C sky130_fd_sc_hd__buf_2
X_2398_ _1442_/Y _2460_/B _2293_/X vssd1 vssd1 vccd1 vccd1 _2398_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1418_ _2786_/Q _2785_/Q _2095_/C vssd1 vssd1 vccd1 vccd1 _1418_/X sky130_fd_sc_hd__and3b_2
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2321_ _2384_/A vssd1 vssd1 vccd1 vccd1 _2321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2183_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2183_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2252_ _2802_/Q _2248_/X _2251_/X vssd1 vssd1 vccd1 vccd1 _2803_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_23_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2937_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1898_ _2671_/Q _1896_/X _1897_/X vssd1 vssd1 vccd1 vccd1 _2672_/D sky130_fd_sc_hd__o21a_1
X_1967_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2519_ _2519_/A vssd1 vssd1 vccd1 vccd1 _2584_/A sky130_fd_sc_hd__buf_2
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2870_ _2875_/CLK _2870_/D vssd1 vssd1 vccd1 vccd1 _2870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1683_ _1681_/Y _2954_/A _1682_/X _2919_/Q vssd1 vssd1 vccd1 vccd1 _1683_/X sky130_fd_sc_hd__o211a_1
X_1821_ _2519_/A vssd1 vssd1 vccd1 vccd1 _2615_/A sky130_fd_sc_hd__buf_2
X_1752_ _1731_/A _1611_/B _1751_/Y vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2304_ _2822_/Q _2301_/X _2290_/X vssd1 vssd1 vccd1 vccd1 _2304_/X sky130_fd_sc_hd__o21ba_1
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2097_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2097_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2235_ _2477_/A vssd1 vssd1 vccd1 vccd1 _2235_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2166_ _2770_/Q _2154_/X _2165_/X vssd1 vssd1 vccd1 vccd1 _2771_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_1_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 repeater1/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2020_ _2717_/Q _2008_/X _2009_/X vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__o21ba_1
X_2922_ _2933_/CLK _2922_/D vssd1 vssd1 vccd1 vccd1 _2922_/Q sky130_fd_sc_hd__dfxtp_1
X_2853_ _2866_/CLK _2853_/D vssd1 vssd1 vccd1 vccd1 _2853_/Q sky130_fd_sc_hd__dfxtp_1
X_1666_ _1663_/X _1764_/B _1665_/Y _2917_/Q vssd1 vssd1 vccd1 vccd1 _1666_/X sky130_fd_sc_hd__o211a_1
X_1804_ _2482_/A vssd1 vssd1 vccd1 vccd1 _1820_/A sky130_fd_sc_hd__clkbuf_2
X_2784_ _2948_/CLK _2784_/D vssd1 vssd1 vccd1 vccd1 _2784_/Q sky130_fd_sc_hd__dfxtp_1
X_1735_ _2939_/Q vssd1 vssd1 vccd1 vccd1 _1735_/Y sky130_fd_sc_hd__inv_2
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _2641_/Q _1597_/B _1597_/C _1570_/Y vssd1 vssd1 vccd1 vccd1 _1598_/C sky130_fd_sc_hd__or4b_1
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2218_ _2789_/Q _2207_/X _2217_/X vssd1 vssd1 vccd1 vccd1 _2790_/D sky130_fd_sc_hd__o21a_1
X_2149_ _2765_/Q _2141_/X _2142_/X vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__o21ba_1
XFILLER_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1520_ _1583_/B _1520_/B vssd1 vssd1 vccd1 vccd1 _1522_/A sky130_fd_sc_hd__nand2_1
X_1451_ _1451_/A _1451_/B vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__and2_2
X_1382_ _1384_/S input1/X vssd1 vssd1 vccd1 vccd1 _1382_/X sky130_fd_sc_hd__and2_1
X_2003_ _2709_/Q _1999_/X _2002_/X vssd1 vssd1 vccd1 vccd1 _2710_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2905_ _2946_/CLK _2905_/D vssd1 vssd1 vccd1 vccd1 _2905_/Q sky130_fd_sc_hd__dfxtp_1
X_2836_ _2891_/CLK _2836_/D vssd1 vssd1 vccd1 vccd1 _2836_/Q sky130_fd_sc_hd__dfxtp_1
X_1649_ _2668_/Q _1639_/Y _1641_/Y _2669_/Q vssd1 vssd1 vccd1 vccd1 _1651_/B sky130_fd_sc_hd__a22o_1
X_2698_ _2914_/CLK _2698_/D vssd1 vssd1 vccd1 vccd1 _2698_/Q sky130_fd_sc_hd__dfxtp_1
X_1718_ _2752_/Q _1724_/B _1724_/C _1714_/A vssd1 vssd1 vccd1 vccd1 _1718_/X sky130_fd_sc_hd__a31o_1
X_2767_ _2815_/CLK _2767_/D vssd1 vssd1 vccd1 vccd1 _2767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2552_ _2915_/Q _2550_/X _2551_/X vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__o21ba_1
X_2483_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2621_ _2945_/Q _2611_/X _2620_/X vssd1 vssd1 vccd1 vccd1 _2942_/D sky130_fd_sc_hd__o21a_1
X_1503_ _1499_/X _1500_/X _1501_/X _1502_/X _2862_/Q _2863_/Q vssd1 vssd1 vccd1 vccd1
+ _1754_/C sky130_fd_sc_hd__mux4_2
XFILLER_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1365_ input13/X input6/X _2846_/Q vssd1 vssd1 vccd1 vccd1 _1365_/X sky130_fd_sc_hd__mux2_1
X_1434_ input16/X input7/X _2849_/Q vssd1 vssd1 vccd1 vccd1 _1434_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2819_ _2822_/CLK _2819_/D vssd1 vssd1 vccd1 vccd1 _2819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput18 bi_u1y0s_L1[3] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1983_ _2742_/Q _2037_/B _1983_/C vssd1 vssd1 vccd1 vccd1 _1984_/A sky130_fd_sc_hd__and3_1
X_2604_ _2934_/Q _2600_/X _2603_/X vssd1 vssd1 vccd1 vccd1 _2935_/D sky130_fd_sc_hd__o21a_1
X_2535_ _2911_/Q _2531_/X _2534_/X vssd1 vssd1 vccd1 vccd1 _2908_/D sky130_fd_sc_hd__o21a_1
X_2466_ _2466_/A vssd1 vssd1 vccd1 vccd1 _2883_/D sky130_fd_sc_hd__clkbuf_1
X_1417_ _2785_/Q vssd1 vssd1 vccd1 vccd1 _1417_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1348_ _2854_/Q _1344_/Y _1347_/Y vssd1 vssd1 vccd1 vccd1 _1605_/C sky130_fd_sc_hd__a21oi_4
X_2397_ _2439_/A vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2251_ _2803_/Q _2240_/X _2241_/X vssd1 vssd1 vccd1 vccd1 _2251_/X sky130_fd_sc_hd__o21ba_1
X_2320_ _2364_/A vssd1 vssd1 vccd1 vccd1 _2384_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2182_ _2776_/Q _2180_/X _2181_/X vssd1 vssd1 vccd1 vccd1 _2777_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1966_ _2696_/Q _1954_/X _1965_/X vssd1 vssd1 vccd1 vccd1 _2697_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1897_ _2672_/Q _1886_/X _1887_/X vssd1 vssd1 vccd1 vccd1 _1897_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2518_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2518_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2449_ _2500_/A vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1820_ _1820_/A vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1682_ _2918_/Q _1753_/B vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__or2_1
X_1751_ _2934_/Q vssd1 vssd1 vccd1 vccd1 _1751_/Y sky130_fd_sc_hd__inv_2
X_2303_ _2820_/Q _2296_/X _2302_/X vssd1 vssd1 vccd1 vccd1 _2821_/D sky130_fd_sc_hd__o21a_1
X_2234_ _2795_/Q _2222_/X _2233_/X vssd1 vssd1 vccd1 vccd1 _2796_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2165_ _2771_/Q _2157_/X _2158_/X vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__o21ba_1
X_2096_ _2096_/A vssd1 vssd1 vccd1 vccd1 _2745_/D sky130_fd_sc_hd__clkbuf_1
X_1949_ _2689_/Q _1941_/X _1948_/X vssd1 vssd1 vccd1 vccd1 _2690_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2921_ _2923_/CLK _2921_/D vssd1 vssd1 vccd1 vccd1 _2921_/Q sky130_fd_sc_hd__dfxtp_1
X_1803_ _2322_/A _2883_/Q vssd1 vssd1 vccd1 vccd1 _2482_/A sky130_fd_sc_hd__and2_1
X_2783_ _2948_/CLK _2783_/D vssd1 vssd1 vccd1 vccd1 _2783_/Q sky130_fd_sc_hd__dfxtp_1
X_2852_ _2866_/CLK _2852_/D vssd1 vssd1 vccd1 vccd1 _2852_/Q sky130_fd_sc_hd__dfxtp_1
X_1596_ _1591_/X _1594_/X _1595_/X _1597_/B vssd1 vssd1 vccd1 vccd1 _1596_/X sky130_fd_sc_hd__a211o_1
X_1665_ _2916_/Q _1786_/A vssd1 vssd1 vccd1 vccd1 _1665_/Y sky130_fd_sc_hd__nand2_1
X_1734_ _1734_/A vssd1 vssd1 vccd1 vccd1 _2037_/C sky130_fd_sc_hd__clkbuf_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2217_ _2790_/Q _2213_/X _2214_/X vssd1 vssd1 vccd1 vccd1 _2217_/X sky130_fd_sc_hd__o21ba_1
X_2079_ _2738_/Q _2066_/X _2078_/X vssd1 vssd1 vccd1 vccd1 _2739_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2148_ _2763_/Q _2137_/X _2147_/X vssd1 vssd1 vccd1 vccd1 _2764_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1450_ _2856_/Q _1448_/X _1449_/X _2857_/Q vssd1 vssd1 vccd1 vccd1 _1451_/B sky130_fd_sc_hd__a211o_1
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1381_ _2834_/Q vssd1 vssd1 vccd1 vccd1 _1384_/S sky130_fd_sc_hd__clkbuf_2
X_2002_ _2710_/Q _1995_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__o21ba_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2904_ _2907_/CLK _2904_/D vssd1 vssd1 vccd1 vccd1 _2904_/Q sky130_fd_sc_hd__dfxtp_1
X_2835_ _2858_/CLK _2835_/D vssd1 vssd1 vccd1 vccd1 _2835_/Q sky130_fd_sc_hd__dfxtp_1
X_2766_ _2766_/CLK _2766_/D vssd1 vssd1 vccd1 vccd1 _2766_/Q sky130_fd_sc_hd__dfxtp_1
X_1648_ _1657_/S vssd1 vssd1 vccd1 vccd1 _1651_/A sky130_fd_sc_hd__clkinv_2
X_2697_ _2914_/CLK _2697_/D vssd1 vssd1 vccd1 vccd1 _2697_/Q sky130_fd_sc_hd__dfxtp_1
X_1717_ _2750_/Q _1708_/Y _1716_/X _2753_/Q vssd1 vssd1 vccd1 vccd1 _1717_/X sky130_fd_sc_hd__a22o_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _2889_/Q _1562_/X _1563_/Y _1564_/X _1698_/B vssd1 vssd1 vccd1 vccd1 _1584_/C
+ sky130_fd_sc_hd__a32oi_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2620_ _2942_/Q _2614_/X _2615_/X vssd1 vssd1 vccd1 vccd1 _2620_/X sky130_fd_sc_hd__o21ba_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2551_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2551_/X sky130_fd_sc_hd__clkbuf_1
X_2482_ _2482_/A vssd1 vssd1 vccd1 vccd1 _2550_/A sky130_fd_sc_hd__clkbuf_2
X_1433_ _1435_/S input4/X vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__and2_1
X_1502_ _1501_/S _1502_/B vssd1 vssd1 vccd1 vccd1 _1502_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_prog_clk clkbuf_2_1_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2933_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1364_ _1366_/S input1/X vssd1 vssd1 vccd1 vccd1 _1364_/X sky130_fd_sc_hd__and2_1
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2749_ _2755_/CLK _2749_/D vssd1 vssd1 vccd1 vccd1 _2749_/Q sky130_fd_sc_hd__dfxtp_1
X_2818_ _2933_/CLK _2818_/D vssd1 vssd1 vccd1 vccd1 _2818_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 bi_u1y0s_L1[4] vssd1 vssd1 vccd1 vccd1 _1385_/B sky130_fd_sc_hd__clkbuf_2
X_1982_ _2701_/Q _1967_/X _1981_/X vssd1 vssd1 vccd1 vccd1 _2702_/D sky130_fd_sc_hd__o21a_1
X_2534_ _2908_/Q _2532_/X _2533_/X vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__o21ba_1
X_2603_ _2935_/Q _2596_/X _2597_/X vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__o21ba_1
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1416_ _2269_/A vssd1 vssd1 vccd1 vccd1 _1420_/A sky130_fd_sc_hd__buf_2
X_2465_ _2268_/A _2633_/S vssd1 vssd1 vccd1 vccd1 _2466_/A sky130_fd_sc_hd__and2b_1
X_1347_ _2853_/Q _1345_/X _1346_/X vssd1 vssd1 vccd1 vccd1 _1347_/Y sky130_fd_sc_hd__a21oi_1
X_2396_ _2860_/Q _2384_/X _2395_/X vssd1 vssd1 vccd1 vccd1 _2855_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ _2801_/Q _2248_/X _2249_/X vssd1 vssd1 vccd1 vccd1 _2802_/D sky130_fd_sc_hd__o21a_1
X_2181_ _2777_/Q _2170_/X _2171_/X vssd1 vssd1 vccd1 vccd1 _2181_/X sky130_fd_sc_hd__o21ba_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1965_ _2697_/Q _1959_/X _1960_/X vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__o21ba_1
X_1896_ _1927_/A vssd1 vssd1 vccd1 vccd1 _1896_/X sky130_fd_sc_hd__clkbuf_2
X_2517_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2379_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2379_/X sky130_fd_sc_hd__clkbuf_1
X_2448_ _2874_/Q _2439_/X _2447_/X vssd1 vssd1 vccd1 vccd1 _2875_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1750_ _2773_/Q _1745_/X _1746_/Y _2771_/Q _1749_/X vssd1 vssd1 vccd1 vccd1 _1750_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1681_ _2918_/Q vssd1 vssd1 vccd1 vccd1 _1681_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2302_ _2821_/Q _2301_/X _2290_/X vssd1 vssd1 vccd1 vccd1 _2302_/X sky130_fd_sc_hd__o21ba_1
X_2233_ _2796_/Q _2227_/X _2228_/X vssd1 vssd1 vccd1 vccd1 _2233_/X sky130_fd_sc_hd__o21ba_1
X_2164_ _2769_/Q _2154_/X _2163_/X vssd1 vssd1 vccd1 vccd1 _2770_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2095_ _2784_/Q _2151_/B _2095_/C vssd1 vssd1 vccd1 vccd1 _2096_/A sky130_fd_sc_hd__and3_1
X_1948_ _2690_/Q _1946_/X _1947_/X vssd1 vssd1 vccd1 vccd1 _1948_/X sky130_fd_sc_hd__o21ba_1
X_1879_ _2665_/Q _1873_/X _1874_/X vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2920_ _2923_/CLK _2920_/D vssd1 vssd1 vccd1 vccd1 _2920_/Q sky130_fd_sc_hd__dfxtp_1
X_1802_ _1849_/A vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2782_ _2948_/CLK _2782_/D vssd1 vssd1 vccd1 vccd1 _2782_/Q sky130_fd_sc_hd__dfxtp_1
X_2851_ _2866_/CLK _2851_/D vssd1 vssd1 vccd1 vccd1 _2851_/Q sky130_fd_sc_hd__dfxtp_1
X_1733_ _2762_/Q _2037_/B _1733_/C vssd1 vssd1 vccd1 vccd1 _1734_/A sky130_fd_sc_hd__and3_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _2645_/Q _1575_/Y _1570_/Y vssd1 vssd1 vccd1 vccd1 _1595_/X sky130_fd_sc_hd__o21a_1
X_1664_ _1664_/A vssd1 vssd1 vccd1 vccd1 _1786_/A sky130_fd_sc_hd__buf_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2216_ _2788_/Q _2207_/X _2215_/X vssd1 vssd1 vccd1 vccd1 _2789_/D sky130_fd_sc_hd__o21a_1
X_2147_ _2764_/Q _2141_/X _2142_/X vssd1 vssd1 vccd1 vccd1 _2147_/X sky130_fd_sc_hd__o21ba_1
X_2078_ _2739_/Q _2068_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _2078_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1380_ _2940_/Q _1380_/B vssd1 vssd1 vccd1 vccd1 _1380_/X sky130_fd_sc_hd__and2_1
X_2001_ _2708_/Q _1999_/X _2000_/X vssd1 vssd1 vccd1 vccd1 _2709_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2903_ _2946_/CLK _2903_/D vssd1 vssd1 vccd1 vccd1 _2903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2696_ _2914_/CLK _2696_/D vssd1 vssd1 vccd1 vccd1 _2696_/Q sky130_fd_sc_hd__dfxtp_1
X_1716_ _1747_/A _1716_/B _1716_/C vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__and3_1
X_2834_ _2858_/CLK _2834_/D vssd1 vssd1 vccd1 vccd1 _2834_/Q sky130_fd_sc_hd__dfxtp_1
X_2765_ _2765_/CLK _2765_/D vssd1 vssd1 vccd1 vccd1 _2765_/Q sky130_fd_sc_hd__dfxtp_1
X_1647_ _1657_/S _1647_/B _1647_/C vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__or3_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1578_ _1593_/B _1593_/C _1589_/D vssd1 vssd1 vccd1 vccd1 _1578_/X sky130_fd_sc_hd__and3_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2550_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2550_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2481_ _2888_/Q _2477_/X _2480_/X vssd1 vssd1 vccd1 vccd1 _2889_/D sky130_fd_sc_hd__o21a_1
X_1363_ _2846_/Q vssd1 vssd1 vccd1 vccd1 _1366_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_1432_ _2849_/Q vssd1 vssd1 vccd1 vccd1 _1435_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_1501_ input18/X input10/X _1501_/S vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__mux2_1
X_2679_ _2687_/CLK _2679_/D vssd1 vssd1 vccd1 vccd1 _2679_/Q sky130_fd_sc_hd__dfxtp_1
X_2748_ _2822_/CLK _2748_/D vssd1 vssd1 vccd1 vccd1 _2748_/Q sky130_fd_sc_hd__dfxtp_1
X_2817_ _2822_/CLK _2817_/D vssd1 vssd1 vccd1 vccd1 _2817_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1981_ _2702_/Q _1977_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__o21ba_1
XFILLER_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2533_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__clkbuf_1
X_2602_ _2937_/Q _2600_/X _2601_/Y vssd1 vssd1 vccd1 vccd1 _2934_/D sky130_fd_sc_hd__o21a_1
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2464_ _2464_/A _2464_/B vssd1 vssd1 vccd1 vccd1 _2633_/S sky130_fd_sc_hd__and2_1
X_1346_ _1340_/Y _1345_/S input5/X _2854_/Q vssd1 vssd1 vccd1 vccd1 _1346_/X sky130_fd_sc_hd__a31o_1
X_2395_ _1449_/B _2387_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _2395_/X sky130_fd_sc_hd__o21ba_1
X_1415_ _2322_/A vssd1 vssd1 vccd1 vccd1 _2269_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_2_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2893_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2180_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1895_ _2670_/Q _1883_/X _1894_/X vssd1 vssd1 vccd1 vccd1 _2671_/D sky130_fd_sc_hd__o21a_1
X_1964_ _2695_/Q _1954_/X _1963_/X vssd1 vssd1 vccd1 vccd1 _2696_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2516_ _2905_/Q _2505_/X _2515_/X vssd1 vssd1 vccd1 vccd1 _2902_/D sky130_fd_sc_hd__o21a_1
X_2447_ _2875_/Q _2444_/X _2436_/X vssd1 vssd1 vccd1 vccd1 _2447_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1329_ _2949_/Q vssd1 vssd1 vccd1 vccd1 _1583_/B sky130_fd_sc_hd__clkbuf_2
X_2378_ _2847_/Q _2370_/X _2377_/X vssd1 vssd1 vccd1 vccd1 _2848_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1680_ _2725_/Q _2726_/Q _2727_/Q _2728_/Q _1672_/X _1692_/B vssd1 vssd1 vccd1 vccd1
+ _1680_/X sky130_fd_sc_hd__mux4_1
X_2301_ _2301_/A vssd1 vssd1 vccd1 vccd1 _2301_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2232_ _2794_/Q _2222_/X _2231_/X vssd1 vssd1 vccd1 vccd1 _2795_/D sky130_fd_sc_hd__o21a_1
X_2163_ _2770_/Q _2157_/X _2158_/X vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__o21ba_1
XFILLER_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2094_ _2743_/Q _2081_/X _2093_/X vssd1 vssd1 vccd1 vccd1 _2744_/D sky130_fd_sc_hd__o21a_1
X_1947_ _1960_/A vssd1 vssd1 vccd1 vccd1 _1947_/X sky130_fd_sc_hd__clkbuf_1
X_1878_ _2663_/Q _1870_/X _1877_/X vssd1 vssd1 vccd1 vccd1 _2664_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2850_ _2866_/CLK _2850_/D vssd1 vssd1 vccd1 vccd1 _2850_/Q sky130_fd_sc_hd__dfxtp_1
X_1663_ _2916_/Q vssd1 vssd1 vccd1 vccd1 _1663_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1801_ _2560_/A vssd1 vssd1 vccd1 vccd1 _1849_/A sky130_fd_sc_hd__clkbuf_4
X_1732_ _1720_/X _1727_/X _1732_/S vssd1 vssd1 vccd1 vccd1 _1733_/C sky130_fd_sc_hd__mux2_1
X_2781_ _2781_/CLK _2781_/D vssd1 vssd1 vccd1 vccd1 _2781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _2643_/Q _1581_/Y _1592_/X _1593_/X vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__a211o_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2077_ _2737_/Q _2066_/X _2076_/X vssd1 vssd1 vccd1 vccd1 _2738_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2215_ _2789_/Q _2213_/X _2214_/X vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__o21ba_1
X_2146_ _2762_/Q _2137_/X _2145_/X vssd1 vssd1 vccd1 vccd1 _2763_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2000_ _2709_/Q _1995_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _2000_/X sky130_fd_sc_hd__o21ba_1
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2902_ _2946_/CLK _2902_/D vssd1 vssd1 vccd1 vccd1 _2902_/Q sky130_fd_sc_hd__dfxtp_1
X_2833_ _2839_/CLK _2833_/D vssd1 vssd1 vccd1 vccd1 _2833_/Q sky130_fd_sc_hd__dfxtp_1
X_2695_ _2881_/CLK _2695_/D vssd1 vssd1 vccd1 vccd1 _2695_/Q sky130_fd_sc_hd__dfxtp_1
X_1646_ _2675_/Q _1644_/Y _1645_/Y _2674_/Q vssd1 vssd1 vccd1 vccd1 _1647_/C sky130_fd_sc_hd__a22o_1
X_1715_ _2746_/Q _1708_/Y _1709_/Y _2747_/Q _1727_/S vssd1 vssd1 vccd1 vccd1 _1715_/X
+ sky130_fd_sc_hd__a221o_1
X_2764_ _2815_/CLK _2764_/D vssd1 vssd1 vccd1 vccd1 _2764_/Q sky130_fd_sc_hd__dfxtp_2
X_1577_ _2949_/Q vssd1 vssd1 vccd1 vccd1 _1593_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2129_ _2757_/Q _2126_/X _2128_/X vssd1 vssd1 vccd1 vccd1 _2129_/X sky130_fd_sc_hd__o21ba_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2480_ _2889_/Q _2469_/X _2470_/X vssd1 vssd1 vccd1 vccd1 _2480_/X sky130_fd_sc_hd__o21ba_1
X_1500_ input13/X input6/X _2861_/Q vssd1 vssd1 vccd1 vccd1 _1500_/X sky130_fd_sc_hd__mux2_1
X_1431_ _1431_/A vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__clkbuf_4
X_1362_ _2944_/Q _1698_/B vssd1 vssd1 vccd1 vccd1 _1362_/X sky130_fd_sc_hd__and2_1
XFILLER_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2816_ _2822_/CLK _2816_/D vssd1 vssd1 vccd1 vccd1 _2816_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_prog_clk clkbuf_2_0_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2949_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2678_ _2687_/CLK _2678_/D vssd1 vssd1 vccd1 vccd1 _2678_/Q sky130_fd_sc_hd__dfxtp_1
X_2747_ _2822_/CLK _2747_/D vssd1 vssd1 vccd1 vccd1 _2747_/Q sky130_fd_sc_hd__dfxtp_1
X_1629_ _2875_/Q _1625_/Y _1628_/Y vssd1 vssd1 vccd1 vccd1 _1630_/B sky130_fd_sc_hd__a21oi_4
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1980_ _2041_/A vssd1 vssd1 vccd1 vccd1 _1980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2532_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2532_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2463_ _2885_/Q _2461_/X _2462_/X vssd1 vssd1 vccd1 vccd1 _2882_/D sky130_fd_sc_hd__o21a_1
X_2601_ _1751_/Y _2542_/X _2313_/X vssd1 vssd1 vccd1 vccd1 _2601_/Y sky130_fd_sc_hd__a21oi_1
X_1414_ _1581_/A vssd1 vssd1 vccd1 vccd1 _2322_/A sky130_fd_sc_hd__clkbuf_2
X_2394_ _2853_/Q _2384_/X _2393_/X vssd1 vssd1 vccd1 vccd1 _2854_/D sky130_fd_sc_hd__o21a_1
X_1345_ input17/X input8/X _1345_/S vssd1 vssd1 vccd1 vccd1 _1345_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1894_ _2671_/Q _1886_/X _1887_/X vssd1 vssd1 vccd1 vccd1 _1894_/X sky130_fd_sc_hd__o21ba_1
X_1963_ _2696_/Q _1959_/X _1960_/X vssd1 vssd1 vccd1 vccd1 _1963_/X sky130_fd_sc_hd__o21ba_1
X_2515_ _2902_/Q _2499_/X _2500_/X vssd1 vssd1 vccd1 vccd1 _2515_/X sky130_fd_sc_hd__o21ba_1
X_2446_ _1626_/S _2439_/X _2445_/X vssd1 vssd1 vccd1 vccd1 _2874_/D sky130_fd_sc_hd__o21a_1
X_1328_ _1328_/A vssd1 vssd1 vccd1 vccd1 _1328_/Y sky130_fd_sc_hd__inv_2
X_2377_ _2848_/Q _2374_/X _2359_/X vssd1 vssd1 vccd1 vccd1 _2377_/X sky130_fd_sc_hd__o21ba_1
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2300_ _2823_/Q _2296_/X _2299_/X vssd1 vssd1 vccd1 vccd1 _2820_/D sky130_fd_sc_hd__o21a_1
X_2231_ _2795_/Q _2227_/X _2228_/X vssd1 vssd1 vccd1 vccd1 _2231_/X sky130_fd_sc_hd__o21ba_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2093_ _2744_/Q _2082_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _2093_/X sky130_fd_sc_hd__o21ba_1
X_2162_ _2768_/Q _2154_/X _2161_/X vssd1 vssd1 vccd1 vccd1 _2769_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1946_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1946_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1877_ _2664_/Q _1873_/X _1874_/X vssd1 vssd1 vccd1 vccd1 _1877_/X sky130_fd_sc_hd__o21ba_1
X_2429_ _1492_/S _2425_/X _2428_/X vssd1 vssd1 vccd1 vccd1 _2868_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1800_ _1868_/A vssd1 vssd1 vccd1 vccd1 _2560_/A sky130_fd_sc_hd__clkbuf_2
X_1662_ _2917_/Q vssd1 vssd1 vccd1 vccd1 _1662_/Y sky130_fd_sc_hd__inv_2
X_1731_ _1731_/A _1731_/B _1731_/C vssd1 vssd1 vccd1 vccd1 _1732_/S sky130_fd_sc_hd__and3_1
X_2780_ _2781_/CLK _2780_/D vssd1 vssd1 vccd1 vccd1 _2780_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _2644_/Q _1593_/B _1593_/C _1593_/D vssd1 vssd1 vccd1 vccd1 _1593_/X sky130_fd_sc_hd__and4_1
X_2214_ _2254_/A vssd1 vssd1 vccd1 vccd1 _2214_/X sky130_fd_sc_hd__clkbuf_1
X_2076_ _2738_/Q _2068_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__o21ba_1
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2145_ _2763_/Q _2141_/X _2142_/X vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__o21ba_1
X_1929_ _2723_/Q _1927_/X _1928_/X vssd1 vssd1 vccd1 vccd1 _2683_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2901_ _2946_/CLK _2901_/D vssd1 vssd1 vccd1 vccd1 _2901_/Q sky130_fd_sc_hd__dfxtp_1
X_2832_ _2893_/CLK _2832_/D vssd1 vssd1 vccd1 vccd1 _2832_/Q sky130_fd_sc_hd__dfxtp_1
X_2763_ _2815_/CLK _2763_/D vssd1 vssd1 vccd1 vccd1 _2763_/Q sky130_fd_sc_hd__dfxtp_1
X_2694_ _2881_/CLK _2694_/D vssd1 vssd1 vccd1 vccd1 _2694_/Q sky130_fd_sc_hd__dfxtp_1
X_1645_ _1645_/A _1645_/B vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__nor2_2
X_1576_ _2653_/Q _1570_/Y _1575_/Y vssd1 vssd1 vccd1 vccd1 _1576_/X sky130_fd_sc_hd__a21o_1
X_1714_ _1714_/A vssd1 vssd1 vccd1 vccd1 _1727_/S sky130_fd_sc_hd__inv_2
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ _2730_/Q _2052_/X _2058_/X vssd1 vssd1 vccd1 vccd1 _2731_/D sky130_fd_sc_hd__o21a_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2128_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2128_/X sky130_fd_sc_hd__clkbuf_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1430_ _1598_/B _1430_/B vssd1 vssd1 vccd1 vccd1 _1431_/A sky130_fd_sc_hd__and2_1
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1361_ _1357_/X _1360_/X _2872_/Q vssd1 vssd1 vccd1 vccd1 _1698_/B sky130_fd_sc_hd__mux2_4
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2746_ _2755_/CLK _2746_/D vssd1 vssd1 vccd1 vccd1 _2746_/Q sky130_fd_sc_hd__dfxtp_1
X_2815_ _2815_/CLK _2815_/D vssd1 vssd1 vccd1 vccd1 _2815_/Q sky130_fd_sc_hd__dfxtp_1
X_2677_ _2677_/CLK _2677_/D vssd1 vssd1 vccd1 vccd1 _2677_/Q sky130_fd_sc_hd__dfxtp_1
X_1559_ _2884_/Q _1754_/C _2885_/Q vssd1 vssd1 vccd1 vccd1 _1559_/X sky130_fd_sc_hd__a21o_1
X_1628_ _2874_/Q _1626_/X _1627_/X vssd1 vssd1 vccd1 vccd1 _1628_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2600_ _2611_/A vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__clkbuf_2
X_1413_ _2949_/Q vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__inv_2
X_2531_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__clkbuf_2
X_2462_ _2882_/Q _2253_/X _2449_/X vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__o21ba_1
X_2393_ _2854_/Q _2387_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _2393_/X sky130_fd_sc_hd__o21ba_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1344_ _1340_/Y _1341_/X _1343_/X vssd1 vssd1 vccd1 vccd1 _1344_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2729_ _2739_/CLK _2729_/D vssd1 vssd1 vccd1 vccd1 _2729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1962_ _2694_/Q _1954_/X _1961_/X vssd1 vssd1 vccd1 vccd1 _2695_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1893_ _2669_/Q _1883_/X _1892_/X vssd1 vssd1 vccd1 vccd1 _2670_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2514_ _2900_/Q _2505_/X _2513_/X vssd1 vssd1 vccd1 vccd1 _2901_/D sky130_fd_sc_hd__o21a_1
X_2445_ _2874_/Q _2444_/X _2436_/X vssd1 vssd1 vccd1 vccd1 _2445_/X sky130_fd_sc_hd__o21ba_1
X_2376_ _1366_/S _2370_/X _2375_/X vssd1 vssd1 vccd1 vccd1 _2847_/D sky130_fd_sc_hd__o21a_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1327_ _1318_/X _1326_/X _2943_/Q vssd1 vssd1 vccd1 vccd1 _1328_/A sky130_fd_sc_hd__mux2_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xclkbuf_leaf_10_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2914_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2230_ _2793_/Q _2222_/X _2229_/X vssd1 vssd1 vccd1 vccd1 _2794_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2092_ _2742_/Q _2081_/X _2091_/Y vssd1 vssd1 vccd1 vccd1 _2743_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2161_ _2769_/Q _2157_/X _2158_/X vssd1 vssd1 vccd1 vccd1 _2161_/X sky130_fd_sc_hd__o21ba_1
X_1945_ _2688_/Q _1941_/X _1944_/X vssd1 vssd1 vccd1 vccd1 _2689_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1876_ _2662_/Q _1870_/X _1875_/X vssd1 vssd1 vccd1 vccd1 _2663_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2428_ _2868_/Q _2417_/X _2422_/X vssd1 vssd1 vccd1 vccd1 _2428_/X sky130_fd_sc_hd__o21ba_1
X_2359_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2359_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1661_ _1486_/Y _2680_/Q _1796_/B _1660_/X vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__a31o_2
X_1592_ _2642_/Q _1593_/B _1584_/C _1593_/D _1597_/C vssd1 vssd1 vccd1 vccd1 _1592_/X
+ sky130_fd_sc_hd__a41o_1
X_1730_ _2924_/Q _1467_/B _1729_/Y _1784_/D vssd1 vssd1 vccd1 vccd1 _1731_/C sky130_fd_sc_hd__o22a_1
XFILLER_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2213_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2144_ _2761_/Q _2137_/X _2143_/X vssd1 vssd1 vccd1 vccd1 _2762_/D sky130_fd_sc_hd__o21a_1
X_2075_ _2736_/Q _2066_/X _2074_/X vssd1 vssd1 vccd1 vccd1 _2737_/D sky130_fd_sc_hd__o21a_1
X_1928_ _2683_/Q _1915_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _1928_/X sky130_fd_sc_hd__o21ba_1
X_1859_ _2658_/Q _1849_/X _1858_/X vssd1 vssd1 vccd1 vccd1 _2659_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_prog_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2900_ _2946_/CLK _2900_/D vssd1 vssd1 vccd1 vccd1 _2900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2831_ _2893_/CLK _2831_/D vssd1 vssd1 vccd1 vccd1 _2831_/Q sky130_fd_sc_hd__dfxtp_1
X_1713_ _2322_/A _1713_/B _1712_/X vssd1 vssd1 vccd1 vccd1 _1714_/A sky130_fd_sc_hd__or3b_2
X_2762_ _2765_/CLK _2762_/D vssd1 vssd1 vccd1 vccd1 _2762_/Q sky130_fd_sc_hd__dfxtp_1
X_2693_ _2881_/CLK _2693_/D vssd1 vssd1 vccd1 vccd1 _2693_/Q sky130_fd_sc_hd__dfxtp_1
X_1644_ _1645_/A _1644_/B vssd1 vssd1 vccd1 vccd1 _1644_/Y sky130_fd_sc_hd__nor2_2
X_1575_ _2887_/Q _1572_/X _1753_/B _1572_/A _1574_/X vssd1 vssd1 vccd1 vccd1 _1575_/Y
+ sky130_fd_sc_hd__o221ai_4
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_0 _2306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2184_/A sky130_fd_sc_hd__clkbuf_2
X_2058_ _2731_/Q _2053_/X _2055_/X vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__o21ba_1
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1360_ _1358_/X _1359_/X _2871_/Q vssd1 vssd1 vccd1 vccd1 _1360_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2676_ _2677_/CLK _2676_/D vssd1 vssd1 vccd1 vccd1 _2676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2745_ _2766_/CLK _2745_/D vssd1 vssd1 vccd1 vccd1 _2745_/Q sky130_fd_sc_hd__dfxtp_1
X_2814_ _2815_/CLK _2814_/D vssd1 vssd1 vccd1 vccd1 _2814_/Q sky130_fd_sc_hd__dfxtp_1
X_1558_ _1430_/B _1557_/Y _2949_/Q vssd1 vssd1 vccd1 vccd1 _1558_/X sky130_fd_sc_hd__o21a_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _2867_/Q vssd1 vssd1 vccd1 vccd1 _1492_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_1627_ _1621_/Y _1626_/S input6/X _2875_/Q vssd1 vssd1 vccd1 vccd1 _1627_/X sky130_fd_sc_hd__a31o_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2530_ _2906_/Q _2517_/X _2529_/X vssd1 vssd1 vccd1 vccd1 _2907_/D sky130_fd_sc_hd__o21a_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2461_ _2477_/A vssd1 vssd1 vccd1 vccd1 _2461_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2392_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2392_/X sky130_fd_sc_hd__clkbuf_1
X_1343_ _1345_/S _1551_/B _2853_/Q vssd1 vssd1 vccd1 vccd1 _1343_/X sky130_fd_sc_hd__and3b_1
X_1412_ _1311_/X _1404_/X _1778_/A vssd1 vssd1 vccd1 vccd1 _2958_/A sky130_fd_sc_hd__o21a_4
XFILLER_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2659_ _2687_/CLK _2659_/D vssd1 vssd1 vccd1 vccd1 _2659_/Q sky130_fd_sc_hd__dfxtp_2
X_2728_ _2739_/CLK _2728_/D vssd1 vssd1 vccd1 vccd1 _2728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1892_ _2670_/Q _1886_/X _1887_/X vssd1 vssd1 vccd1 vccd1 _1892_/X sky130_fd_sc_hd__o21ba_1
X_1961_ _2695_/Q _1959_/X _1960_/X vssd1 vssd1 vccd1 vccd1 _1961_/X sky130_fd_sc_hd__o21ba_1
X_2513_ _2901_/Q _2499_/X _2500_/X vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__o21ba_1
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1326_ _1613_/B _1784_/D _2942_/Q vssd1 vssd1 vccd1 vccd1 _1326_/X sky130_fd_sc_hd__mux2_1
X_2444_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2444_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2375_ _2847_/Q _2374_/X _2359_/X vssd1 vssd1 vccd1 vccd1 _2375_/X sky130_fd_sc_hd__o21ba_1
XFILLER_24_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2160_ _2767_/Q _2154_/X _2159_/X vssd1 vssd1 vccd1 vccd1 _2768_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_prog_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_2091_ _1427_/Y _2090_/X _1972_/X vssd1 vssd1 vccd1 vccd1 _2091_/Y sky130_fd_sc_hd__a21oi_1
X_1944_ _2689_/Q _1932_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _1944_/X sky130_fd_sc_hd__o21ba_1
X_1875_ _2663_/Q _1873_/X _1874_/X vssd1 vssd1 vccd1 vccd1 _1875_/X sky130_fd_sc_hd__o21ba_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2427_ _2872_/Q _2425_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _2867_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2289_ _2819_/Q _2282_/X _2288_/X vssd1 vssd1 vccd1 vccd1 _2816_/D sky130_fd_sc_hd__o21a_1
X_2358_ _2519_/A vssd1 vssd1 vccd1 vccd1 _2422_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _2680_/Q _2640_/Q _2681_/Q vssd1 vssd1 vccd1 vccd1 _1660_/X sky130_fd_sc_hd__and3b_1
X_1591_ _2647_/Q _1581_/Y _1589_/X _1590_/X vssd1 vssd1 vccd1 vccd1 _1591_/X sky130_fd_sc_hd__a211o_1
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2212_ _2212_/A vssd1 vssd1 vccd1 vccd1 _2469_/A sky130_fd_sc_hd__clkbuf_2
X_2143_ _2762_/Q _2141_/X _2142_/X vssd1 vssd1 vccd1 vccd1 _2143_/X sky130_fd_sc_hd__o21ba_1
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2074_ _2737_/Q _2068_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _2074_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1927_ _1927_/A vssd1 vssd1 vccd1 vccd1 _1927_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1858_ _2659_/Q _1850_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _1858_/X sky130_fd_sc_hd__o21ba_1
X_1789_ _2822_/Q _1786_/A _2823_/Q vssd1 vssd1 vccd1 vccd1 _1791_/B sky130_fd_sc_hd__o21ai_1
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2830_ _2943_/CLK _2830_/D vssd1 vssd1 vccd1 vccd1 _2830_/Q sky130_fd_sc_hd__dfxtp_1
X_2692_ _2881_/CLK _2692_/D vssd1 vssd1 vccd1 vccd1 _2692_/Q sky130_fd_sc_hd__dfxtp_1
X_1643_ _1643_/A _1643_/B vssd1 vssd1 vccd1 vccd1 _1645_/A sky130_fd_sc_hd__and2_1
X_1712_ _2926_/Q _1613_/B _1430_/B _1711_/Y vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__o22a_1
X_2761_ _2765_/CLK _2761_/D vssd1 vssd1 vccd1 vccd1 _2761_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 _1792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _2959_/A _1573_/Y _2949_/Q vssd1 vssd1 vccd1 vccd1 _1574_/X sky130_fd_sc_hd__o21a_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2057_ _2729_/Q _2052_/X _2056_/X vssd1 vssd1 vccd1 vccd1 _2730_/D sky130_fd_sc_hd__o21a_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _2126_/A vssd1 vssd1 vccd1 vccd1 _2126_/X sky130_fd_sc_hd__clkbuf_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2959_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2959_/X sky130_fd_sc_hd__clkbuf_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_prog_clk clkbuf_2_2_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2677_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2813_ _2948_/CLK _2813_/D vssd1 vssd1 vccd1 vccd1 _2813_/Q sky130_fd_sc_hd__dfxtp_1
X_2675_ _2677_/CLK _2675_/D vssd1 vssd1 vccd1 vccd1 _2675_/Q sky130_fd_sc_hd__dfxtp_1
X_2744_ _2755_/CLK _2744_/D vssd1 vssd1 vccd1 vccd1 _2744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1626_ input18/X input10/X _1626_/S vssd1 vssd1 vccd1 vccd1 _1626_/X sky130_fd_sc_hd__mux2_1
X_1488_ _2699_/Q vssd1 vssd1 vccd1 vccd1 _1867_/B sky130_fd_sc_hd__inv_2
X_1557_ _2885_/Q _2884_/Q vssd1 vssd1 vccd1 vccd1 _1557_/Y sky130_fd_sc_hd__nand2_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ _2749_/Q _2097_/X _2108_/X vssd1 vssd1 vccd1 vccd1 _2750_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2460_ _2460_/A _2460_/B vssd1 vssd1 vccd1 vccd1 _2881_/D sky130_fd_sc_hd__nor2_2
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2391_ _1345_/S _2384_/X _2390_/X vssd1 vssd1 vccd1 vccd1 _2853_/D sky130_fd_sc_hd__o21a_1
X_1411_ _2151_/B vssd1 vssd1 vccd1 vccd1 _1778_/A sky130_fd_sc_hd__clkbuf_4
X_1342_ _2852_/Q vssd1 vssd1 vccd1 vccd1 _1345_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1609_ _2701_/Q _2661_/Q _2702_/Q vssd1 vssd1 vccd1 vccd1 _1609_/Y sky130_fd_sc_hd__nand3b_1
X_2658_ _2687_/CLK _2658_/D vssd1 vssd1 vccd1 vccd1 _2658_/Q sky130_fd_sc_hd__dfxtp_1
X_2727_ _2739_/CLK _2727_/D vssd1 vssd1 vccd1 vccd1 _2727_/Q sky130_fd_sc_hd__dfxtp_1
X_2589_ _2928_/Q _2587_/X _2588_/X vssd1 vssd1 vccd1 vccd1 _2929_/D sky130_fd_sc_hd__o21a_1
XFILLER_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1891_ _2668_/Q _1883_/X _1890_/X vssd1 vssd1 vccd1 vccd1 _2669_/D sky130_fd_sc_hd__o21a_1
X_1960_ _1960_/A vssd1 vssd1 vccd1 vccd1 _1960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2512_ _2903_/Q _2505_/X _2511_/Y vssd1 vssd1 vccd1 vccd1 _2900_/D sky130_fd_sc_hd__o21a_1
X_2443_ _2878_/Q _2439_/X _2442_/X vssd1 vssd1 vccd1 vccd1 _2873_/D sky130_fd_sc_hd__o21a_1
X_2374_ _2430_/A vssd1 vssd1 vccd1 vccd1 _2374_/X sky130_fd_sc_hd__clkbuf_2
X_1325_ _2955_/A vssd1 vssd1 vccd1 vccd1 _1784_/D sky130_fd_sc_hd__buf_2
XFILLER_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2090_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2090_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1943_ _2687_/Q _1941_/X _1942_/X vssd1 vssd1 vccd1 vccd1 _2688_/D sky130_fd_sc_hd__o21a_1
X_1874_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1874_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2426_ _1492_/S _2417_/X _2422_/X vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2288_ _2816_/Q _2285_/X _2277_/X vssd1 vssd1 vccd1 vccd1 _2288_/X sky130_fd_sc_hd__o21ba_1
X_2357_ _1322_/S _2352_/X _2356_/X vssd1 vssd1 vccd1 vccd1 _2841_/D sky130_fd_sc_hd__o21a_1
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _2646_/Q _1583_/B _1584_/C _1593_/D _1575_/Y vssd1 vssd1 vccd1 vccd1 _1590_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2073_ _2735_/Q _2066_/X _2072_/X vssd1 vssd1 vccd1 vccd1 _2736_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2211_ _2787_/Q _2207_/X _2210_/X vssd1 vssd1 vccd1 vccd1 _2788_/D sky130_fd_sc_hd__o21a_1
X_2142_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1857_ _2657_/Q _1849_/X _1856_/X vssd1 vssd1 vccd1 vccd1 _2658_/D sky130_fd_sc_hd__o21a_1
X_1926_ _1926_/A vssd1 vssd1 vccd1 vccd1 _2682_/D sky130_fd_sc_hd__clkbuf_1
X_1788_ _1786_/X _1787_/X _1420_/A vssd1 vssd1 vccd1 vccd1 _1788_/Y sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_29_prog_clk clkbuf_2_0_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2866_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2409_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2409_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2691_ _2907_/CLK _2691_/D vssd1 vssd1 vccd1 vccd1 _2691_/Q sky130_fd_sc_hd__dfxtp_1
X_1642_ _2676_/Q _1639_/Y _1641_/Y _2677_/Q vssd1 vssd1 vccd1 vccd1 _1647_/B sky130_fd_sc_hd__a22o_1
X_1711_ _2927_/Q _2926_/Q vssd1 vssd1 vccd1 vccd1 _1711_/Y sky130_fd_sc_hd__nand2_1
X_2760_ _2822_/CLK _2760_/D vssd1 vssd1 vccd1 vccd1 _2760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _2887_/Q _2886_/Q vssd1 vssd1 vccd1 vccd1 _1573_/Y sky130_fd_sc_hd__nand2_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2056_ _2730_/Q _2053_/X _2055_/X vssd1 vssd1 vccd1 vccd1 _2056_/X sky130_fd_sc_hd__o21ba_1
X_2125_ _2755_/Q _2123_/X _2124_/X vssd1 vssd1 vccd1 vccd1 _2756_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1909_ _2675_/Q _1896_/X _1908_/X vssd1 vssd1 vccd1 vccd1 _2676_/D sky130_fd_sc_hd__o21a_1
X_2958_ _2958_/A vssd1 vssd1 vccd1 vccd1 _2958_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2889_ _2891_/CLK _2889_/D vssd1 vssd1 vccd1 vccd1 _2889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput50 _1775_/Y vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[7] sky130_fd_sc_hd__clkbuf_1
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2743_ _2931_/CLK _2743_/D vssd1 vssd1 vccd1 vccd1 _2743_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2812_ _2815_/CLK _2812_/D vssd1 vssd1 vccd1 vccd1 _2812_/Q sky130_fd_sc_hd__dfxtp_1
X_2674_ _2677_/CLK _2674_/D vssd1 vssd1 vccd1 vccd1 _2674_/Q sky130_fd_sc_hd__dfxtp_1
X_1556_ _2833_/Q _1552_/Y _1555_/Y vssd1 vssd1 vccd1 vccd1 _1764_/B sky130_fd_sc_hd__a21oi_4
X_1625_ _1621_/Y _1622_/X _1624_/X vssd1 vssd1 vccd1 vccd1 _1625_/Y sky130_fd_sc_hd__a21oi_1
X_1487_ _2894_/Q vssd1 vssd1 vccd1 vccd1 _1487_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2039_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2108_ _2750_/Q _2100_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _2108_/X sky130_fd_sc_hd__o21ba_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1410_ _1697_/A vssd1 vssd1 vccd1 vccd1 _2151_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2390_ _2853_/Q _2387_/X _2379_/X vssd1 vssd1 vccd1 vccd1 _2390_/X sky130_fd_sc_hd__o21ba_1
X_1341_ input20/X input2/X _2852_/Q vssd1 vssd1 vccd1 vccd1 _1341_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2726_ _2739_/CLK _2726_/D vssd1 vssd1 vccd1 vccd1 _2726_/Q sky130_fd_sc_hd__dfxtp_1
X_1608_ _2702_/Q _2701_/Q vssd1 vssd1 vccd1 vccd1 _1608_/X sky130_fd_sc_hd__or2b_2
X_1539_ _1524_/X _1526_/X _1539_/S vssd1 vssd1 vccd1 vccd1 _1540_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2657_ _2668_/CLK _2657_/D vssd1 vssd1 vccd1 vccd1 _2657_/Q sky130_fd_sc_hd__dfxtp_1
X_2588_ _2929_/Q _2583_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__o21ba_1
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1890_ _2669_/Q _1886_/X _1887_/X vssd1 vssd1 vccd1 vccd1 _1890_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2511_ _1547_/Y _2090_/X _2510_/X vssd1 vssd1 vccd1 vccd1 _2511_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2373_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2430_/A sky130_fd_sc_hd__clkbuf_2
X_2442_ _1626_/S _2430_/X _2436_/X vssd1 vssd1 vccd1 vccd1 _2442_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1324_ _1320_/X _1321_/X _1322_/X _1323_/X _2841_/Q _2842_/Q vssd1 vssd1 vccd1 vccd1
+ _1613_/B sky130_fd_sc_hd__mux4_2
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2709_ _2721_/CLK _2709_/D vssd1 vssd1 vccd1 vccd1 _2709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1942_ _2688_/Q _1932_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _1942_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1873_ _1899_/A vssd1 vssd1 vccd1 vccd1 _1873_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2356_ _2841_/Q _2353_/X _2345_/X vssd1 vssd1 vccd1 vccd1 _2356_/X sky130_fd_sc_hd__o21ba_1
X_2425_ _2439_/A vssd1 vssd1 vccd1 vccd1 _2425_/X sky130_fd_sc_hd__clkbuf_2
X_2287_ _2814_/Q _2282_/X _2286_/X vssd1 vssd1 vccd1 vccd1 _2815_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2210_ _2788_/Q _2196_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _2210_/X sky130_fd_sc_hd__o21ba_1
X_2072_ _2736_/Q _2068_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _2072_/X sky130_fd_sc_hd__o21ba_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2141_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2141_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1925_ _2721_/Q _1925_/B vssd1 vssd1 vccd1 vccd1 _1926_/A sky130_fd_sc_hd__and2_1
X_1856_ _2658_/Q _1850_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _1856_/X sky130_fd_sc_hd__o21ba_1
X_1787_ _2820_/Q _1794_/B _2821_/Q vssd1 vssd1 vccd1 vccd1 _1787_/X sky130_fd_sc_hd__or3b_1
X_2339_ _2384_/A vssd1 vssd1 vccd1 vccd1 _2339_/X sky130_fd_sc_hd__clkbuf_2
X_2408_ _2859_/Q _2397_/X _2407_/X vssd1 vssd1 vccd1 vccd1 _2860_/D sky130_fd_sc_hd__o21a_1
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2690_ _2907_/CLK _2690_/D vssd1 vssd1 vccd1 vccd1 _2690_/Q sky130_fd_sc_hd__dfxtp_1
X_1641_ _1641_/A _1644_/B vssd1 vssd1 vccd1 vccd1 _1641_/Y sky130_fd_sc_hd__nor2_2
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1710_ _2926_/Q _1572_/B _2927_/Q vssd1 vssd1 vccd1 vccd1 _1713_/B sky130_fd_sc_hd__a21oi_1
X_1572_ _1572_/A _1572_/B vssd1 vssd1 vccd1 vccd1 _1572_/X sky130_fd_sc_hd__and2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _2756_/Q _2113_/X _2114_/X vssd1 vssd1 vccd1 vccd1 _2124_/X sky130_fd_sc_hd__o21ba_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ _2114_/A vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1908_ _2676_/Q _1899_/X _1901_/X vssd1 vssd1 vccd1 vccd1 _1908_/X sky130_fd_sc_hd__o21ba_1
X_1839_ _2651_/Q _1837_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _1839_/X sky130_fd_sc_hd__o21ba_1
X_2888_ _2891_/CLK _2888_/D vssd1 vssd1 vccd1 vccd1 _2888_/Q sky130_fd_sc_hd__dfxtp_1
X_2957_ _2960_/A vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput40 _2959_/A vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[9] sky130_fd_sc_hd__clkbuf_1
Xoutput51 _1772_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_prog_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2742_ _2755_/CLK _2742_/D vssd1 vssd1 vccd1 vccd1 _2742_/Q sky130_fd_sc_hd__dfxtp_1
X_2811_ _2951_/CLK _2811_/D vssd1 vssd1 vccd1 vccd1 _2811_/Q sky130_fd_sc_hd__dfxtp_1
X_2673_ _2677_/CLK _2673_/D vssd1 vssd1 vccd1 vccd1 _2673_/Q sky130_fd_sc_hd__dfxtp_1
X_1555_ _2832_/Q _1553_/X _1554_/X vssd1 vssd1 vccd1 vccd1 _1555_/Y sky130_fd_sc_hd__a21oi_1
X_1624_ _1626_/S _1624_/B _2874_/Q vssd1 vssd1 vccd1 vccd1 _1624_/X sky130_fd_sc_hd__and3b_1
X_1486_ _2681_/Q vssd1 vssd1 vccd1 vccd1 _1486_/Y sky130_fd_sc_hd__inv_2
X_2107_ _2748_/Q _2097_/X _2106_/X vssd1 vssd1 vccd1 vccd1 _2749_/D sky130_fd_sc_hd__o21a_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _2038_/A vssd1 vssd1 vccd1 vccd1 _2724_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_13_prog_clk clkbuf_2_3_0_prog_clk/X vssd1 vssd1 vccd1 vccd1 _2735_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1340_ _2853_/Q vssd1 vssd1 vccd1 vccd1 _1340_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2656_ _2668_/CLK _2656_/D vssd1 vssd1 vccd1 vccd1 _2656_/Q sky130_fd_sc_hd__dfxtp_1
X_2725_ _2739_/CLK _2725_/D vssd1 vssd1 vccd1 vccd1 _2725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1469_ _1476_/A vssd1 vssd1 vccd1 vccd1 _1469_/Y sky130_fd_sc_hd__inv_2
X_1607_ _1540_/Y _1546_/X _1607_/S vssd1 vssd1 vccd1 vccd1 _1867_/D sky130_fd_sc_hd__mux2_1
X_1538_ _1538_/A _1538_/B vssd1 vssd1 vccd1 vccd1 _1539_/S sky130_fd_sc_hd__nand2_1
X_2587_ _2611_/A vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2510_ _2510_/A vssd1 vssd1 vccd1 vccd1 _2510_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1323_ _1322_/S _1624_/B vssd1 vssd1 vccd1 vccd1 _1323_/X sky130_fd_sc_hd__and2b_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2441_ _2871_/Q _2439_/X _2440_/X vssd1 vssd1 vccd1 vccd1 _2872_/D sky130_fd_sc_hd__o21a_1
X_2372_ _2851_/Q _2370_/X _2371_/X vssd1 vssd1 vccd1 vccd1 _2846_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2708_ _2721_/CLK _2708_/D vssd1 vssd1 vccd1 vccd1 _2708_/Q sky130_fd_sc_hd__dfxtp_1
X_2639_ _2639_/A _2639_/B vssd1 vssd1 vccd1 vccd1 _2951_/D sky130_fd_sc_hd__nor2_1
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1941_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1941_/X sky130_fd_sc_hd__clkbuf_2
X_1872_ _2702_/Q _1870_/X _1871_/X vssd1 vssd1 vccd1 vccd1 _2662_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2355_ _2845_/Q _2352_/X _2354_/X vssd1 vssd1 vccd1 vccd1 _2840_/D sky130_fd_sc_hd__o21a_1
X_2424_ _2865_/Q _2412_/X _2423_/X vssd1 vssd1 vccd1 vccd1 _2866_/D sky130_fd_sc_hd__o21a_1
X_2286_ _2815_/Q _2285_/X _2277_/X vssd1 vssd1 vccd1 vccd1 _2286_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2140_ _2212_/A vssd1 vssd1 vccd1 vccd1 _2196_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2071_ _2734_/Q _2066_/X _2070_/X vssd1 vssd1 vccd1 vccd1 _2735_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1924_ _2680_/Q _1910_/X _1923_/Y vssd1 vssd1 vccd1 vccd1 _2681_/D sky130_fd_sc_hd__o21a_1
X_1855_ _2656_/Q _1849_/X _1854_/X vssd1 vssd1 vccd1 vccd1 _2657_/D sky130_fd_sc_hd__o21a_1
X_1786_ _1786_/A _2821_/Q _2820_/Q vssd1 vssd1 vccd1 vccd1 _1786_/X sky130_fd_sc_hd__or3b_1
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2338_ _2839_/Q _2321_/X _2337_/X vssd1 vssd1 vccd1 vccd1 _2834_/D sky130_fd_sc_hd__o21a_1
X_2407_ _2860_/Q _2404_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _2407_/X sky130_fd_sc_hd__o21ba_1
X_2269_ _2269_/A _2951_/Q vssd1 vssd1 vccd1 vccd1 _2314_/S sky130_fd_sc_hd__nand2_1
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_prog_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1640_ _1739_/A _1640_/B vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__nand2_1
X_1571_ _2886_/Q vssd1 vssd1 vccd1 vccd1 _1572_/A sky130_fd_sc_hd__clkbuf_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2123_/X sky130_fd_sc_hd__clkbuf_2
X_2054_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2114_/A sky130_fd_sc_hd__clkbuf_2
X_1907_ _2674_/Q _1896_/X _1906_/X vssd1 vssd1 vccd1 vccd1 _2675_/D sky130_fd_sc_hd__o21a_1
X_1838_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1838_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2887_ _2891_/CLK _2887_/D vssd1 vssd1 vccd1 vccd1 _2887_/Q sky130_fd_sc_hd__dfxtp_2
X_2956_ _2961_/A vssd1 vssd1 vccd1 vccd1 _2956_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1769_ _1769_/A vssd1 vssd1 vccd1 vccd1 _2095_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput30 _2960_/A vssd1 vssd1 vccd1 vccd1 cu_x0y0n_L1[10] sky130_fd_sc_hd__clkbuf_1
Xoutput52 _2959_/X vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_31_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput41 _1782_/Y vssd1 vssd1 vccd1 vccd1 cu_x0y0s_L1[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2672_ _2677_/CLK _2672_/D vssd1 vssd1 vccd1 vccd1 _2672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2741_ _2755_/CLK _2741_/D vssd1 vssd1 vccd1 vccd1 _2741_/Q sky130_fd_sc_hd__dfxtp_1
X_2810_ _2815_/CLK _2810_/D vssd1 vssd1 vccd1 vccd1 _2810_/Q sky130_fd_sc_hd__dfxtp_1
X_1485_ _1485_/A vssd1 vssd1 vccd1 vccd1 _2955_/A sky130_fd_sc_hd__buf_4
X_1554_ _1548_/Y _1553_/S input10/X _2833_/Q vssd1 vssd1 vccd1 vccd1 _1554_/X sky130_fd_sc_hd__a31o_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1623_ _2873_/Q vssd1 vssd1 vccd1 vccd1 _1626_/S sky130_fd_sc_hd__dlymetal6s2s_1
.ends

