// SPDX-FileCopyrightText: 2022 Princeton University
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// Automatically generated by PRGA's RTL generator
module tile_clb (
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif
    output wire [11:0] cu_x0y0n_L1
    , output wire [11:0] cu_x0y0s_L1
    , input wire [11:0] bi_u1y0n_L1
    , input wire [11:0] bi_u1y0s_L1
    , input wire [0:0] clk
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [7:0] _i_blk__out;
    wire [0:0] _i_blk__prog_dout;
    wire [0:0] _i_blk__prog_we_o;
    wire [11:0] _i_cbox_e0__cu_x0y0n_L1;
    wire [11:0] _i_cbox_e0__cu_x0y0s_L1;
    wire [0:0] _i_cbox_e0__prog_dout;
    wire [0:0] _i_cbox_e0__prog_we_o;
    wire [15:0] _i_cbox_w0__bp_x0y0i0_in;
    wire [0:0] _i_cbox_w0__prog_dout;
    wire [0:0] _i_cbox_w0__prog_we_o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_buf_prog_rst_l1__Q;
    wire [0:0] _i_buf_prog_done_l1__Q;
        
    clb i_blk (
        .clk(clk)
        ,.in(_i_cbox_w0__bp_x0y0i0_in)
        ,.out(_i_blk__out)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_blk__prog_dout)
        ,.prog_we_o(_i_blk__prog_we_o)
        );
    cbox_tile_clb_e0 i_cbox_e0 (
        .bp_x0y0i0_out(_i_blk__out)
        ,.cu_x0y0n_L1(_i_cbox_e0__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_cbox_e0__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_blk__prog_we_o)
        ,.prog_din(_i_blk__prog_dout)
        ,.prog_dout(_i_cbox_e0__prog_dout)
        ,.prog_we_o(_i_cbox_e0__prog_we_o)
        );
    cbox_tile_clb_w0 i_cbox_w0 (
        .bp_x0y0i0_in(_i_cbox_w0__bp_x0y0i0_in)
        ,.bi_u1y0n_L1(bi_u1y0n_L1)
        ,.bi_u1y0s_L1(bi_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_cbox_e0__prog_we_o)
        ,.prog_din(_i_cbox_e0__prog_dout)
        ,.prog_dout(_i_cbox_w0__prog_dout)
        ,.prog_we_o(_i_cbox_w0__prog_we_o)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(_i_buf_prog_rst_l1__Q)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(_i_buf_prog_done_l1__Q)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    prga_simple_buf i_buf_prog_rst_l1 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l1__Q)
        );
    prga_simple_bufr i_buf_prog_done_l1 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l1__Q)
        );
        
    assign cu_x0y0n_L1 = _i_cbox_e0__cu_x0y0n_L1;
    assign cu_x0y0s_L1 = _i_cbox_e0__cu_x0y0s_L1;
    assign prog_dout = _i_cbox_w0__prog_dout;
    assign prog_we_o = _i_cbox_w0__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module clb (
    input wire [0:0] clk
    , input wire [15:0] in
    , output wire [7:0] out
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _cluster_i0__o;
    wire [0:0] _cluster_i0__prog_dout;
    wire [0:0] _cluster_i1__o;
    wire [0:0] _cluster_i1__prog_dout;
    wire [0:0] _cluster_i2__o;
    wire [0:0] _cluster_i2__prog_dout;
    wire [0:0] _cluster_i3__o;
    wire [0:0] _cluster_i3__prog_dout;
    wire [0:0] _cluster_i4__o;
    wire [0:0] _cluster_i4__prog_dout;
    wire [0:0] _cluster_i5__o;
    wire [0:0] _cluster_i5__prog_dout;
    wire [0:0] _cluster_i6__o;
    wire [0:0] _cluster_i6__prog_dout;
    wire [0:0] _cluster_i7__o;
    wire [0:0] _cluster_i7__prog_dout;
    wire [0:0] _i_sw_cluster_i0_i_0__o;
    wire [0:0] _i_sw_cluster_i0_i_1__o;
    wire [0:0] _i_sw_cluster_i0_i_2__o;
    wire [0:0] _i_sw_cluster_i0_i_3__o;
    wire [0:0] _i_sw_cluster_i1_i_0__o;
    wire [0:0] _i_sw_cluster_i1_i_1__o;
    wire [0:0] _i_sw_cluster_i1_i_2__o;
    wire [0:0] _i_sw_cluster_i1_i_3__o;
    wire [0:0] _i_sw_cluster_i2_i_0__o;
    wire [0:0] _i_sw_cluster_i2_i_1__o;
    wire [0:0] _i_sw_cluster_i2_i_2__o;
    wire [0:0] _i_sw_cluster_i2_i_3__o;
    wire [0:0] _i_sw_cluster_i3_i_0__o;
    wire [0:0] _i_sw_cluster_i3_i_1__o;
    wire [0:0] _i_sw_cluster_i3_i_2__o;
    wire [0:0] _i_sw_cluster_i3_i_3__o;
    wire [0:0] _i_sw_cluster_i4_i_0__o;
    wire [0:0] _i_sw_cluster_i4_i_1__o;
    wire [0:0] _i_sw_cluster_i4_i_2__o;
    wire [0:0] _i_sw_cluster_i4_i_3__o;
    wire [0:0] _i_sw_cluster_i5_i_0__o;
    wire [0:0] _i_sw_cluster_i5_i_1__o;
    wire [0:0] _i_sw_cluster_i5_i_2__o;
    wire [0:0] _i_sw_cluster_i5_i_3__o;
    wire [0:0] _i_sw_cluster_i6_i_0__o;
    wire [0:0] _i_sw_cluster_i6_i_1__o;
    wire [0:0] _i_sw_cluster_i6_i_2__o;
    wire [0:0] _i_sw_cluster_i6_i_3__o;
    wire [0:0] _i_sw_cluster_i7_i_0__o;
    wire [0:0] _i_sw_cluster_i7_i_1__o;
    wire [0:0] _i_sw_cluster_i7_i_2__o;
    wire [0:0] _i_sw_cluster_i7_i_3__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_cluster_i0_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i0_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i0_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i0_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i0_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i0_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i0_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i0_i_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i1_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i1_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i1_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i1_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i1_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i1_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i1_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i1_i_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i2_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i2_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i2_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i2_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i2_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i2_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i2_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i2_i_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i3_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i3_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i3_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i3_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i3_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i3_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i3_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i3_i_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i4_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i4_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i4_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i4_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i4_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i4_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i4_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i4_i_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i5_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i5_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i5_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i5_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i5_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i5_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i5_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i5_i_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i6_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i6_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i6_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i6_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i6_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i6_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i6_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i6_i_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i7_i_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i7_i_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i7_i_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i7_i_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i7_i_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i7_i_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cluster_i7_i_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cluster_i7_i_3__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    slice cluster_i0 (
        .clk(clk)
        ,.i({_i_sw_cluster_i0_i_3__o,
            _i_sw_cluster_i0_i_2__o,
            _i_sw_cluster_i0_i_1__o,
            _i_sw_cluster_i0_i_0__o})
        ,.o(_cluster_i0__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_cluster_i0__prog_dout)
        );
    slice cluster_i1 (
        .clk(clk)
        ,.i({_i_sw_cluster_i1_i_3__o,
            _i_sw_cluster_i1_i_2__o,
            _i_sw_cluster_i1_i_1__o,
            _i_sw_cluster_i1_i_0__o})
        ,.o(_cluster_i1__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i0__prog_dout)
        ,.prog_dout(_cluster_i1__prog_dout)
        );
    slice cluster_i2 (
        .clk(clk)
        ,.i({_i_sw_cluster_i2_i_3__o,
            _i_sw_cluster_i2_i_2__o,
            _i_sw_cluster_i2_i_1__o,
            _i_sw_cluster_i2_i_0__o})
        ,.o(_cluster_i2__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i1__prog_dout)
        ,.prog_dout(_cluster_i2__prog_dout)
        );
    slice cluster_i3 (
        .clk(clk)
        ,.i({_i_sw_cluster_i3_i_3__o,
            _i_sw_cluster_i3_i_2__o,
            _i_sw_cluster_i3_i_1__o,
            _i_sw_cluster_i3_i_0__o})
        ,.o(_cluster_i3__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i2__prog_dout)
        ,.prog_dout(_cluster_i3__prog_dout)
        );
    slice cluster_i4 (
        .clk(clk)
        ,.i({_i_sw_cluster_i4_i_3__o,
            _i_sw_cluster_i4_i_2__o,
            _i_sw_cluster_i4_i_1__o,
            _i_sw_cluster_i4_i_0__o})
        ,.o(_cluster_i4__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i3__prog_dout)
        ,.prog_dout(_cluster_i4__prog_dout)
        );
    slice cluster_i5 (
        .clk(clk)
        ,.i({_i_sw_cluster_i5_i_3__o,
            _i_sw_cluster_i5_i_2__o,
            _i_sw_cluster_i5_i_1__o,
            _i_sw_cluster_i5_i_0__o})
        ,.o(_cluster_i5__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i4__prog_dout)
        ,.prog_dout(_cluster_i5__prog_dout)
        );
    slice cluster_i6 (
        .clk(clk)
        ,.i({_i_sw_cluster_i6_i_3__o,
            _i_sw_cluster_i6_i_2__o,
            _i_sw_cluster_i6_i_1__o,
            _i_sw_cluster_i6_i_0__o})
        ,.o(_cluster_i6__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i5__prog_dout)
        ,.prog_dout(_cluster_i6__prog_dout)
        );
    slice cluster_i7 (
        .clk(clk)
        ,.i({_i_sw_cluster_i7_i_3__o,
            _i_sw_cluster_i7_i_2__o,
            _i_sw_cluster_i7_i_1__o,
            _i_sw_cluster_i7_i_0__o})
        ,.o(_cluster_i7__o)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i6__prog_dout)
        ,.prog_dout(_cluster_i7__prog_dout)
        );
    sw3 i_sw_cluster_i0_i_0 (
        .i({_cluster_i0__o,
            in[8],
            in[0]})
        ,.o(_i_sw_cluster_i0_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_0__prog_data)
        );
    sw3 i_sw_cluster_i0_i_1 (
        .i({_cluster_i2__o,
            in[10],
            in[2]})
        ,.o(_i_sw_cluster_i0_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_1__prog_data)
        );
    sw3 i_sw_cluster_i0_i_2 (
        .i({_cluster_i4__o,
            in[12],
            in[4]})
        ,.o(_i_sw_cluster_i0_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_2__prog_data)
        );
    sw3 i_sw_cluster_i0_i_3 (
        .i({_cluster_i6__o,
            in[14],
            in[6]})
        ,.o(_i_sw_cluster_i0_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_3__prog_data)
        );
    sw3 i_sw_cluster_i1_i_0 (
        .i({_cluster_i1__o,
            in[9],
            in[1]})
        ,.o(_i_sw_cluster_i1_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_0__prog_data)
        );
    sw3 i_sw_cluster_i1_i_1 (
        .i({_cluster_i4__o,
            in[11],
            in[3]})
        ,.o(_i_sw_cluster_i1_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_1__prog_data)
        );
    sw3 i_sw_cluster_i1_i_2 (
        .i({_cluster_i5__o,
            in[13],
            in[5]})
        ,.o(_i_sw_cluster_i1_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_2__prog_data)
        );
    sw3 i_sw_cluster_i1_i_3 (
        .i({_cluster_i7__o,
            in[15],
            in[8]})
        ,.o(_i_sw_cluster_i1_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_3__prog_data)
        );
    sw3 i_sw_cluster_i2_i_0 (
        .i({_cluster_i0__o,
            in[7],
            in[0]})
        ,.o(_i_sw_cluster_i2_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_0__prog_data)
        );
    sw3 i_sw_cluster_i2_i_1 (
        .i({_cluster_i2__o,
            in[10],
            in[2]})
        ,.o(_i_sw_cluster_i2_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_1__prog_data)
        );
    sw3 i_sw_cluster_i2_i_2 (
        .i({_cluster_i3__o,
            in[12],
            in[4]})
        ,.o(_i_sw_cluster_i2_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_2__prog_data)
        );
    sw3 i_sw_cluster_i2_i_3 (
        .i({_cluster_i4__o,
            in[14],
            in[6]})
        ,.o(_i_sw_cluster_i2_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_3__prog_data)
        );
    sw3 i_sw_cluster_i3_i_0 (
        .i({_cluster_i0__o,
            in[9],
            in[1]})
        ,.o(_i_sw_cluster_i3_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_0__prog_data)
        );
    sw3 i_sw_cluster_i3_i_1 (
        .i({_cluster_i1__o,
            in[11],
            in[3]})
        ,.o(_i_sw_cluster_i3_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_1__prog_data)
        );
    sw3 i_sw_cluster_i3_i_2 (
        .i({_cluster_i5__o,
            in[13],
            in[5]})
        ,.o(_i_sw_cluster_i3_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_2__prog_data)
        );
    sw3 i_sw_cluster_i3_i_3 (
        .i({_cluster_i6__o,
            in[15],
            in[8]})
        ,.o(_i_sw_cluster_i3_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_3__prog_data)
        );
    sw3 i_sw_cluster_i4_i_0 (
        .i({_cluster_i2__o,
            in[7],
            in[0]})
        ,.o(_i_sw_cluster_i4_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_0__prog_data)
        );
    sw3 i_sw_cluster_i4_i_1 (
        .i({_cluster_i3__o,
            in[9],
            in[2]})
        ,.o(_i_sw_cluster_i4_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_1__prog_data)
        );
    sw3 i_sw_cluster_i4_i_2 (
        .i({_cluster_i4__o,
            in[12],
            in[4]})
        ,.o(_i_sw_cluster_i4_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_2__prog_data)
        );
    sw3 i_sw_cluster_i4_i_3 (
        .i({_cluster_i6__o,
            in[14],
            in[6]})
        ,.o(_i_sw_cluster_i4_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_3__prog_data)
        );
    sw3 i_sw_cluster_i5_i_0 (
        .i({_cluster_i2__o,
            in[10],
            in[3]})
        ,.o(_i_sw_cluster_i5_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_0__prog_data)
        );
    sw3 i_sw_cluster_i5_i_1 (
        .i({_cluster_i4__o,
            in[11],
            in[5]})
        ,.o(_i_sw_cluster_i5_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_1__prog_data)
        );
    sw3 i_sw_cluster_i5_i_2 (
        .i({_cluster_i6__o,
            in[13],
            in[6]})
        ,.o(_i_sw_cluster_i5_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_2__prog_data)
        );
    sw3 i_sw_cluster_i5_i_3 (
        .i({_cluster_i7__o,
            in[15],
            in[8]})
        ,.o(_i_sw_cluster_i5_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_3__prog_data)
        );
    sw3 i_sw_cluster_i6_i_0 (
        .i({_cluster_i1__o,
            in[8],
            in[0]})
        ,.o(_i_sw_cluster_i6_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_0__prog_data)
        );
    sw3 i_sw_cluster_i6_i_1 (
        .i({_cluster_i4__o,
            in[10],
            in[1]})
        ,.o(_i_sw_cluster_i6_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_1__prog_data)
        );
    sw3 i_sw_cluster_i6_i_2 (
        .i({_cluster_i5__o,
            in[12],
            in[5]})
        ,.o(_i_sw_cluster_i6_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_2__prog_data)
        );
    sw3 i_sw_cluster_i6_i_3 (
        .i({_cluster_i7__o,
            in[14],
            in[7]})
        ,.o(_i_sw_cluster_i6_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_3__prog_data)
        );
    sw3 i_sw_cluster_i7_i_0 (
        .i({_cluster_i0__o,
            in[7],
            in[0]})
        ,.o(_i_sw_cluster_i7_i_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_0__prog_data)
        );
    sw3 i_sw_cluster_i7_i_1 (
        .i({_cluster_i1__o,
            in[11],
            in[2]})
        ,.o(_i_sw_cluster_i7_i_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_1__prog_data)
        );
    sw3 i_sw_cluster_i7_i_2 (
        .i({_cluster_i2__o,
            in[13],
            in[4]})
        ,.o(_i_sw_cluster_i7_i_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_2__prog_data)
        );
    sw3 i_sw_cluster_i7_i_3 (
        .i({_cluster_i3__o,
            in[15],
            in[5]})
        ,.o(_i_sw_cluster_i7_i_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_3__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i0_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_cluster_i7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i0_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i0_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i0_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i0_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i0_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i0_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i0_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i0_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i0_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i0_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i0_i_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i1_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i0_i_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i1_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i1_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i1_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i1_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i1_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i1_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i1_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i1_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i1_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i1_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i1_i_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i2_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i1_i_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i2_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i2_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i2_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i2_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i2_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i2_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i2_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i2_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i2_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i2_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i2_i_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i3_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i2_i_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i3_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i3_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i3_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i3_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i3_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i3_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i3_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i3_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i3_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i3_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i3_i_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i4_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i3_i_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i4_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i4_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i4_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i4_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i4_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i4_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i4_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i4_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i4_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i4_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i4_i_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i5_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i4_i_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i5_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i5_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i5_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i5_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i5_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i5_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i5_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i5_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i5_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i5_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i5_i_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i6_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i5_i_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i6_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i6_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i6_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i6_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i6_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i6_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i6_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i6_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i6_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i6_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i6_i_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i7_i_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i6_i_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i7_i_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i7_i_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i7_i_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i7_i_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i7_i_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i7_i_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i7_i_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cluster_i7_i_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i7_i_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cluster_i7_i_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cluster_i7_i_3__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cluster_i7_i_3__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign out = {_cluster_i7__o,
        _cluster_i6__o,
        _cluster_i5__o,
        _cluster_i4__o,
        _cluster_i3__o,
        _cluster_i2__o,
        _cluster_i1__o,
        _cluster_i0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module cbox_tile_clb_e0 (
    input wire [7:0] bp_x0y0i0_out
    , output wire [11:0] cu_x0y0n_L1
    , output wire [11:0] cu_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_cu_x0y0n_L1_0__o;
    wire [0:0] _i_sw_cu_x0y0n_L1_2__o;
    wire [0:0] _i_sw_cu_x0y0n_L1_7__o;
    wire [0:0] _i_sw_cu_x0y0n_L1_8__o;
    wire [0:0] _i_sw_cu_x0y0s_L1_0__o;
    wire [0:0] _i_sw_cu_x0y0s_L1_2__o;
    wire [0:0] _i_sw_cu_x0y0s_L1_7__o;
    wire [0:0] _i_sw_cu_x0y0s_L1_8__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0n_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0n_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0n_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0n_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0n_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0n_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0n_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0n_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0s_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0s_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0s_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0s_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0s_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0s_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0s_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0s_L1_8__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_cu_x0y0n_L1_0 (
        .i({bp_x0y0i0_out[7],
            bp_x0y0i0_out[0]})
        ,.o(_i_sw_cu_x0y0n_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_0__prog_data)
        );
    sw2 i_sw_cu_x0y0n_L1_2 (
        .i({bp_x0y0i0_out[6],
            bp_x0y0i0_out[2]})
        ,.o(_i_sw_cu_x0y0n_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_2__prog_data)
        );
    sw2 i_sw_cu_x0y0n_L1_7 (
        .i(bp_x0y0i0_out[7:6])
        ,.o(_i_sw_cu_x0y0n_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_7__prog_data)
        );
    sw2 i_sw_cu_x0y0n_L1_8 (
        .i(bp_x0y0i0_out[5:4])
        ,.o(_i_sw_cu_x0y0n_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_8__prog_data)
        );
    sw2 i_sw_cu_x0y0s_L1_0 (
        .i({bp_x0y0i0_out[7],
            bp_x0y0i0_out[0]})
        ,.o(_i_sw_cu_x0y0s_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_0__prog_data)
        );
    sw2 i_sw_cu_x0y0s_L1_2 (
        .i({bp_x0y0i0_out[6],
            bp_x0y0i0_out[2]})
        ,.o(_i_sw_cu_x0y0s_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_2__prog_data)
        );
    sw2 i_sw_cu_x0y0s_L1_7 (
        .i(bp_x0y0i0_out[7:6])
        ,.o(_i_sw_cu_x0y0s_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_7__prog_data)
        );
    sw2 i_sw_cu_x0y0s_L1_8 (
        .i(bp_x0y0i0_out[5:4])
        ,.o(_i_sw_cu_x0y0s_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_8__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0n_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0n_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0n_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0n_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0n_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0n_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0n_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0n_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0n_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0n_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0n_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0s_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0n_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0s_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0s_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0s_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0s_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0s_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0s_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0s_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0s_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0s_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0s_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_8__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0s_L1_8__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign cu_x0y0n_L1 = {bp_x0y0i0_out[1],
        bp_x0y0i0_out[3:2],
        _i_sw_cu_x0y0n_L1_8__o,
        _i_sw_cu_x0y0n_L1_7__o,
        bp_x0y0i0_out[0],
        bp_x0y0i0_out[3],
        bp_x0y0i0_out[1],
        bp_x0y0i0_out[4],
        _i_sw_cu_x0y0n_L1_2__o,
        bp_x0y0i0_out[5],
        _i_sw_cu_x0y0n_L1_0__o};
    assign cu_x0y0s_L1 = {bp_x0y0i0_out[1],
        bp_x0y0i0_out[3:2],
        _i_sw_cu_x0y0s_L1_8__o,
        _i_sw_cu_x0y0s_L1_7__o,
        bp_x0y0i0_out[0],
        bp_x0y0i0_out[3],
        bp_x0y0i0_out[1],
        bp_x0y0i0_out[4],
        _i_sw_cu_x0y0s_L1_2__o,
        bp_x0y0i0_out[5],
        _i_sw_cu_x0y0s_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module cbox_tile_clb_w0 (
    output wire [15:0] bp_x0y0i0_in
    , input wire [11:0] bi_u1y0n_L1
    , input wire [11:0] bi_u1y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_bp_x0y0i0_in_0__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_1__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_2__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_3__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_4__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_5__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_6__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_7__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_8__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_9__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_10__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_11__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_12__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_13__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_14__o;
    wire [0:0] _i_sw_bp_x0y0i0_in_15__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_0__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_1__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_2__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_3__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_4__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_5__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_6__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_7__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_8__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_9__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_10__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_11__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_11__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_12__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_12__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_13__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_13__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_14__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_14__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_in_15__prog_dout;
    wire [2:0] _i_prog_data_i_sw_bp_x0y0i0_in_15__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw6 i_sw_bp_x0y0i0_in_0 (
        .i({bi_u1y0s_L1[8],
            bi_u1y0n_L1[8],
            bi_u1y0s_L1[4],
            bi_u1y0n_L1[4],
            bi_u1y0s_L1[0],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_bp_x0y0i0_in_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_0__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_1 (
        .i({bi_u1y0s_L1[11],
            bi_u1y0n_L1[11],
            bi_u1y0s_L1[7],
            bi_u1y0n_L1[7],
            bi_u1y0s_L1[3],
            bi_u1y0n_L1[3]})
        ,.o(_i_sw_bp_x0y0i0_in_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_1__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_2 (
        .i({bi_u1y0s_L1[10],
            bi_u1y0n_L1[10],
            bi_u1y0s_L1[6],
            bi_u1y0n_L1[6],
            bi_u1y0s_L1[2],
            bi_u1y0n_L1[2]})
        ,.o(_i_sw_bp_x0y0i0_in_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_2__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_3 (
        .i({bi_u1y0s_L1[9],
            bi_u1y0n_L1[9],
            bi_u1y0s_L1[5],
            bi_u1y0n_L1[5],
            bi_u1y0s_L1[1],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_bp_x0y0i0_in_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_3__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_4 (
        .i({bi_u1y0s_L1[9],
            bi_u1y0n_L1[9],
            bi_u1y0s_L1[4],
            bi_u1y0n_L1[4],
            bi_u1y0s_L1[1],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_bp_x0y0i0_in_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_4__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_5 (
        .i({bi_u1y0s_L1[7],
            bi_u1y0n_L1[7],
            bi_u1y0s_L1[3],
            bi_u1y0n_L1[3],
            bi_u1y0s_L1[0],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_bp_x0y0i0_in_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_5__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_6 (
        .i({bi_u1y0s_L1[11],
            bi_u1y0n_L1[11],
            bi_u1y0s_L1[8],
            bi_u1y0n_L1[8],
            bi_u1y0s_L1[5],
            bi_u1y0n_L1[5]})
        ,.o(_i_sw_bp_x0y0i0_in_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_6__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_7 (
        .i({bi_u1y0s_L1[10],
            bi_u1y0n_L1[10],
            bi_u1y0s_L1[6],
            bi_u1y0n_L1[6],
            bi_u1y0s_L1[2],
            bi_u1y0n_L1[2]})
        ,.o(_i_sw_bp_x0y0i0_in_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_7__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_8 (
        .i({bi_u1y0s_L1[10],
            bi_u1y0n_L1[10],
            bi_u1y0s_L1[5],
            bi_u1y0n_L1[5],
            bi_u1y0s_L1[2],
            bi_u1y0n_L1[2]})
        ,.o(_i_sw_bp_x0y0i0_in_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_8__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_9 (
        .i({bi_u1y0s_L1[9],
            bi_u1y0n_L1[9],
            bi_u1y0s_L1[4],
            bi_u1y0n_L1[4],
            bi_u1y0s_L1[1],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_bp_x0y0i0_in_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_9__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_10 (
        .i({bi_u1y0s_L1[7],
            bi_u1y0n_L1[7],
            bi_u1y0s_L1[3],
            bi_u1y0n_L1[3],
            bi_u1y0s_L1[0],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_bp_x0y0i0_in_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_10__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_11 (
        .i({bi_u1y0s_L1[11],
            bi_u1y0n_L1[11],
            bi_u1y0s_L1[8],
            bi_u1y0n_L1[8],
            bi_u1y0s_L1[5],
            bi_u1y0n_L1[5]})
        ,.o(_i_sw_bp_x0y0i0_in_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_11__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_12 (
        .i({bi_u1y0s_L1[11],
            bi_u1y0n_L1[11],
            bi_u1y0s_L1[6],
            bi_u1y0n_L1[6],
            bi_u1y0s_L1[3],
            bi_u1y0n_L1[3]})
        ,.o(_i_sw_bp_x0y0i0_in_12__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_12__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_13 (
        .i({bi_u1y0s_L1[9],
            bi_u1y0n_L1[9],
            bi_u1y0s_L1[6],
            bi_u1y0n_L1[6],
            bi_u1y0s_L1[1],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_bp_x0y0i0_in_13__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_13__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_14 (
        .i({bi_u1y0s_L1[4],
            bi_u1y0n_L1[4],
            bi_u1y0s_L1[2],
            bi_u1y0n_L1[2],
            bi_u1y0s_L1[0],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_bp_x0y0i0_in_14__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_14__prog_data)
        );
    sw6 i_sw_bp_x0y0i0_in_15 (
        .i({bi_u1y0s_L1[10],
            bi_u1y0n_L1[10],
            bi_u1y0s_L1[8],
            bi_u1y0n_L1[8],
            bi_u1y0s_L1[7],
            bi_u1y0n_L1[7]})
        ,.o(_i_sw_bp_x0y0i0_in_15__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_15__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_0__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_1__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_2__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_3__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_4__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_5__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_6__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_7__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_8__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_9__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_10__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_11__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_12 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_11__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_12__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_12__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_13 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_12__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_13__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_13__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_14 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_13__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_14__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_14__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_bp_x0y0i0_in_15 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_14__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_in_15__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_in_15__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_in_15__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign bp_x0y0i0_in = {_i_sw_bp_x0y0i0_in_15__o,
        _i_sw_bp_x0y0i0_in_14__o,
        _i_sw_bp_x0y0i0_in_13__o,
        _i_sw_bp_x0y0i0_in_12__o,
        _i_sw_bp_x0y0i0_in_11__o,
        _i_sw_bp_x0y0i0_in_10__o,
        _i_sw_bp_x0y0i0_in_9__o,
        _i_sw_bp_x0y0i0_in_8__o,
        _i_sw_bp_x0y0i0_in_7__o,
        _i_sw_bp_x0y0i0_in_6__o,
        _i_sw_bp_x0y0i0_in_5__o,
        _i_sw_bp_x0y0i0_in_4__o,
        _i_sw_bp_x0y0i0_in_3__o,
        _i_sw_bp_x0y0i0_in_2__o,
        _i_sw_bp_x0y0i0_in_1__o,
        _i_sw_bp_x0y0i0_in_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module prga_simple_buf (
    input wire [0:0] C,
    input wire [0:0] D,
    output reg [0:0] Q
    );

    always @(posedge C) begin
        Q <= D;
    end

endmodule// Automatically generated by PRGA's RTL generator
module prga_simple_bufr (
    input wire [0:0] C,
    input wire [0:0] R,
    input wire [0:0] D,
    output reg [0:0] Q
    );

    always @(posedge C) begin
        if (R) begin
            Q <= 1'b0;
        end else begin
            Q <= D;
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module slice (
    input wire [0:0] clk
    , input wire [3:0] i
    , output wire [0:0] o
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    );
    
        
    wire [0:0] _lut__out;
    wire [0:0] _ff__Q;
    wire [0:0] _i_sw_o__o;
    wire [0:0] _i_prog_data_lut__prog_dout;
    wire [16:0] _i_prog_data_lut__prog_data;
    wire [0:0] _i_prog_data_ff__prog_dout;
    wire [0:0] _i_prog_data_ff__prog_data;
    wire [0:0] _i_prog_data_i_sw_o__prog_dout;
    wire [1:0] _i_prog_data_i_sw_o__prog_data;
        
    lut4 lut (
        .in(i)
        ,.out(_lut__out)
        ,.prog_done(prog_done)
        ,.prog_data(_i_prog_data_lut__prog_data)
        );
    flipflop ff (
        .clk(clk)
        ,.D(_lut__out)
        ,.Q(_ff__Q)
        ,.prog_done(prog_done)
        ,.prog_data(_i_prog_data_ff__prog_data)
        );
    sw2 i_sw_o (
        .i({_ff__Q,
            _lut__out})
        ,.o(_i_sw_o__o)
        ,.prog_done(prog_done)
        ,.prog_data(_i_prog_data_i_sw_o__prog_data)
        );
    scanchain_data_d17 i_prog_data_lut (
        .prog_clk(prog_clk)
        ,.prog_rst(prog_rst)
        ,.prog_done(prog_done)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_prog_data_lut__prog_dout)
        ,.prog_data(_i_prog_data_lut__prog_data)
        );
    scanchain_data_d1 i_prog_data_ff (
        .prog_clk(prog_clk)
        ,.prog_rst(prog_rst)
        ,.prog_done(prog_done)
        ,.prog_we(prog_we)
        ,.prog_din(_i_prog_data_lut__prog_dout)
        ,.prog_dout(_i_prog_data_ff__prog_dout)
        ,.prog_data(_i_prog_data_ff__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_o (
        .prog_clk(prog_clk)
        ,.prog_rst(prog_rst)
        ,.prog_done(prog_done)
        ,.prog_we(prog_we)
        ,.prog_din(_i_prog_data_ff__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_o__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_o__prog_data)
        );
        
    assign o = _i_sw_o__o;
    assign prog_dout = _i_prog_data_i_sw_o__prog_dout;

endmodule
// Automatically generated by PRGA's RTL generator
module sw3 (
    input wire [2:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [1:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                2'd1: o = i[0];
                2'd2: o = i[1];
                2'd3: o = i[2];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_delim (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [0:0] prog_we_o
    , output reg [1 - 1:0] prog_dout
    );

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_we_o <= 1'b0;
            prog_dout <= 1'b0;
        end else if (~prog_done && prog_we) begin
            prog_we_o <= 1'b1;
            prog_dout <= prog_din;
        end else begin
            prog_we_o <= 1'b0;
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d2 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [2 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 2;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule// Automatically generated by PRGA's RTL generator
module sw2 (
    input wire [1:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [1:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                2'd1: o = i[0];
                2'd2: o = i[1];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module sw6 (
    input wire [5:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [2:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                3'd1: o = i[0];
                3'd2: o = i[1];
                3'd3: o = i[2];
                3'd4: o = i[3];
                3'd5: o = i[4];
                3'd6: o = i[5];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d3 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [3 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 3;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule// Automatically generated by PRGA's RTL generator
module lut4 (
    input wire [3:0] in
    , output reg [0:0] out

    , input wire [0:0] prog_done
    , input wire [16:0] prog_data
        // prog_data[ 0 +: 15]: LUT content
        // prog_data[16]: LUT enabled (not disabled)
    );

    localparam  IDX_LUT_ENABLE = 16;

    always @* begin
        if (~prog_done || ~prog_data[IDX_LUT_ENABLE]) begin
            out = 1'b0;
        end else begin
            case (in)
                4'd0: out = prog_data[0];
                4'd1: out = prog_data[1];
                4'd2: out = prog_data[2];
                4'd3: out = prog_data[3];
                4'd4: out = prog_data[4];
                4'd5: out = prog_data[5];
                4'd6: out = prog_data[6];
                4'd7: out = prog_data[7];
                4'd8: out = prog_data[8];
                4'd9: out = prog_data[9];
                4'd10: out = prog_data[10];
                4'd11: out = prog_data[11];
                4'd12: out = prog_data[12];
                4'd13: out = prog_data[13];
                4'd14: out = prog_data[14];
                4'd15: out = prog_data[15];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module flipflop (
    input wire [0:0] clk
    , input wire [0:0] D
    , output reg [0:0] Q

    , input wire [0:0] prog_done    // programming finished
    , input wire [0:0] prog_data    // mode: enabled (not disabled)
    );

    always @(posedge clk) begin
        if (~prog_done || ~prog_data) begin
            Q <= 1'b0;
        end else begin
            Q <= D;
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d17 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [17 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 17;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d1 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [1 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 1;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule
