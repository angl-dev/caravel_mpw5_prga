// SPDX-FileCopyrightText: 2022 Princeton University
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// Automatically generated by PRGA's RTL generator
module top (
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif
    input wire [0:0] ipin_x0y1_0
    , output wire [0:0] opin_x0y1_0
    , output wire [0:0] oe_x0y1_0
    , input wire [0:0] ipin_x0y1_1
    , output wire [0:0] opin_x0y1_1
    , output wire [0:0] oe_x0y1_1
    , input wire [0:0] ipin_x0y2_0
    , output wire [0:0] opin_x0y2_0
    , output wire [0:0] oe_x0y2_0
    , input wire [0:0] ipin_x0y2_1
    , output wire [0:0] opin_x0y2_1
    , output wire [0:0] oe_x0y2_1
    , input wire [0:0] ipin_x0y3_0
    , output wire [0:0] opin_x0y3_0
    , output wire [0:0] oe_x0y3_0
    , input wire [0:0] ipin_x0y3_1
    , output wire [0:0] opin_x0y3_1
    , output wire [0:0] oe_x0y3_1
    , input wire [0:0] ipin_x0y4_0
    , output wire [0:0] opin_x0y4_0
    , output wire [0:0] oe_x0y4_0
    , input wire [0:0] ipin_x0y4_1
    , output wire [0:0] opin_x0y4_1
    , output wire [0:0] oe_x0y4_1
    , input wire [0:0] ipin_x0y5_0
    , output wire [0:0] opin_x0y5_0
    , output wire [0:0] oe_x0y5_0
    , input wire [0:0] ipin_x0y5_1
    , output wire [0:0] opin_x0y5_1
    , output wire [0:0] oe_x0y5_1
    , input wire [0:0] ipin_x0y6_0
    , output wire [0:0] opin_x0y6_0
    , output wire [0:0] oe_x0y6_0
    , input wire [0:0] ipin_x0y6_1
    , output wire [0:0] opin_x0y6_1
    , output wire [0:0] oe_x0y6_1
    , input wire [0:0] ipin_x0y7_0
    , output wire [0:0] opin_x0y7_0
    , output wire [0:0] oe_x0y7_0
    , input wire [0:0] ipin_x0y7_1
    , output wire [0:0] opin_x0y7_1
    , output wire [0:0] oe_x0y7_1
    , input wire [0:0] ipin_x0y8_0
    , output wire [0:0] opin_x0y8_0
    , output wire [0:0] oe_x0y8_0
    , input wire [0:0] ipin_x0y8_1
    , output wire [0:0] opin_x0y8_1
    , output wire [0:0] oe_x0y8_1
    , input wire [0:0] ipin_x1y9_0
    , output wire [0:0] opin_x1y9_0
    , output wire [0:0] oe_x1y9_0
    , input wire [0:0] ipin_x1y9_1
    , output wire [0:0] opin_x1y9_1
    , output wire [0:0] oe_x1y9_1
    , input wire [0:0] ipin_x2y9_0
    , output wire [0:0] opin_x2y9_0
    , output wire [0:0] oe_x2y9_0
    , input wire [0:0] ipin_x2y9_1
    , output wire [0:0] opin_x2y9_1
    , output wire [0:0] oe_x2y9_1
    , input wire [0:0] ipin_x3y9_0
    , output wire [0:0] opin_x3y9_0
    , output wire [0:0] oe_x3y9_0
    , input wire [0:0] ipin_x3y9_1
    , output wire [0:0] opin_x3y9_1
    , output wire [0:0] oe_x3y9_1
    , input wire [0:0] ipin_x4y9_0
    , output wire [0:0] opin_x4y9_0
    , output wire [0:0] oe_x4y9_0
    , input wire [0:0] ipin_x4y9_1
    , output wire [0:0] opin_x4y9_1
    , output wire [0:0] oe_x4y9_1
    , input wire [0:0] ipin_x5y9_0
    , output wire [0:0] opin_x5y9_0
    , output wire [0:0] oe_x5y9_0
    , input wire [0:0] ipin_x5y9_1
    , output wire [0:0] opin_x5y9_1
    , output wire [0:0] oe_x5y9_1
    , input wire [0:0] ipin_x6y9_0
    , output wire [0:0] opin_x6y9_0
    , output wire [0:0] oe_x6y9_0
    , input wire [0:0] ipin_x6y9_1
    , output wire [0:0] opin_x6y9_1
    , output wire [0:0] oe_x6y9_1
    , input wire [0:0] ipin_x7y9_0
    , output wire [0:0] opin_x7y9_0
    , output wire [0:0] oe_x7y9_0
    , input wire [0:0] ipin_x7y9_1
    , output wire [0:0] opin_x7y9_1
    , output wire [0:0] oe_x7y9_1
    , input wire [0:0] ipin_x8y9_0
    , output wire [0:0] opin_x8y9_0
    , output wire [0:0] oe_x8y9_0
    , input wire [0:0] ipin_x8y9_1
    , output wire [0:0] opin_x8y9_1
    , output wire [0:0] oe_x8y9_1
    , input wire [0:0] ipin_x9y1_0
    , output wire [0:0] opin_x9y1_0
    , output wire [0:0] oe_x9y1_0
    , input wire [0:0] ipin_x9y1_1
    , output wire [0:0] opin_x9y1_1
    , output wire [0:0] oe_x9y1_1
    , input wire [0:0] ipin_x9y2_0
    , output wire [0:0] opin_x9y2_0
    , output wire [0:0] oe_x9y2_0
    , input wire [0:0] ipin_x9y2_1
    , output wire [0:0] opin_x9y2_1
    , output wire [0:0] oe_x9y2_1
    , input wire [0:0] ipin_x9y3_0
    , output wire [0:0] opin_x9y3_0
    , output wire [0:0] oe_x9y3_0
    , input wire [0:0] ipin_x9y3_1
    , output wire [0:0] opin_x9y3_1
    , output wire [0:0] oe_x9y3_1
    , input wire [0:0] ipin_x9y4_0
    , output wire [0:0] opin_x9y4_0
    , output wire [0:0] oe_x9y4_0
    , input wire [0:0] ipin_x9y4_1
    , output wire [0:0] opin_x9y4_1
    , output wire [0:0] oe_x9y4_1
    , input wire [0:0] ipin_x9y5_0
    , output wire [0:0] opin_x9y5_0
    , output wire [0:0] oe_x9y5_0
    , input wire [0:0] ipin_x9y5_1
    , output wire [0:0] opin_x9y5_1
    , output wire [0:0] oe_x9y5_1
    , input wire [0:0] ipin_x9y6_0
    , output wire [0:0] opin_x9y6_0
    , output wire [0:0] oe_x9y6_0
    , input wire [0:0] ipin_x9y6_1
    , output wire [0:0] opin_x9y6_1
    , output wire [0:0] oe_x9y6_1
    , input wire [0:0] ipin_x9y7_0
    , output wire [0:0] opin_x9y7_0
    , output wire [0:0] oe_x9y7_0
    , input wire [0:0] ipin_x9y7_1
    , output wire [0:0] opin_x9y7_1
    , output wire [0:0] oe_x9y7_1
    , input wire [0:0] ipin_x9y8_0
    , output wire [0:0] opin_x9y8_0
    , output wire [0:0] oe_x9y8_0
    , input wire [0:0] ipin_x9y8_1
    , output wire [0:0] opin_x9y8_1
    , output wire [0:0] oe_x9y8_1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
endmodule
