VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2750.000 BY 3400.000 ;
  PIN ipin_x0y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END ipin_x0y1_0
  PIN ipin_x0y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END ipin_x0y1_1
  PIN ipin_x0y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END ipin_x0y2_0
  PIN ipin_x0y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END ipin_x0y2_1
  PIN ipin_x0y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END ipin_x0y3_0
  PIN ipin_x0y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END ipin_x0y3_1
  PIN ipin_x0y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END ipin_x0y4_0
  PIN ipin_x0y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END ipin_x0y4_1
  PIN ipin_x0y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END ipin_x0y5_0
  PIN ipin_x0y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END ipin_x0y5_1
  PIN ipin_x0y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END ipin_x0y6_0
  PIN ipin_x0y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.000 4.000 814.600 ;
    END
  END ipin_x0y6_1
  PIN ipin_x0y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.400 4.000 886.000 ;
    END
  END ipin_x0y7_0
  PIN ipin_x0y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.120 4.000 956.720 ;
    END
  END ipin_x0y7_1
  PIN ipin_x0y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END ipin_x0y8_0
  PIN ipin_x0y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1097.560 4.000 1098.160 ;
    END
  END ipin_x0y8_1
  PIN ipin_x1y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 3396.000 28.890 3400.000 ;
    END
  END ipin_x1y9_0
  PIN ipin_x1y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 3396.000 85.930 3400.000 ;
    END
  END ipin_x1y9_1
  PIN ipin_x2y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 3396.000 143.430 3400.000 ;
    END
  END ipin_x2y9_0
  PIN ipin_x2y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 3396.000 200.470 3400.000 ;
    END
  END ipin_x2y9_1
  PIN ipin_x3y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 3396.000 257.970 3400.000 ;
    END
  END ipin_x3y9_0
  PIN ipin_x3y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 3396.000 315.010 3400.000 ;
    END
  END ipin_x3y9_1
  PIN ipin_x4y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 3396.000 372.510 3400.000 ;
    END
  END ipin_x4y9_0
  PIN ipin_x4y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 3396.000 429.550 3400.000 ;
    END
  END ipin_x4y9_1
  PIN ipin_x5y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 3396.000 487.050 3400.000 ;
    END
  END ipin_x5y9_0
  PIN ipin_x5y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 3396.000 544.090 3400.000 ;
    END
  END ipin_x5y9_1
  PIN ipin_x6y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 3396.000 601.590 3400.000 ;
    END
  END ipin_x6y9_0
  PIN ipin_x6y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 3396.000 658.630 3400.000 ;
    END
  END ipin_x6y9_1
  PIN ipin_x7y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 3396.000 716.130 3400.000 ;
    END
  END ipin_x7y9_0
  PIN ipin_x7y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 3396.000 773.630 3400.000 ;
    END
  END ipin_x7y9_1
  PIN ipin_x8y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 3396.000 830.670 3400.000 ;
    END
  END ipin_x8y9_0
  PIN ipin_x8y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 3396.000 888.170 3400.000 ;
    END
  END ipin_x8y9_1
  PIN ipin_x9y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 35.400 2750.000 36.000 ;
    END
  END ipin_x9y1_0
  PIN ipin_x9y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 106.120 2750.000 106.720 ;
    END
  END ipin_x9y1_1
  PIN ipin_x9y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 176.840 2750.000 177.440 ;
    END
  END ipin_x9y2_0
  PIN ipin_x9y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 247.560 2750.000 248.160 ;
    END
  END ipin_x9y2_1
  PIN ipin_x9y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 318.280 2750.000 318.880 ;
    END
  END ipin_x9y3_0
  PIN ipin_x9y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 389.000 2750.000 389.600 ;
    END
  END ipin_x9y3_1
  PIN ipin_x9y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 460.400 2750.000 461.000 ;
    END
  END ipin_x9y4_0
  PIN ipin_x9y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 531.120 2750.000 531.720 ;
    END
  END ipin_x9y4_1
  PIN ipin_x9y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 601.840 2750.000 602.440 ;
    END
  END ipin_x9y5_0
  PIN ipin_x9y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 672.560 2750.000 673.160 ;
    END
  END ipin_x9y5_1
  PIN ipin_x9y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 743.280 2750.000 743.880 ;
    END
  END ipin_x9y6_0
  PIN ipin_x9y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 814.000 2750.000 814.600 ;
    END
  END ipin_x9y6_1
  PIN ipin_x9y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 885.400 2750.000 886.000 ;
    END
  END ipin_x9y7_0
  PIN ipin_x9y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 956.120 2750.000 956.720 ;
    END
  END ipin_x9y7_1
  PIN ipin_x9y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1026.840 2750.000 1027.440 ;
    END
  END ipin_x9y8_0
  PIN ipin_x9y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1097.560 2750.000 1098.160 ;
    END
  END ipin_x9y8_1
  PIN oe_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2301.840 4.000 2302.440 ;
    END
  END oe_x0y1_0
  PIN oe_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2372.560 4.000 2373.160 ;
    END
  END oe_x0y1_1
  PIN oe_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2443.280 4.000 2443.880 ;
    END
  END oe_x0y2_0
  PIN oe_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2514.000 4.000 2514.600 ;
    END
  END oe_x0y2_1
  PIN oe_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2585.400 4.000 2586.000 ;
    END
  END oe_x0y3_0
  PIN oe_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2656.120 4.000 2656.720 ;
    END
  END oe_x0y3_1
  PIN oe_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2726.840 4.000 2727.440 ;
    END
  END oe_x0y4_0
  PIN oe_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2797.560 4.000 2798.160 ;
    END
  END oe_x0y4_1
  PIN oe_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2868.280 4.000 2868.880 ;
    END
  END oe_x0y5_0
  PIN oe_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2939.000 4.000 2939.600 ;
    END
  END oe_x0y5_1
  PIN oe_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3010.400 4.000 3011.000 ;
    END
  END oe_x0y6_0
  PIN oe_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3081.120 4.000 3081.720 ;
    END
  END oe_x0y6_1
  PIN oe_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3151.840 4.000 3152.440 ;
    END
  END oe_x0y7_0
  PIN oe_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3222.560 4.000 3223.160 ;
    END
  END oe_x0y7_1
  PIN oe_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3293.280 4.000 3293.880 ;
    END
  END oe_x0y8_0
  PIN oe_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3364.000 4.000 3364.600 ;
    END
  END oe_x0y8_1
  PIN oe_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 3396.000 1861.990 3400.000 ;
    END
  END oe_x1y9_0
  PIN oe_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.750 3396.000 1919.030 3400.000 ;
    END
  END oe_x1y9_1
  PIN oe_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.250 3396.000 1976.530 3400.000 ;
    END
  END oe_x2y9_0
  PIN oe_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.290 3396.000 2033.570 3400.000 ;
    END
  END oe_x2y9_1
  PIN oe_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.790 3396.000 2091.070 3400.000 ;
    END
  END oe_x3y9_0
  PIN oe_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.290 3396.000 2148.570 3400.000 ;
    END
  END oe_x3y9_1
  PIN oe_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.330 3396.000 2205.610 3400.000 ;
    END
  END oe_x4y9_0
  PIN oe_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.830 3396.000 2263.110 3400.000 ;
    END
  END oe_x4y9_1
  PIN oe_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.870 3396.000 2320.150 3400.000 ;
    END
  END oe_x5y9_0
  PIN oe_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2377.370 3396.000 2377.650 3400.000 ;
    END
  END oe_x5y9_1
  PIN oe_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.410 3396.000 2434.690 3400.000 ;
    END
  END oe_x6y9_0
  PIN oe_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.910 3396.000 2492.190 3400.000 ;
    END
  END oe_x6y9_1
  PIN oe_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2548.950 3396.000 2549.230 3400.000 ;
    END
  END oe_x7y9_0
  PIN oe_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2606.450 3396.000 2606.730 3400.000 ;
    END
  END oe_x7y9_1
  PIN oe_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2663.490 3396.000 2663.770 3400.000 ;
    END
  END oe_x8y9_0
  PIN oe_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.990 3396.000 2721.270 3400.000 ;
    END
  END oe_x8y9_1
  PIN oe_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2301.840 2750.000 2302.440 ;
    END
  END oe_x9y1_0
  PIN oe_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2372.560 2750.000 2373.160 ;
    END
  END oe_x9y1_1
  PIN oe_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2443.280 2750.000 2443.880 ;
    END
  END oe_x9y2_0
  PIN oe_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2514.000 2750.000 2514.600 ;
    END
  END oe_x9y2_1
  PIN oe_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2585.400 2750.000 2586.000 ;
    END
  END oe_x9y3_0
  PIN oe_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2656.120 2750.000 2656.720 ;
    END
  END oe_x9y3_1
  PIN oe_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2726.840 2750.000 2727.440 ;
    END
  END oe_x9y4_0
  PIN oe_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2797.560 2750.000 2798.160 ;
    END
  END oe_x9y4_1
  PIN oe_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2868.280 2750.000 2868.880 ;
    END
  END oe_x9y5_0
  PIN oe_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2939.000 2750.000 2939.600 ;
    END
  END oe_x9y5_1
  PIN oe_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3010.400 2750.000 3011.000 ;
    END
  END oe_x9y6_0
  PIN oe_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3081.120 2750.000 3081.720 ;
    END
  END oe_x9y6_1
  PIN oe_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3151.840 2750.000 3152.440 ;
    END
  END oe_x9y7_0
  PIN oe_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3222.560 2750.000 3223.160 ;
    END
  END oe_x9y7_1
  PIN oe_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3293.280 2750.000 3293.880 ;
    END
  END oe_x9y8_0
  PIN oe_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3364.000 2750.000 3364.600 ;
    END
  END oe_x9y8_1
  PIN opin_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END opin_x0y1_0
  PIN opin_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.000 4.000 1239.600 ;
    END
  END opin_x0y1_1
  PIN opin_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1310.400 4.000 1311.000 ;
    END
  END opin_x0y2_0
  PIN opin_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.120 4.000 1381.720 ;
    END
  END opin_x0y2_1
  PIN opin_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END opin_x0y3_0
  PIN opin_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1522.560 4.000 1523.160 ;
    END
  END opin_x0y3_1
  PIN opin_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1593.280 4.000 1593.880 ;
    END
  END opin_x0y4_0
  PIN opin_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1664.000 4.000 1664.600 ;
    END
  END opin_x0y4_1
  PIN opin_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1735.400 4.000 1736.000 ;
    END
  END opin_x0y5_0
  PIN opin_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1806.120 4.000 1806.720 ;
    END
  END opin_x0y5_1
  PIN opin_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1876.840 4.000 1877.440 ;
    END
  END opin_x0y6_0
  PIN opin_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1947.560 4.000 1948.160 ;
    END
  END opin_x0y6_1
  PIN opin_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2018.280 4.000 2018.880 ;
    END
  END opin_x0y7_0
  PIN opin_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2089.000 4.000 2089.600 ;
    END
  END opin_x0y7_1
  PIN opin_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2160.400 4.000 2161.000 ;
    END
  END opin_x0y8_0
  PIN opin_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2231.120 4.000 2231.720 ;
    END
  END opin_x0y8_1
  PIN opin_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 3396.000 945.210 3400.000 ;
    END
  END opin_x1y9_0
  PIN opin_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 3396.000 1002.710 3400.000 ;
    END
  END opin_x1y9_1
  PIN opin_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 3396.000 1059.750 3400.000 ;
    END
  END opin_x2y9_0
  PIN opin_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 3396.000 1117.250 3400.000 ;
    END
  END opin_x2y9_1
  PIN opin_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 3396.000 1174.290 3400.000 ;
    END
  END opin_x3y9_0
  PIN opin_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.510 3396.000 1231.790 3400.000 ;
    END
  END opin_x3y9_1
  PIN opin_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.550 3396.000 1288.830 3400.000 ;
    END
  END opin_x4y9_0
  PIN opin_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 3396.000 1346.330 3400.000 ;
    END
  END opin_x4y9_1
  PIN opin_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.550 3396.000 1403.830 3400.000 ;
    END
  END opin_x5y9_0
  PIN opin_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.590 3396.000 1460.870 3400.000 ;
    END
  END opin_x5y9_1
  PIN opin_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 3396.000 1518.370 3400.000 ;
    END
  END opin_x6y9_0
  PIN opin_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 3396.000 1575.410 3400.000 ;
    END
  END opin_x6y9_1
  PIN opin_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 3396.000 1632.910 3400.000 ;
    END
  END opin_x7y9_0
  PIN opin_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 3396.000 1689.950 3400.000 ;
    END
  END opin_x7y9_1
  PIN opin_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 3396.000 1747.450 3400.000 ;
    END
  END opin_x8y9_0
  PIN opin_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.210 3396.000 1804.490 3400.000 ;
    END
  END opin_x8y9_1
  PIN opin_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1168.280 2750.000 1168.880 ;
    END
  END opin_x9y1_0
  PIN opin_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1239.000 2750.000 1239.600 ;
    END
  END opin_x9y1_1
  PIN opin_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1310.400 2750.000 1311.000 ;
    END
  END opin_x9y2_0
  PIN opin_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1381.120 2750.000 1381.720 ;
    END
  END opin_x9y2_1
  PIN opin_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1451.840 2750.000 1452.440 ;
    END
  END opin_x9y3_0
  PIN opin_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1522.560 2750.000 1523.160 ;
    END
  END opin_x9y3_1
  PIN opin_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1593.280 2750.000 1593.880 ;
    END
  END opin_x9y4_0
  PIN opin_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1664.000 2750.000 1664.600 ;
    END
  END opin_x9y4_1
  PIN opin_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1735.400 2750.000 1736.000 ;
    END
  END opin_x9y5_0
  PIN opin_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1806.120 2750.000 1806.720 ;
    END
  END opin_x9y5_1
  PIN opin_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1876.840 2750.000 1877.440 ;
    END
  END opin_x9y6_0
  PIN opin_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1947.560 2750.000 1948.160 ;
    END
  END opin_x9y6_1
  PIN opin_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2018.280 2750.000 2018.880 ;
    END
  END opin_x9y7_0
  PIN opin_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2089.000 2750.000 2089.600 ;
    END
  END opin_x9y7_1
  PIN opin_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2160.400 2750.000 2161.000 ;
    END
  END opin_x9y8_0
  PIN opin_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2231.120 2750.000 2231.720 ;
    END
  END opin_x9y8_1
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END prog_clk
  PIN prog_din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END prog_din
  PIN prog_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END prog_done
  PIN prog_dout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END prog_dout
  PIN prog_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 0.000 1768.150 4.000 ;
    END
  END prog_rst
  PIN prog_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.710 0.000 2160.990 4.000 ;
    END
  END prog_we
  PIN prog_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2553.550 0.000 2553.830 4.000 ;
    END
  END prog_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 3389.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 3389.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 3389.360 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2744.360 3389.205 ;
      LAYER met1 ;
        RECT 5.520 10.640 2744.360 3389.360 ;
      LAYER met2 ;
        RECT 6.990 3395.720 28.330 3396.330 ;
        RECT 29.170 3395.720 85.370 3396.330 ;
        RECT 86.210 3395.720 142.870 3396.330 ;
        RECT 143.710 3395.720 199.910 3396.330 ;
        RECT 200.750 3395.720 257.410 3396.330 ;
        RECT 258.250 3395.720 314.450 3396.330 ;
        RECT 315.290 3395.720 371.950 3396.330 ;
        RECT 372.790 3395.720 428.990 3396.330 ;
        RECT 429.830 3395.720 486.490 3396.330 ;
        RECT 487.330 3395.720 543.530 3396.330 ;
        RECT 544.370 3395.720 601.030 3396.330 ;
        RECT 601.870 3395.720 658.070 3396.330 ;
        RECT 658.910 3395.720 715.570 3396.330 ;
        RECT 716.410 3395.720 773.070 3396.330 ;
        RECT 773.910 3395.720 830.110 3396.330 ;
        RECT 830.950 3395.720 887.610 3396.330 ;
        RECT 888.450 3395.720 944.650 3396.330 ;
        RECT 945.490 3395.720 1002.150 3396.330 ;
        RECT 1002.990 3395.720 1059.190 3396.330 ;
        RECT 1060.030 3395.720 1116.690 3396.330 ;
        RECT 1117.530 3395.720 1173.730 3396.330 ;
        RECT 1174.570 3395.720 1231.230 3396.330 ;
        RECT 1232.070 3395.720 1288.270 3396.330 ;
        RECT 1289.110 3395.720 1345.770 3396.330 ;
        RECT 1346.610 3395.720 1403.270 3396.330 ;
        RECT 1404.110 3395.720 1460.310 3396.330 ;
        RECT 1461.150 3395.720 1517.810 3396.330 ;
        RECT 1518.650 3395.720 1574.850 3396.330 ;
        RECT 1575.690 3395.720 1632.350 3396.330 ;
        RECT 1633.190 3395.720 1689.390 3396.330 ;
        RECT 1690.230 3395.720 1746.890 3396.330 ;
        RECT 1747.730 3395.720 1803.930 3396.330 ;
        RECT 1804.770 3395.720 1861.430 3396.330 ;
        RECT 1862.270 3395.720 1918.470 3396.330 ;
        RECT 1919.310 3395.720 1975.970 3396.330 ;
        RECT 1976.810 3395.720 2033.010 3396.330 ;
        RECT 2033.850 3395.720 2090.510 3396.330 ;
        RECT 2091.350 3395.720 2148.010 3396.330 ;
        RECT 2148.850 3395.720 2205.050 3396.330 ;
        RECT 2205.890 3395.720 2262.550 3396.330 ;
        RECT 2263.390 3395.720 2319.590 3396.330 ;
        RECT 2320.430 3395.720 2377.090 3396.330 ;
        RECT 2377.930 3395.720 2434.130 3396.330 ;
        RECT 2434.970 3395.720 2491.630 3396.330 ;
        RECT 2492.470 3395.720 2548.670 3396.330 ;
        RECT 2549.510 3395.720 2606.170 3396.330 ;
        RECT 2607.010 3395.720 2663.210 3396.330 ;
        RECT 2664.050 3395.720 2720.710 3396.330 ;
        RECT 2721.550 3395.720 2741.050 3396.330 ;
        RECT 6.990 4.280 2741.050 3395.720 ;
        RECT 6.990 4.000 196.230 4.280 ;
        RECT 197.070 4.000 589.070 4.280 ;
        RECT 589.910 4.000 981.910 4.280 ;
        RECT 982.750 4.000 1374.750 4.280 ;
        RECT 1375.590 4.000 1767.590 4.280 ;
        RECT 1768.430 4.000 2160.430 4.280 ;
        RECT 2161.270 4.000 2553.270 4.280 ;
        RECT 2554.110 4.000 2741.050 4.280 ;
      LAYER met3 ;
        RECT 4.000 3365.000 2746.000 3389.285 ;
        RECT 4.400 3363.600 2745.600 3365.000 ;
        RECT 4.000 3294.280 2746.000 3363.600 ;
        RECT 4.400 3292.880 2745.600 3294.280 ;
        RECT 4.000 3223.560 2746.000 3292.880 ;
        RECT 4.400 3222.160 2745.600 3223.560 ;
        RECT 4.000 3152.840 2746.000 3222.160 ;
        RECT 4.400 3151.440 2745.600 3152.840 ;
        RECT 4.000 3082.120 2746.000 3151.440 ;
        RECT 4.400 3080.720 2745.600 3082.120 ;
        RECT 4.000 3011.400 2746.000 3080.720 ;
        RECT 4.400 3010.000 2745.600 3011.400 ;
        RECT 4.000 2940.000 2746.000 3010.000 ;
        RECT 4.400 2938.600 2745.600 2940.000 ;
        RECT 4.000 2869.280 2746.000 2938.600 ;
        RECT 4.400 2867.880 2745.600 2869.280 ;
        RECT 4.000 2798.560 2746.000 2867.880 ;
        RECT 4.400 2797.160 2745.600 2798.560 ;
        RECT 4.000 2727.840 2746.000 2797.160 ;
        RECT 4.400 2726.440 2745.600 2727.840 ;
        RECT 4.000 2657.120 2746.000 2726.440 ;
        RECT 4.400 2655.720 2745.600 2657.120 ;
        RECT 4.000 2586.400 2746.000 2655.720 ;
        RECT 4.400 2585.000 2745.600 2586.400 ;
        RECT 4.000 2515.000 2746.000 2585.000 ;
        RECT 4.400 2513.600 2745.600 2515.000 ;
        RECT 4.000 2444.280 2746.000 2513.600 ;
        RECT 4.400 2442.880 2745.600 2444.280 ;
        RECT 4.000 2373.560 2746.000 2442.880 ;
        RECT 4.400 2372.160 2745.600 2373.560 ;
        RECT 4.000 2302.840 2746.000 2372.160 ;
        RECT 4.400 2301.440 2745.600 2302.840 ;
        RECT 4.000 2232.120 2746.000 2301.440 ;
        RECT 4.400 2230.720 2745.600 2232.120 ;
        RECT 4.000 2161.400 2746.000 2230.720 ;
        RECT 4.400 2160.000 2745.600 2161.400 ;
        RECT 4.000 2090.000 2746.000 2160.000 ;
        RECT 4.400 2088.600 2745.600 2090.000 ;
        RECT 4.000 2019.280 2746.000 2088.600 ;
        RECT 4.400 2017.880 2745.600 2019.280 ;
        RECT 4.000 1948.560 2746.000 2017.880 ;
        RECT 4.400 1947.160 2745.600 1948.560 ;
        RECT 4.000 1877.840 2746.000 1947.160 ;
        RECT 4.400 1876.440 2745.600 1877.840 ;
        RECT 4.000 1807.120 2746.000 1876.440 ;
        RECT 4.400 1805.720 2745.600 1807.120 ;
        RECT 4.000 1736.400 2746.000 1805.720 ;
        RECT 4.400 1735.000 2745.600 1736.400 ;
        RECT 4.000 1665.000 2746.000 1735.000 ;
        RECT 4.400 1663.600 2745.600 1665.000 ;
        RECT 4.000 1594.280 2746.000 1663.600 ;
        RECT 4.400 1592.880 2745.600 1594.280 ;
        RECT 4.000 1523.560 2746.000 1592.880 ;
        RECT 4.400 1522.160 2745.600 1523.560 ;
        RECT 4.000 1452.840 2746.000 1522.160 ;
        RECT 4.400 1451.440 2745.600 1452.840 ;
        RECT 4.000 1382.120 2746.000 1451.440 ;
        RECT 4.400 1380.720 2745.600 1382.120 ;
        RECT 4.000 1311.400 2746.000 1380.720 ;
        RECT 4.400 1310.000 2745.600 1311.400 ;
        RECT 4.000 1240.000 2746.000 1310.000 ;
        RECT 4.400 1238.600 2745.600 1240.000 ;
        RECT 4.000 1169.280 2746.000 1238.600 ;
        RECT 4.400 1167.880 2745.600 1169.280 ;
        RECT 4.000 1098.560 2746.000 1167.880 ;
        RECT 4.400 1097.160 2745.600 1098.560 ;
        RECT 4.000 1027.840 2746.000 1097.160 ;
        RECT 4.400 1026.440 2745.600 1027.840 ;
        RECT 4.000 957.120 2746.000 1026.440 ;
        RECT 4.400 955.720 2745.600 957.120 ;
        RECT 4.000 886.400 2746.000 955.720 ;
        RECT 4.400 885.000 2745.600 886.400 ;
        RECT 4.000 815.000 2746.000 885.000 ;
        RECT 4.400 813.600 2745.600 815.000 ;
        RECT 4.000 744.280 2746.000 813.600 ;
        RECT 4.400 742.880 2745.600 744.280 ;
        RECT 4.000 673.560 2746.000 742.880 ;
        RECT 4.400 672.160 2745.600 673.560 ;
        RECT 4.000 602.840 2746.000 672.160 ;
        RECT 4.400 601.440 2745.600 602.840 ;
        RECT 4.000 532.120 2746.000 601.440 ;
        RECT 4.400 530.720 2745.600 532.120 ;
        RECT 4.000 461.400 2746.000 530.720 ;
        RECT 4.400 460.000 2745.600 461.400 ;
        RECT 4.000 390.000 2746.000 460.000 ;
        RECT 4.400 388.600 2745.600 390.000 ;
        RECT 4.000 319.280 2746.000 388.600 ;
        RECT 4.400 317.880 2745.600 319.280 ;
        RECT 4.000 248.560 2746.000 317.880 ;
        RECT 4.400 247.160 2745.600 248.560 ;
        RECT 4.000 177.840 2746.000 247.160 ;
        RECT 4.400 176.440 2745.600 177.840 ;
        RECT 4.000 107.120 2746.000 176.440 ;
        RECT 4.400 105.720 2745.600 107.120 ;
        RECT 4.000 36.400 2746.000 105.720 ;
        RECT 4.400 35.000 2745.600 36.400 ;
        RECT 4.000 10.715 2746.000 35.000 ;
      LAYER met4 ;
        RECT 135.535 11.735 174.240 3388.265 ;
        RECT 176.640 11.735 251.040 3388.265 ;
        RECT 253.440 11.735 327.840 3388.265 ;
        RECT 330.240 11.735 404.640 3388.265 ;
        RECT 407.040 11.735 481.440 3388.265 ;
        RECT 483.840 11.735 558.240 3388.265 ;
        RECT 560.640 11.735 635.040 3388.265 ;
        RECT 637.440 11.735 711.840 3388.265 ;
        RECT 714.240 11.735 788.640 3388.265 ;
        RECT 791.040 11.735 865.440 3388.265 ;
        RECT 867.840 11.735 942.240 3388.265 ;
        RECT 944.640 11.735 1019.040 3388.265 ;
        RECT 1021.440 11.735 1095.840 3388.265 ;
        RECT 1098.240 11.735 1172.640 3388.265 ;
        RECT 1175.040 11.735 1249.440 3388.265 ;
        RECT 1251.840 11.735 1326.240 3388.265 ;
        RECT 1328.640 11.735 1403.040 3388.265 ;
        RECT 1405.440 11.735 1479.840 3388.265 ;
        RECT 1482.240 11.735 1556.640 3388.265 ;
        RECT 1559.040 11.735 1633.440 3388.265 ;
        RECT 1635.840 11.735 1710.240 3388.265 ;
        RECT 1712.640 11.735 1787.040 3388.265 ;
        RECT 1789.440 11.735 1863.840 3388.265 ;
        RECT 1866.240 11.735 1940.640 3388.265 ;
        RECT 1943.040 11.735 2017.440 3388.265 ;
        RECT 2019.840 11.735 2094.240 3388.265 ;
        RECT 2096.640 11.735 2171.040 3388.265 ;
        RECT 2173.440 11.735 2247.840 3388.265 ;
        RECT 2250.240 11.735 2324.640 3388.265 ;
        RECT 2327.040 11.735 2401.440 3388.265 ;
        RECT 2403.840 11.735 2478.240 3388.265 ;
        RECT 2480.640 11.735 2481.865 3388.265 ;
  END
END top
END LIBRARY

