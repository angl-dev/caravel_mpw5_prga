VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2750.000 BY 3600.000 ;
  PIN ipin_x0y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END ipin_x0y1_0
  PIN ipin_x0y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END ipin_x0y1_1
  PIN ipin_x0y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END ipin_x0y2_0
  PIN ipin_x0y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END ipin_x0y2_1
  PIN ipin_x0y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END ipin_x0y3_0
  PIN ipin_x0y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END ipin_x0y3_1
  PIN ipin_x0y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END ipin_x0y4_0
  PIN ipin_x0y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END ipin_x0y4_1
  PIN ipin_x0y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END ipin_x0y5_0
  PIN ipin_x0y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END ipin_x0y5_1
  PIN ipin_x0y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.800 4.000 787.400 ;
    END
  END ipin_x0y6_0
  PIN ipin_x0y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END ipin_x0y6_1
  PIN ipin_x0y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END ipin_x0y7_0
  PIN ipin_x0y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END ipin_x0y7_1
  PIN ipin_x0y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1087.360 4.000 1087.960 ;
    END
  END ipin_x0y8_0
  PIN ipin_x0y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END ipin_x0y8_1
  PIN ipin_x1y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 3596.000 28.890 3600.000 ;
    END
  END ipin_x1y9_0
  PIN ipin_x1y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 3596.000 85.930 3600.000 ;
    END
  END ipin_x1y9_1
  PIN ipin_x2y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 3596.000 143.430 3600.000 ;
    END
  END ipin_x2y9_0
  PIN ipin_x2y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 3596.000 200.470 3600.000 ;
    END
  END ipin_x2y9_1
  PIN ipin_x3y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 3596.000 257.970 3600.000 ;
    END
  END ipin_x3y9_0
  PIN ipin_x3y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 3596.000 315.010 3600.000 ;
    END
  END ipin_x3y9_1
  PIN ipin_x4y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 3596.000 372.510 3600.000 ;
    END
  END ipin_x4y9_0
  PIN ipin_x4y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 3596.000 429.550 3600.000 ;
    END
  END ipin_x4y9_1
  PIN ipin_x5y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 3596.000 487.050 3600.000 ;
    END
  END ipin_x5y9_0
  PIN ipin_x5y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 3596.000 544.090 3600.000 ;
    END
  END ipin_x5y9_1
  PIN ipin_x6y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 3596.000 601.590 3600.000 ;
    END
  END ipin_x6y9_0
  PIN ipin_x6y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 3596.000 658.630 3600.000 ;
    END
  END ipin_x6y9_1
  PIN ipin_x7y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 3596.000 716.130 3600.000 ;
    END
  END ipin_x7y9_0
  PIN ipin_x7y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 3596.000 773.630 3600.000 ;
    END
  END ipin_x7y9_1
  PIN ipin_x8y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 3596.000 830.670 3600.000 ;
    END
  END ipin_x8y9_0
  PIN ipin_x8y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 3596.000 888.170 3600.000 ;
    END
  END ipin_x8y9_1
  PIN ipin_x9y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 37.440 2750.000 38.040 ;
    END
  END ipin_x9y1_0
  PIN ipin_x9y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 112.240 2750.000 112.840 ;
    END
  END ipin_x9y1_1
  PIN ipin_x9y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 187.040 2750.000 187.640 ;
    END
  END ipin_x9y2_0
  PIN ipin_x9y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 261.840 2750.000 262.440 ;
    END
  END ipin_x9y2_1
  PIN ipin_x9y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 337.320 2750.000 337.920 ;
    END
  END ipin_x9y3_0
  PIN ipin_x9y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 412.120 2750.000 412.720 ;
    END
  END ipin_x9y3_1
  PIN ipin_x9y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 486.920 2750.000 487.520 ;
    END
  END ipin_x9y4_0
  PIN ipin_x9y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 562.400 2750.000 563.000 ;
    END
  END ipin_x9y4_1
  PIN ipin_x9y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 637.200 2750.000 637.800 ;
    END
  END ipin_x9y5_0
  PIN ipin_x9y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 712.000 2750.000 712.600 ;
    END
  END ipin_x9y5_1
  PIN ipin_x9y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 786.800 2750.000 787.400 ;
    END
  END ipin_x9y6_0
  PIN ipin_x9y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 862.280 2750.000 862.880 ;
    END
  END ipin_x9y6_1
  PIN ipin_x9y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 937.080 2750.000 937.680 ;
    END
  END ipin_x9y7_0
  PIN ipin_x9y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1011.880 2750.000 1012.480 ;
    END
  END ipin_x9y7_1
  PIN ipin_x9y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1087.360 2750.000 1087.960 ;
    END
  END ipin_x9y8_0
  PIN ipin_x9y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1162.160 2750.000 1162.760 ;
    END
  END ipin_x9y8_1
  PIN oe_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2437.160 4.000 2437.760 ;
    END
  END oe_x0y1_0
  PIN oe_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2511.960 4.000 2512.560 ;
    END
  END oe_x0y1_1
  PIN oe_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2586.760 4.000 2587.360 ;
    END
  END oe_x0y2_0
  PIN oe_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2662.240 4.000 2662.840 ;
    END
  END oe_x0y2_1
  PIN oe_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2737.040 4.000 2737.640 ;
    END
  END oe_x0y3_0
  PIN oe_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2811.840 4.000 2812.440 ;
    END
  END oe_x0y3_1
  PIN oe_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2887.320 4.000 2887.920 ;
    END
  END oe_x0y4_0
  PIN oe_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2962.120 4.000 2962.720 ;
    END
  END oe_x0y4_1
  PIN oe_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3036.920 4.000 3037.520 ;
    END
  END oe_x0y5_0
  PIN oe_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3111.720 4.000 3112.320 ;
    END
  END oe_x0y5_1
  PIN oe_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3187.200 4.000 3187.800 ;
    END
  END oe_x0y6_0
  PIN oe_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3262.000 4.000 3262.600 ;
    END
  END oe_x0y6_1
  PIN oe_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3336.800 4.000 3337.400 ;
    END
  END oe_x0y7_0
  PIN oe_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3412.280 4.000 3412.880 ;
    END
  END oe_x0y7_1
  PIN oe_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3487.080 4.000 3487.680 ;
    END
  END oe_x0y8_0
  PIN oe_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3561.880 4.000 3562.480 ;
    END
  END oe_x0y8_1
  PIN oe_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 3596.000 1861.990 3600.000 ;
    END
  END oe_x1y9_0
  PIN oe_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.750 3596.000 1919.030 3600.000 ;
    END
  END oe_x1y9_1
  PIN oe_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.250 3596.000 1976.530 3600.000 ;
    END
  END oe_x2y9_0
  PIN oe_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.290 3596.000 2033.570 3600.000 ;
    END
  END oe_x2y9_1
  PIN oe_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.790 3596.000 2091.070 3600.000 ;
    END
  END oe_x3y9_0
  PIN oe_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.290 3596.000 2148.570 3600.000 ;
    END
  END oe_x3y9_1
  PIN oe_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.330 3596.000 2205.610 3600.000 ;
    END
  END oe_x4y9_0
  PIN oe_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.830 3596.000 2263.110 3600.000 ;
    END
  END oe_x4y9_1
  PIN oe_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.870 3596.000 2320.150 3600.000 ;
    END
  END oe_x5y9_0
  PIN oe_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2377.370 3596.000 2377.650 3600.000 ;
    END
  END oe_x5y9_1
  PIN oe_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.410 3596.000 2434.690 3600.000 ;
    END
  END oe_x6y9_0
  PIN oe_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.910 3596.000 2492.190 3600.000 ;
    END
  END oe_x6y9_1
  PIN oe_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2548.950 3596.000 2549.230 3600.000 ;
    END
  END oe_x7y9_0
  PIN oe_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2606.450 3596.000 2606.730 3600.000 ;
    END
  END oe_x7y9_1
  PIN oe_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2663.490 3596.000 2663.770 3600.000 ;
    END
  END oe_x8y9_0
  PIN oe_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.990 3596.000 2721.270 3600.000 ;
    END
  END oe_x8y9_1
  PIN oe_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2437.160 2750.000 2437.760 ;
    END
  END oe_x9y1_0
  PIN oe_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2511.960 2750.000 2512.560 ;
    END
  END oe_x9y1_1
  PIN oe_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2586.760 2750.000 2587.360 ;
    END
  END oe_x9y2_0
  PIN oe_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2662.240 2750.000 2662.840 ;
    END
  END oe_x9y2_1
  PIN oe_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2737.040 2750.000 2737.640 ;
    END
  END oe_x9y3_0
  PIN oe_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2811.840 2750.000 2812.440 ;
    END
  END oe_x9y3_1
  PIN oe_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2887.320 2750.000 2887.920 ;
    END
  END oe_x9y4_0
  PIN oe_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2962.120 2750.000 2962.720 ;
    END
  END oe_x9y4_1
  PIN oe_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3036.920 2750.000 3037.520 ;
    END
  END oe_x9y5_0
  PIN oe_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3111.720 2750.000 3112.320 ;
    END
  END oe_x9y5_1
  PIN oe_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3187.200 2750.000 3187.800 ;
    END
  END oe_x9y6_0
  PIN oe_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3262.000 2750.000 3262.600 ;
    END
  END oe_x9y6_1
  PIN oe_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3336.800 2750.000 3337.400 ;
    END
  END oe_x9y7_0
  PIN oe_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3412.280 2750.000 3412.880 ;
    END
  END oe_x9y7_1
  PIN oe_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3487.080 2750.000 3487.680 ;
    END
  END oe_x9y8_0
  PIN oe_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 3561.880 2750.000 3562.480 ;
    END
  END oe_x9y8_1
  PIN opin_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.960 4.000 1237.560 ;
    END
  END opin_x0y1_0
  PIN opin_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.760 4.000 1312.360 ;
    END
  END opin_x0y1_1
  PIN opin_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END opin_x0y2_0
  PIN opin_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END opin_x0y2_1
  PIN opin_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END opin_x0y3_0
  PIN opin_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1612.320 4.000 1612.920 ;
    END
  END opin_x0y3_1
  PIN opin_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1687.120 4.000 1687.720 ;
    END
  END opin_x0y4_0
  PIN opin_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1761.920 4.000 1762.520 ;
    END
  END opin_x0y4_1
  PIN opin_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1837.400 4.000 1838.000 ;
    END
  END opin_x0y5_0
  PIN opin_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1912.200 4.000 1912.800 ;
    END
  END opin_x0y5_1
  PIN opin_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1987.000 4.000 1987.600 ;
    END
  END opin_x0y6_0
  PIN opin_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2061.800 4.000 2062.400 ;
    END
  END opin_x0y6_1
  PIN opin_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2137.280 4.000 2137.880 ;
    END
  END opin_x0y7_0
  PIN opin_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2212.080 4.000 2212.680 ;
    END
  END opin_x0y7_1
  PIN opin_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2286.880 4.000 2287.480 ;
    END
  END opin_x0y8_0
  PIN opin_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2362.360 4.000 2362.960 ;
    END
  END opin_x0y8_1
  PIN opin_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 3596.000 945.210 3600.000 ;
    END
  END opin_x1y9_0
  PIN opin_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 3596.000 1002.710 3600.000 ;
    END
  END opin_x1y9_1
  PIN opin_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 3596.000 1059.750 3600.000 ;
    END
  END opin_x2y9_0
  PIN opin_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 3596.000 1117.250 3600.000 ;
    END
  END opin_x2y9_1
  PIN opin_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 3596.000 1174.290 3600.000 ;
    END
  END opin_x3y9_0
  PIN opin_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.510 3596.000 1231.790 3600.000 ;
    END
  END opin_x3y9_1
  PIN opin_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.550 3596.000 1288.830 3600.000 ;
    END
  END opin_x4y9_0
  PIN opin_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 3596.000 1346.330 3600.000 ;
    END
  END opin_x4y9_1
  PIN opin_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.550 3596.000 1403.830 3600.000 ;
    END
  END opin_x5y9_0
  PIN opin_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.590 3596.000 1460.870 3600.000 ;
    END
  END opin_x5y9_1
  PIN opin_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 3596.000 1518.370 3600.000 ;
    END
  END opin_x6y9_0
  PIN opin_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 3596.000 1575.410 3600.000 ;
    END
  END opin_x6y9_1
  PIN opin_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 3596.000 1632.910 3600.000 ;
    END
  END opin_x7y9_0
  PIN opin_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 3596.000 1689.950 3600.000 ;
    END
  END opin_x7y9_1
  PIN opin_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 3596.000 1747.450 3600.000 ;
    END
  END opin_x8y9_0
  PIN opin_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.210 3596.000 1804.490 3600.000 ;
    END
  END opin_x8y9_1
  PIN opin_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1236.960 2750.000 1237.560 ;
    END
  END opin_x9y1_0
  PIN opin_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1311.760 2750.000 1312.360 ;
    END
  END opin_x9y1_1
  PIN opin_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1387.240 2750.000 1387.840 ;
    END
  END opin_x9y2_0
  PIN opin_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1462.040 2750.000 1462.640 ;
    END
  END opin_x9y2_1
  PIN opin_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1536.840 2750.000 1537.440 ;
    END
  END opin_x9y3_0
  PIN opin_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1612.320 2750.000 1612.920 ;
    END
  END opin_x9y3_1
  PIN opin_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1687.120 2750.000 1687.720 ;
    END
  END opin_x9y4_0
  PIN opin_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1761.920 2750.000 1762.520 ;
    END
  END opin_x9y4_1
  PIN opin_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1837.400 2750.000 1838.000 ;
    END
  END opin_x9y5_0
  PIN opin_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1912.200 2750.000 1912.800 ;
    END
  END opin_x9y5_1
  PIN opin_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 1987.000 2750.000 1987.600 ;
    END
  END opin_x9y6_0
  PIN opin_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2061.800 2750.000 2062.400 ;
    END
  END opin_x9y6_1
  PIN opin_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2137.280 2750.000 2137.880 ;
    END
  END opin_x9y7_0
  PIN opin_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2212.080 2750.000 2212.680 ;
    END
  END opin_x9y7_1
  PIN opin_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2286.880 2750.000 2287.480 ;
    END
  END opin_x9y8_0
  PIN opin_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2746.000 2362.360 2750.000 2362.960 ;
    END
  END opin_x9y8_1
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END prog_clk
  PIN prog_din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END prog_din
  PIN prog_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END prog_done
  PIN prog_dout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END prog_dout
  PIN prog_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 0.000 1768.150 4.000 ;
    END
  END prog_rst
  PIN prog_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.710 0.000 2160.990 4.000 ;
    END
  END prog_we
  PIN prog_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2553.550 0.000 2553.830 4.000 ;
    END
  END prog_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 3587.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 3587.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 3587.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2744.360 3587.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 2744.360 3587.920 ;
      LAYER met2 ;
        RECT 6.990 3595.720 28.330 3596.250 ;
        RECT 29.170 3595.720 85.370 3596.250 ;
        RECT 86.210 3595.720 142.870 3596.250 ;
        RECT 143.710 3595.720 199.910 3596.250 ;
        RECT 200.750 3595.720 257.410 3596.250 ;
        RECT 258.250 3595.720 314.450 3596.250 ;
        RECT 315.290 3595.720 371.950 3596.250 ;
        RECT 372.790 3595.720 428.990 3596.250 ;
        RECT 429.830 3595.720 486.490 3596.250 ;
        RECT 487.330 3595.720 543.530 3596.250 ;
        RECT 544.370 3595.720 601.030 3596.250 ;
        RECT 601.870 3595.720 658.070 3596.250 ;
        RECT 658.910 3595.720 715.570 3596.250 ;
        RECT 716.410 3595.720 773.070 3596.250 ;
        RECT 773.910 3595.720 830.110 3596.250 ;
        RECT 830.950 3595.720 887.610 3596.250 ;
        RECT 888.450 3595.720 944.650 3596.250 ;
        RECT 945.490 3595.720 1002.150 3596.250 ;
        RECT 1002.990 3595.720 1059.190 3596.250 ;
        RECT 1060.030 3595.720 1116.690 3596.250 ;
        RECT 1117.530 3595.720 1173.730 3596.250 ;
        RECT 1174.570 3595.720 1231.230 3596.250 ;
        RECT 1232.070 3595.720 1288.270 3596.250 ;
        RECT 1289.110 3595.720 1345.770 3596.250 ;
        RECT 1346.610 3595.720 1403.270 3596.250 ;
        RECT 1404.110 3595.720 1460.310 3596.250 ;
        RECT 1461.150 3595.720 1517.810 3596.250 ;
        RECT 1518.650 3595.720 1574.850 3596.250 ;
        RECT 1575.690 3595.720 1632.350 3596.250 ;
        RECT 1633.190 3595.720 1689.390 3596.250 ;
        RECT 1690.230 3595.720 1746.890 3596.250 ;
        RECT 1747.730 3595.720 1803.930 3596.250 ;
        RECT 1804.770 3595.720 1861.430 3596.250 ;
        RECT 1862.270 3595.720 1918.470 3596.250 ;
        RECT 1919.310 3595.720 1975.970 3596.250 ;
        RECT 1976.810 3595.720 2033.010 3596.250 ;
        RECT 2033.850 3595.720 2090.510 3596.250 ;
        RECT 2091.350 3595.720 2148.010 3596.250 ;
        RECT 2148.850 3595.720 2205.050 3596.250 ;
        RECT 2205.890 3595.720 2262.550 3596.250 ;
        RECT 2263.390 3595.720 2319.590 3596.250 ;
        RECT 2320.430 3595.720 2377.090 3596.250 ;
        RECT 2377.930 3595.720 2434.130 3596.250 ;
        RECT 2434.970 3595.720 2491.630 3596.250 ;
        RECT 2492.470 3595.720 2548.670 3596.250 ;
        RECT 2549.510 3595.720 2606.170 3596.250 ;
        RECT 2607.010 3595.720 2663.210 3596.250 ;
        RECT 2664.050 3595.720 2720.710 3596.250 ;
        RECT 2721.550 3595.720 2741.050 3596.250 ;
        RECT 6.990 4.280 2741.050 3595.720 ;
        RECT 6.990 4.000 196.230 4.280 ;
        RECT 197.070 4.000 589.070 4.280 ;
        RECT 589.910 4.000 981.910 4.280 ;
        RECT 982.750 4.000 1374.750 4.280 ;
        RECT 1375.590 4.000 1767.590 4.280 ;
        RECT 1768.430 4.000 2160.430 4.280 ;
        RECT 2161.270 4.000 2553.270 4.280 ;
        RECT 2554.110 4.000 2741.050 4.280 ;
      LAYER met3 ;
        RECT 4.000 3562.880 2746.000 3587.845 ;
        RECT 4.400 3561.480 2745.600 3562.880 ;
        RECT 4.000 3488.080 2746.000 3561.480 ;
        RECT 4.400 3486.680 2745.600 3488.080 ;
        RECT 4.000 3413.280 2746.000 3486.680 ;
        RECT 4.400 3411.880 2745.600 3413.280 ;
        RECT 4.000 3337.800 2746.000 3411.880 ;
        RECT 4.400 3336.400 2745.600 3337.800 ;
        RECT 4.000 3263.000 2746.000 3336.400 ;
        RECT 4.400 3261.600 2745.600 3263.000 ;
        RECT 4.000 3188.200 2746.000 3261.600 ;
        RECT 4.400 3186.800 2745.600 3188.200 ;
        RECT 4.000 3112.720 2746.000 3186.800 ;
        RECT 4.400 3111.320 2745.600 3112.720 ;
        RECT 4.000 3037.920 2746.000 3111.320 ;
        RECT 4.400 3036.520 2745.600 3037.920 ;
        RECT 4.000 2963.120 2746.000 3036.520 ;
        RECT 4.400 2961.720 2745.600 2963.120 ;
        RECT 4.000 2888.320 2746.000 2961.720 ;
        RECT 4.400 2886.920 2745.600 2888.320 ;
        RECT 4.000 2812.840 2746.000 2886.920 ;
        RECT 4.400 2811.440 2745.600 2812.840 ;
        RECT 4.000 2738.040 2746.000 2811.440 ;
        RECT 4.400 2736.640 2745.600 2738.040 ;
        RECT 4.000 2663.240 2746.000 2736.640 ;
        RECT 4.400 2661.840 2745.600 2663.240 ;
        RECT 4.000 2587.760 2746.000 2661.840 ;
        RECT 4.400 2586.360 2745.600 2587.760 ;
        RECT 4.000 2512.960 2746.000 2586.360 ;
        RECT 4.400 2511.560 2745.600 2512.960 ;
        RECT 4.000 2438.160 2746.000 2511.560 ;
        RECT 4.400 2436.760 2745.600 2438.160 ;
        RECT 4.000 2363.360 2746.000 2436.760 ;
        RECT 4.400 2361.960 2745.600 2363.360 ;
        RECT 4.000 2287.880 2746.000 2361.960 ;
        RECT 4.400 2286.480 2745.600 2287.880 ;
        RECT 4.000 2213.080 2746.000 2286.480 ;
        RECT 4.400 2211.680 2745.600 2213.080 ;
        RECT 4.000 2138.280 2746.000 2211.680 ;
        RECT 4.400 2136.880 2745.600 2138.280 ;
        RECT 4.000 2062.800 2746.000 2136.880 ;
        RECT 4.400 2061.400 2745.600 2062.800 ;
        RECT 4.000 1988.000 2746.000 2061.400 ;
        RECT 4.400 1986.600 2745.600 1988.000 ;
        RECT 4.000 1913.200 2746.000 1986.600 ;
        RECT 4.400 1911.800 2745.600 1913.200 ;
        RECT 4.000 1838.400 2746.000 1911.800 ;
        RECT 4.400 1837.000 2745.600 1838.400 ;
        RECT 4.000 1762.920 2746.000 1837.000 ;
        RECT 4.400 1761.520 2745.600 1762.920 ;
        RECT 4.000 1688.120 2746.000 1761.520 ;
        RECT 4.400 1686.720 2745.600 1688.120 ;
        RECT 4.000 1613.320 2746.000 1686.720 ;
        RECT 4.400 1611.920 2745.600 1613.320 ;
        RECT 4.000 1537.840 2746.000 1611.920 ;
        RECT 4.400 1536.440 2745.600 1537.840 ;
        RECT 4.000 1463.040 2746.000 1536.440 ;
        RECT 4.400 1461.640 2745.600 1463.040 ;
        RECT 4.000 1388.240 2746.000 1461.640 ;
        RECT 4.400 1386.840 2745.600 1388.240 ;
        RECT 4.000 1312.760 2746.000 1386.840 ;
        RECT 4.400 1311.360 2745.600 1312.760 ;
        RECT 4.000 1237.960 2746.000 1311.360 ;
        RECT 4.400 1236.560 2745.600 1237.960 ;
        RECT 4.000 1163.160 2746.000 1236.560 ;
        RECT 4.400 1161.760 2745.600 1163.160 ;
        RECT 4.000 1088.360 2746.000 1161.760 ;
        RECT 4.400 1086.960 2745.600 1088.360 ;
        RECT 4.000 1012.880 2746.000 1086.960 ;
        RECT 4.400 1011.480 2745.600 1012.880 ;
        RECT 4.000 938.080 2746.000 1011.480 ;
        RECT 4.400 936.680 2745.600 938.080 ;
        RECT 4.000 863.280 2746.000 936.680 ;
        RECT 4.400 861.880 2745.600 863.280 ;
        RECT 4.000 787.800 2746.000 861.880 ;
        RECT 4.400 786.400 2745.600 787.800 ;
        RECT 4.000 713.000 2746.000 786.400 ;
        RECT 4.400 711.600 2745.600 713.000 ;
        RECT 4.000 638.200 2746.000 711.600 ;
        RECT 4.400 636.800 2745.600 638.200 ;
        RECT 4.000 563.400 2746.000 636.800 ;
        RECT 4.400 562.000 2745.600 563.400 ;
        RECT 4.000 487.920 2746.000 562.000 ;
        RECT 4.400 486.520 2745.600 487.920 ;
        RECT 4.000 413.120 2746.000 486.520 ;
        RECT 4.400 411.720 2745.600 413.120 ;
        RECT 4.000 338.320 2746.000 411.720 ;
        RECT 4.400 336.920 2745.600 338.320 ;
        RECT 4.000 262.840 2746.000 336.920 ;
        RECT 4.400 261.440 2745.600 262.840 ;
        RECT 4.000 188.040 2746.000 261.440 ;
        RECT 4.400 186.640 2745.600 188.040 ;
        RECT 4.000 113.240 2746.000 186.640 ;
        RECT 4.400 111.840 2745.600 113.240 ;
        RECT 4.000 38.440 2746.000 111.840 ;
        RECT 4.400 37.040 2745.600 38.440 ;
        RECT 4.000 10.715 2746.000 37.040 ;
      LAYER met4 ;
        RECT 164.975 11.735 174.240 3586.145 ;
        RECT 176.640 11.735 251.040 3586.145 ;
        RECT 253.440 11.735 327.840 3586.145 ;
        RECT 330.240 11.735 404.640 3586.145 ;
        RECT 407.040 11.735 481.440 3586.145 ;
        RECT 483.840 11.735 558.240 3586.145 ;
        RECT 560.640 11.735 635.040 3586.145 ;
        RECT 637.440 11.735 711.840 3586.145 ;
        RECT 714.240 11.735 788.640 3586.145 ;
        RECT 791.040 11.735 865.440 3586.145 ;
        RECT 867.840 11.735 942.240 3586.145 ;
        RECT 944.640 11.735 1019.040 3586.145 ;
        RECT 1021.440 11.735 1095.840 3586.145 ;
        RECT 1098.240 11.735 1172.640 3586.145 ;
        RECT 1175.040 11.735 1249.440 3586.145 ;
        RECT 1251.840 11.735 1326.240 3586.145 ;
        RECT 1328.640 11.735 1403.040 3586.145 ;
        RECT 1405.440 11.735 1479.840 3586.145 ;
        RECT 1482.240 11.735 1556.640 3586.145 ;
        RECT 1559.040 11.735 1633.440 3586.145 ;
        RECT 1635.840 11.735 1710.240 3586.145 ;
        RECT 1712.640 11.735 1787.040 3586.145 ;
        RECT 1789.440 11.735 1863.840 3586.145 ;
        RECT 1866.240 11.735 1940.640 3586.145 ;
        RECT 1943.040 11.735 2017.440 3586.145 ;
        RECT 2019.840 11.735 2094.240 3586.145 ;
        RECT 2096.640 11.735 2171.040 3586.145 ;
        RECT 2173.440 11.735 2247.840 3586.145 ;
        RECT 2250.240 11.735 2324.640 3586.145 ;
        RECT 2327.040 11.735 2401.440 3586.145 ;
        RECT 2403.840 11.735 2478.240 3586.145 ;
        RECT 2480.640 11.735 2481.865 3586.145 ;
  END
END top
END LIBRARY

