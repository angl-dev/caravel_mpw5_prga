magic
tech sky130A
magscale 1 2
timestamp 1653704188
<< obsli1 >>
rect 30424 29159 548200 664585
<< obsm1 >>
rect 2774 20612 580690 703044
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 2778 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 580686 703610
rect 2778 19751 580686 703464
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 560 697140 583440 697237
rect 480 697004 583440 697140
rect 480 684484 583520 697004
rect 560 684084 583520 684484
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19755 583440 19988
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 6914 -1894 7534 705830
rect 9234 -5734 9854 709670
rect 10634 -3814 11254 707750
rect 12034 -1894 12654 705830
rect 12954 -7654 13574 711590
rect 14354 -5734 14974 709670
rect 15754 -3814 16374 707750
rect 17154 -1894 17774 705830
rect 18074 -7654 18694 711590
rect 19474 -5734 20094 709670
rect 20874 -3814 21494 707750
rect 22274 -1894 22894 705830
rect 23194 -7654 23814 711590
rect 24594 -5734 25214 709670
rect 25994 -3814 26614 707750
rect 27394 669000 28014 705830
rect 28314 669000 28934 711590
rect 29714 669000 30334 709670
rect 31114 669000 31734 707750
rect 32514 669000 33134 705830
rect 33434 669000 34054 711590
rect 34834 669000 35454 709670
rect 36234 669000 36854 707750
rect 37634 669000 38254 705830
rect 38554 669000 39174 711590
rect 39954 669000 40574 709670
rect 41354 669000 41974 707750
rect 42754 669000 43374 705830
rect 43674 669000 44294 711590
rect 45074 669000 45694 709670
rect 46474 669000 47094 707750
rect 47874 669000 48494 705830
rect 48794 669000 49414 711590
rect 50194 669000 50814 709670
rect 51594 669000 52214 707750
rect 52994 669000 53614 705830
rect 53914 669000 54534 711590
rect 55314 669000 55934 709670
rect 56714 669000 57334 707750
rect 58114 669000 58734 705830
rect 59034 669000 59654 711590
rect 60434 669000 61054 709670
rect 61834 669000 62454 707750
rect 63234 669000 63854 705830
rect 64154 669000 64774 711590
rect 65554 669000 66174 709670
rect 66954 669000 67574 707750
rect 68354 669000 68974 705830
rect 69274 669000 69894 711590
rect 70674 669000 71294 709670
rect 72074 669000 72694 707750
rect 73474 669000 74094 705830
rect 74394 669000 75014 711590
rect 75794 669000 76414 709670
rect 77194 669000 77814 707750
rect 78594 669000 79214 705830
rect 79514 669000 80134 711590
rect 80914 669000 81534 709670
rect 82314 669000 82934 707750
rect 83714 669000 84334 705830
rect 84634 669000 85254 711590
rect 86034 669000 86654 709670
rect 87434 669000 88054 707750
rect 88834 669000 89454 705830
rect 89754 669000 90374 711590
rect 91154 669000 91774 709670
rect 92554 669000 93174 707750
rect 93954 669000 94574 705830
rect 94874 669000 95494 711590
rect 96274 669000 96894 709670
rect 97674 669000 98294 707750
rect 99074 669000 99694 705830
rect 99994 669000 100614 711590
rect 101394 669000 102014 709670
rect 102794 669000 103414 707750
rect 104194 669000 104814 705830
rect 105114 669000 105734 711590
rect 106514 669000 107134 709670
rect 107914 669000 108534 707750
rect 109314 669000 109934 705830
rect 110234 669000 110854 711590
rect 111634 669000 112254 709670
rect 113034 669000 113654 707750
rect 114434 669000 115054 705830
rect 115354 669000 115974 711590
rect 116754 669000 117374 709670
rect 118154 669000 118774 707750
rect 119554 669000 120174 705830
rect 120474 669000 121094 711590
rect 121874 669000 122494 709670
rect 123274 669000 123894 707750
rect 124674 669000 125294 705830
rect 125594 669000 126214 711590
rect 126994 669000 127614 709670
rect 128394 669000 129014 707750
rect 129794 669000 130414 705830
rect 130714 669000 131334 711590
rect 132114 669000 132734 709670
rect 133514 669000 134134 707750
rect 134914 669000 135534 705830
rect 135834 669000 136454 711590
rect 137234 669000 137854 709670
rect 138634 669000 139254 707750
rect 140034 669000 140654 705830
rect 140954 669000 141574 711590
rect 142354 669000 142974 709670
rect 143754 669000 144374 707750
rect 145154 669000 145774 705830
rect 146074 669000 146694 711590
rect 147474 669000 148094 709670
rect 148874 669000 149494 707750
rect 150274 669000 150894 705830
rect 151194 669000 151814 711590
rect 152594 669000 153214 709670
rect 153994 669000 154614 707750
rect 155394 669000 156014 705830
rect 156314 669000 156934 711590
rect 157714 669000 158334 709670
rect 159114 669000 159734 707750
rect 160514 669000 161134 705830
rect 161434 669000 162054 711590
rect 162834 669000 163454 709670
rect 164234 669000 164854 707750
rect 165634 669000 166254 705830
rect 166554 669000 167174 711590
rect 167954 669000 168574 709670
rect 169354 669000 169974 707750
rect 170754 669000 171374 705830
rect 171674 669000 172294 711590
rect 173074 669000 173694 709670
rect 174474 669000 175094 707750
rect 175874 669000 176494 705830
rect 176794 669000 177414 711590
rect 178194 669000 178814 709670
rect 179594 669000 180214 707750
rect 180994 669000 181614 705830
rect 181914 669000 182534 711590
rect 183314 669000 183934 709670
rect 184714 669000 185334 707750
rect 186114 669000 186734 705830
rect 187034 669000 187654 711590
rect 188434 669000 189054 709670
rect 189834 669000 190454 707750
rect 191234 669000 191854 705830
rect 192154 669000 192774 711590
rect 193554 669000 194174 709670
rect 194954 669000 195574 707750
rect 196354 669000 196974 705830
rect 197274 669000 197894 711590
rect 198674 669000 199294 709670
rect 200074 669000 200694 707750
rect 201474 669000 202094 705830
rect 202394 669000 203014 711590
rect 203794 669000 204414 709670
rect 205194 669000 205814 707750
rect 206594 669000 207214 705830
rect 207514 669000 208134 711590
rect 208914 669000 209534 709670
rect 210314 669000 210934 707750
rect 211714 669000 212334 705830
rect 212634 669000 213254 711590
rect 214034 669000 214654 709670
rect 215434 669000 216054 707750
rect 216834 669000 217454 705830
rect 217754 669000 218374 711590
rect 219154 669000 219774 709670
rect 220554 669000 221174 707750
rect 221954 669000 222574 705830
rect 222874 669000 223494 711590
rect 224274 669000 224894 709670
rect 225674 669000 226294 707750
rect 227074 669000 227694 705830
rect 227994 669000 228614 711590
rect 229394 669000 230014 709670
rect 230794 669000 231414 707750
rect 232194 669000 232814 705830
rect 233114 669000 233734 711590
rect 234514 669000 235134 709670
rect 235914 669000 236534 707750
rect 237314 669000 237934 705830
rect 238234 669000 238854 711590
rect 239634 669000 240254 709670
rect 241034 669000 241654 707750
rect 242434 669000 243054 705830
rect 243354 669000 243974 711590
rect 244754 669000 245374 709670
rect 246154 669000 246774 707750
rect 247554 669000 248174 705830
rect 248474 669000 249094 711590
rect 249874 669000 250494 709670
rect 251274 669000 251894 707750
rect 252674 669000 253294 705830
rect 253594 669000 254214 711590
rect 254994 669000 255614 709670
rect 256394 669000 257014 707750
rect 257794 669000 258414 705830
rect 258714 669000 259334 711590
rect 260114 669000 260734 709670
rect 261514 669000 262134 707750
rect 262914 669000 263534 705830
rect 263834 669000 264454 711590
rect 265234 669000 265854 709670
rect 266634 669000 267254 707750
rect 268034 669000 268654 705830
rect 268954 669000 269574 711590
rect 270354 669000 270974 709670
rect 271754 669000 272374 707750
rect 273154 669000 273774 705830
rect 274074 669000 274694 711590
rect 275474 669000 276094 709670
rect 276874 669000 277494 707750
rect 278274 669000 278894 705830
rect 279194 669000 279814 711590
rect 280594 669000 281214 709670
rect 281994 669000 282614 707750
rect 283394 669000 284014 705830
rect 284314 669000 284934 711590
rect 285714 669000 286334 709670
rect 287114 669000 287734 707750
rect 288514 669000 289134 705830
rect 289434 669000 290054 711590
rect 290834 669000 291454 709670
rect 292234 669000 292854 707750
rect 293634 669000 294254 705830
rect 294554 669000 295174 711590
rect 295954 669000 296574 709670
rect 297354 669000 297974 707750
rect 298754 669000 299374 705830
rect 299674 669000 300294 711590
rect 301074 669000 301694 709670
rect 302474 669000 303094 707750
rect 303874 669000 304494 705830
rect 304794 669000 305414 711590
rect 306194 669000 306814 709670
rect 307594 669000 308214 707750
rect 308994 669000 309614 705830
rect 309914 669000 310534 711590
rect 311314 669000 311934 709670
rect 312714 669000 313334 707750
rect 314114 669000 314734 705830
rect 315034 669000 315654 711590
rect 316434 669000 317054 709670
rect 317834 669000 318454 707750
rect 319234 669000 319854 705830
rect 320154 669000 320774 711590
rect 321554 669000 322174 709670
rect 322954 669000 323574 707750
rect 324354 669000 324974 705830
rect 325274 669000 325894 711590
rect 326674 669000 327294 709670
rect 328074 669000 328694 707750
rect 329474 669000 330094 705830
rect 330394 669000 331014 711590
rect 331794 669000 332414 709670
rect 333194 669000 333814 707750
rect 334594 669000 335214 705830
rect 335514 669000 336134 711590
rect 336914 669000 337534 709670
rect 338314 669000 338934 707750
rect 339714 669000 340334 705830
rect 340634 669000 341254 711590
rect 342034 669000 342654 709670
rect 343434 669000 344054 707750
rect 344834 669000 345454 705830
rect 345754 669000 346374 711590
rect 347154 669000 347774 709670
rect 348554 669000 349174 707750
rect 349954 669000 350574 705830
rect 350874 669000 351494 711590
rect 352274 669000 352894 709670
rect 353674 669000 354294 707750
rect 355074 669000 355694 705830
rect 355994 669000 356614 711590
rect 357394 669000 358014 709670
rect 358794 669000 359414 707750
rect 360194 669000 360814 705830
rect 361114 669000 361734 711590
rect 362514 669000 363134 709670
rect 363914 669000 364534 707750
rect 365314 669000 365934 705830
rect 366234 669000 366854 711590
rect 367634 669000 368254 709670
rect 369034 669000 369654 707750
rect 370434 669000 371054 705830
rect 371354 669000 371974 711590
rect 372754 669000 373374 709670
rect 374154 669000 374774 707750
rect 375554 669000 376174 705830
rect 376474 669000 377094 711590
rect 377874 669000 378494 709670
rect 379274 669000 379894 707750
rect 380674 669000 381294 705830
rect 381594 669000 382214 711590
rect 382994 669000 383614 709670
rect 384394 669000 385014 707750
rect 385794 669000 386414 705830
rect 386714 669000 387334 711590
rect 388114 669000 388734 709670
rect 389514 669000 390134 707750
rect 390914 669000 391534 705830
rect 391834 669000 392454 711590
rect 393234 669000 393854 709670
rect 394634 669000 395254 707750
rect 396034 669000 396654 705830
rect 396954 669000 397574 711590
rect 398354 669000 398974 709670
rect 399754 669000 400374 707750
rect 401154 669000 401774 705830
rect 402074 669000 402694 711590
rect 403474 669000 404094 709670
rect 404874 669000 405494 707750
rect 406274 669000 406894 705830
rect 407194 669000 407814 711590
rect 408594 669000 409214 709670
rect 409994 669000 410614 707750
rect 411394 669000 412014 705830
rect 412314 669000 412934 711590
rect 413714 669000 414334 709670
rect 415114 669000 415734 707750
rect 416514 669000 417134 705830
rect 417434 669000 418054 711590
rect 418834 669000 419454 709670
rect 420234 669000 420854 707750
rect 421634 669000 422254 705830
rect 422554 669000 423174 711590
rect 423954 669000 424574 709670
rect 425354 669000 425974 707750
rect 426754 669000 427374 705830
rect 427674 669000 428294 711590
rect 429074 669000 429694 709670
rect 430474 669000 431094 707750
rect 431874 669000 432494 705830
rect 432794 669000 433414 711590
rect 434194 669000 434814 709670
rect 435594 669000 436214 707750
rect 436994 669000 437614 705830
rect 437914 669000 438534 711590
rect 439314 669000 439934 709670
rect 440714 669000 441334 707750
rect 442114 669000 442734 705830
rect 443034 669000 443654 711590
rect 444434 669000 445054 709670
rect 445834 669000 446454 707750
rect 447234 669000 447854 705830
rect 448154 669000 448774 711590
rect 449554 669000 450174 709670
rect 450954 669000 451574 707750
rect 452354 669000 452974 705830
rect 453274 669000 453894 711590
rect 454674 669000 455294 709670
rect 456074 669000 456694 707750
rect 457474 669000 458094 705830
rect 458394 669000 459014 711590
rect 459794 669000 460414 709670
rect 461194 669000 461814 707750
rect 462594 669000 463214 705830
rect 463514 669000 464134 711590
rect 464914 669000 465534 709670
rect 466314 669000 466934 707750
rect 467714 669000 468334 705830
rect 468634 669000 469254 711590
rect 470034 669000 470654 709670
rect 471434 669000 472054 707750
rect 472834 669000 473454 705830
rect 473754 669000 474374 711590
rect 475154 669000 475774 709670
rect 476554 669000 477174 707750
rect 477954 669000 478574 705830
rect 478874 669000 479494 711590
rect 480274 669000 480894 709670
rect 481674 669000 482294 707750
rect 483074 669000 483694 705830
rect 483994 669000 484614 711590
rect 485394 669000 486014 709670
rect 486794 669000 487414 707750
rect 488194 669000 488814 705830
rect 489114 669000 489734 711590
rect 490514 669000 491134 709670
rect 491914 669000 492534 707750
rect 493314 669000 493934 705830
rect 494234 669000 494854 711590
rect 495634 669000 496254 709670
rect 497034 669000 497654 707750
rect 498434 669000 499054 705830
rect 499354 669000 499974 711590
rect 500754 669000 501374 709670
rect 502154 669000 502774 707750
rect 503554 669000 504174 705830
rect 504474 669000 505094 711590
rect 505874 669000 506494 709670
rect 507274 669000 507894 707750
rect 508674 669000 509294 705830
rect 509594 669000 510214 711590
rect 510994 669000 511614 709670
rect 512394 669000 513014 707750
rect 513794 669000 514414 705830
rect 514714 669000 515334 711590
rect 516114 669000 516734 709670
rect 517514 669000 518134 707750
rect 518914 669000 519534 705830
rect 519834 669000 520454 711590
rect 521234 669000 521854 709670
rect 522634 669000 523254 707750
rect 524034 669000 524654 705830
rect 524954 669000 525574 711590
rect 526354 669000 526974 709670
rect 527754 669000 528374 707750
rect 529154 669000 529774 705830
rect 530074 669000 530694 711590
rect 531474 669000 532094 709670
rect 532874 669000 533494 707750
rect 534274 669000 534894 705830
rect 535194 669000 535814 711590
rect 536594 669000 537214 709670
rect 537994 669000 538614 707750
rect 539394 669000 540014 705830
rect 540314 669000 540934 711590
rect 541714 669000 542334 709670
rect 543114 669000 543734 707750
rect 544514 669000 545134 705830
rect 545434 669000 546054 711590
rect 546834 669000 547454 709670
rect 548234 669000 548854 707750
rect 549634 669000 550254 705830
rect 550554 669000 551174 711590
rect 27394 -1894 28014 25000
rect 28314 -7654 28934 25000
rect 29714 -5734 30334 25000
rect 31114 -3814 31734 25000
rect 32514 -1894 33134 25000
rect 33434 -7654 34054 25000
rect 34834 -5734 35454 25000
rect 36234 -3814 36854 25000
rect 37634 -1894 38254 25000
rect 38554 -7654 39174 25000
rect 39954 -5734 40574 25000
rect 41354 -3814 41974 25000
rect 42754 -1894 43374 25000
rect 43674 -7654 44294 25000
rect 45074 -5734 45694 25000
rect 46474 -3814 47094 25000
rect 47874 -1894 48494 25000
rect 48794 -7654 49414 25000
rect 50194 -5734 50814 25000
rect 51594 -3814 52214 25000
rect 52994 -1894 53614 25000
rect 53914 -7654 54534 25000
rect 55314 -5734 55934 25000
rect 56714 -3814 57334 25000
rect 58114 -1894 58734 25000
rect 59034 -7654 59654 25000
rect 60434 -5734 61054 25000
rect 61834 -3814 62454 25000
rect 63234 -1894 63854 25000
rect 64154 -7654 64774 25000
rect 65554 -5734 66174 25000
rect 66954 -3814 67574 25000
rect 68354 -1894 68974 25000
rect 69274 -7654 69894 25000
rect 70674 -5734 71294 25000
rect 72074 -3814 72694 25000
rect 73474 -1894 74094 25000
rect 74394 -7654 75014 25000
rect 75794 -5734 76414 25000
rect 77194 -3814 77814 25000
rect 78594 -1894 79214 25000
rect 79514 -7654 80134 25000
rect 80914 -5734 81534 25000
rect 82314 -3814 82934 25000
rect 83714 -1894 84334 25000
rect 84634 -7654 85254 25000
rect 86034 -5734 86654 25000
rect 87434 -3814 88054 25000
rect 88834 -1894 89454 25000
rect 89754 -7654 90374 25000
rect 91154 -5734 91774 25000
rect 92554 -3814 93174 25000
rect 93954 -1894 94574 25000
rect 94874 -7654 95494 25000
rect 96274 -5734 96894 25000
rect 97674 -3814 98294 25000
rect 99074 -1894 99694 25000
rect 99994 -7654 100614 25000
rect 101394 -5734 102014 25000
rect 102794 -3814 103414 25000
rect 104194 -1894 104814 25000
rect 105114 -7654 105734 25000
rect 106514 -5734 107134 25000
rect 107914 -3814 108534 25000
rect 109314 -1894 109934 25000
rect 110234 -7654 110854 25000
rect 111634 -5734 112254 25000
rect 113034 -3814 113654 25000
rect 114434 -1894 115054 25000
rect 115354 -7654 115974 25000
rect 116754 -5734 117374 25000
rect 118154 -3814 118774 25000
rect 119554 -1894 120174 25000
rect 120474 -7654 121094 25000
rect 121874 -5734 122494 25000
rect 123274 -3814 123894 25000
rect 124674 -1894 125294 25000
rect 125594 -7654 126214 25000
rect 126994 -5734 127614 25000
rect 128394 -3814 129014 25000
rect 129794 -1894 130414 25000
rect 130714 -7654 131334 25000
rect 132114 -5734 132734 25000
rect 133514 -3814 134134 25000
rect 134914 -1894 135534 25000
rect 135834 -7654 136454 25000
rect 137234 -5734 137854 25000
rect 138634 -3814 139254 25000
rect 140034 -1894 140654 25000
rect 140954 -7654 141574 25000
rect 142354 -5734 142974 25000
rect 143754 -3814 144374 25000
rect 145154 -1894 145774 25000
rect 146074 -7654 146694 25000
rect 147474 -5734 148094 25000
rect 148874 -3814 149494 25000
rect 150274 -1894 150894 25000
rect 151194 -7654 151814 25000
rect 152594 -5734 153214 25000
rect 153994 -3814 154614 25000
rect 155394 -1894 156014 25000
rect 156314 -7654 156934 25000
rect 157714 -5734 158334 25000
rect 159114 -3814 159734 25000
rect 160514 -1894 161134 25000
rect 161434 -7654 162054 25000
rect 162834 -5734 163454 25000
rect 164234 -3814 164854 25000
rect 165634 -1894 166254 25000
rect 166554 -7654 167174 25000
rect 167954 -5734 168574 25000
rect 169354 -3814 169974 25000
rect 170754 -1894 171374 25000
rect 171674 -7654 172294 25000
rect 173074 -5734 173694 25000
rect 174474 -3814 175094 25000
rect 175874 -1894 176494 25000
rect 176794 -7654 177414 25000
rect 178194 -5734 178814 25000
rect 179594 -3814 180214 25000
rect 180994 -1894 181614 25000
rect 181914 -7654 182534 25000
rect 183314 -5734 183934 25000
rect 184714 -3814 185334 25000
rect 186114 -1894 186734 25000
rect 187034 -7654 187654 25000
rect 188434 -5734 189054 25000
rect 189834 -3814 190454 25000
rect 191234 -1894 191854 25000
rect 192154 -7654 192774 25000
rect 193554 -5734 194174 25000
rect 194954 -3814 195574 25000
rect 196354 -1894 196974 25000
rect 197274 -7654 197894 25000
rect 198674 -5734 199294 25000
rect 200074 -3814 200694 25000
rect 201474 -1894 202094 25000
rect 202394 -7654 203014 25000
rect 203794 -5734 204414 25000
rect 205194 -3814 205814 25000
rect 206594 -1894 207214 25000
rect 207514 -7654 208134 25000
rect 208914 -5734 209534 25000
rect 210314 -3814 210934 25000
rect 211714 -1894 212334 25000
rect 212634 -7654 213254 25000
rect 214034 -5734 214654 25000
rect 215434 -3814 216054 25000
rect 216834 -1894 217454 25000
rect 217754 -7654 218374 25000
rect 219154 -5734 219774 25000
rect 220554 -3814 221174 25000
rect 221954 -1894 222574 25000
rect 222874 -7654 223494 25000
rect 224274 -5734 224894 25000
rect 225674 -3814 226294 25000
rect 227074 -1894 227694 25000
rect 227994 -7654 228614 25000
rect 229394 -5734 230014 25000
rect 230794 -3814 231414 25000
rect 232194 -1894 232814 25000
rect 233114 -7654 233734 25000
rect 234514 -5734 235134 25000
rect 235914 -3814 236534 25000
rect 237314 -1894 237934 25000
rect 238234 -7654 238854 25000
rect 239634 -5734 240254 25000
rect 241034 -3814 241654 25000
rect 242434 -1894 243054 25000
rect 243354 -7654 243974 25000
rect 244754 -5734 245374 25000
rect 246154 -3814 246774 25000
rect 247554 -1894 248174 25000
rect 248474 -7654 249094 25000
rect 249874 -5734 250494 25000
rect 251274 -3814 251894 25000
rect 252674 -1894 253294 25000
rect 253594 -7654 254214 25000
rect 254994 -5734 255614 25000
rect 256394 -3814 257014 25000
rect 257794 -1894 258414 25000
rect 258714 -7654 259334 25000
rect 260114 -5734 260734 25000
rect 261514 -3814 262134 25000
rect 262914 -1894 263534 25000
rect 263834 -7654 264454 25000
rect 265234 -5734 265854 25000
rect 266634 -3814 267254 25000
rect 268034 -1894 268654 25000
rect 268954 -7654 269574 25000
rect 270354 -5734 270974 25000
rect 271754 -3814 272374 25000
rect 273154 -1894 273774 25000
rect 274074 -7654 274694 25000
rect 275474 -5734 276094 25000
rect 276874 -3814 277494 25000
rect 278274 -1894 278894 25000
rect 279194 -7654 279814 25000
rect 280594 -5734 281214 25000
rect 281994 -3814 282614 25000
rect 283394 -1894 284014 25000
rect 284314 -7654 284934 25000
rect 285714 -5734 286334 25000
rect 287114 -3814 287734 25000
rect 288514 -1894 289134 25000
rect 289434 -7654 290054 25000
rect 290834 -5734 291454 25000
rect 292234 -3814 292854 25000
rect 293634 -1894 294254 25000
rect 294554 -7654 295174 25000
rect 295954 -5734 296574 25000
rect 297354 -3814 297974 25000
rect 298754 -1894 299374 25000
rect 299674 -7654 300294 25000
rect 301074 -5734 301694 25000
rect 302474 -3814 303094 25000
rect 303874 -1894 304494 25000
rect 304794 -7654 305414 25000
rect 306194 -5734 306814 25000
rect 307594 -3814 308214 25000
rect 308994 -1894 309614 25000
rect 309914 -7654 310534 25000
rect 311314 -5734 311934 25000
rect 312714 -3814 313334 25000
rect 314114 -1894 314734 25000
rect 315034 -7654 315654 25000
rect 316434 -5734 317054 25000
rect 317834 -3814 318454 25000
rect 319234 -1894 319854 25000
rect 320154 -7654 320774 25000
rect 321554 -5734 322174 25000
rect 322954 -3814 323574 25000
rect 324354 -1894 324974 25000
rect 325274 -7654 325894 25000
rect 326674 -5734 327294 25000
rect 328074 -3814 328694 25000
rect 329474 -1894 330094 25000
rect 330394 -7654 331014 25000
rect 331794 -5734 332414 25000
rect 333194 -3814 333814 25000
rect 334594 -1894 335214 25000
rect 335514 -7654 336134 25000
rect 336914 -5734 337534 25000
rect 338314 -3814 338934 25000
rect 339714 -1894 340334 25000
rect 340634 -7654 341254 25000
rect 342034 -5734 342654 25000
rect 343434 -3814 344054 25000
rect 344834 -1894 345454 25000
rect 345754 -7654 346374 25000
rect 347154 -5734 347774 25000
rect 348554 -3814 349174 25000
rect 349954 -1894 350574 25000
rect 350874 -7654 351494 25000
rect 352274 -5734 352894 25000
rect 353674 -3814 354294 25000
rect 355074 -1894 355694 25000
rect 355994 -7654 356614 25000
rect 357394 -5734 358014 25000
rect 358794 -3814 359414 25000
rect 360194 -1894 360814 25000
rect 361114 -7654 361734 25000
rect 362514 -5734 363134 25000
rect 363914 -3814 364534 25000
rect 365314 -1894 365934 25000
rect 366234 -7654 366854 25000
rect 367634 -5734 368254 25000
rect 369034 -3814 369654 25000
rect 370434 -1894 371054 25000
rect 371354 -7654 371974 25000
rect 372754 -5734 373374 25000
rect 374154 -3814 374774 25000
rect 375554 -1894 376174 25000
rect 376474 -7654 377094 25000
rect 377874 -5734 378494 25000
rect 379274 -3814 379894 25000
rect 380674 -1894 381294 25000
rect 381594 -7654 382214 25000
rect 382994 -5734 383614 25000
rect 384394 -3814 385014 25000
rect 385794 -1894 386414 25000
rect 386714 -7654 387334 25000
rect 388114 -5734 388734 25000
rect 389514 -3814 390134 25000
rect 390914 -1894 391534 25000
rect 391834 -7654 392454 25000
rect 393234 -5734 393854 25000
rect 394634 -3814 395254 25000
rect 396034 -1894 396654 25000
rect 396954 -7654 397574 25000
rect 398354 -5734 398974 25000
rect 399754 -3814 400374 25000
rect 401154 -1894 401774 25000
rect 402074 -7654 402694 25000
rect 403474 -5734 404094 25000
rect 404874 -3814 405494 25000
rect 406274 -1894 406894 25000
rect 407194 -7654 407814 25000
rect 408594 -5734 409214 25000
rect 409994 -3814 410614 25000
rect 411394 -1894 412014 25000
rect 412314 -7654 412934 25000
rect 413714 -5734 414334 25000
rect 415114 -3814 415734 25000
rect 416514 -1894 417134 25000
rect 417434 -7654 418054 25000
rect 418834 -5734 419454 25000
rect 420234 -3814 420854 25000
rect 421634 -1894 422254 25000
rect 422554 -7654 423174 25000
rect 423954 -5734 424574 25000
rect 425354 -3814 425974 25000
rect 426754 -1894 427374 25000
rect 427674 -7654 428294 25000
rect 429074 -5734 429694 25000
rect 430474 -3814 431094 25000
rect 431874 -1894 432494 25000
rect 432794 -7654 433414 25000
rect 434194 -5734 434814 25000
rect 435594 -3814 436214 25000
rect 436994 -1894 437614 25000
rect 437914 -7654 438534 25000
rect 439314 -5734 439934 25000
rect 440714 -3814 441334 25000
rect 442114 -1894 442734 25000
rect 443034 -7654 443654 25000
rect 444434 -5734 445054 25000
rect 445834 -3814 446454 25000
rect 447234 -1894 447854 25000
rect 448154 -7654 448774 25000
rect 449554 -5734 450174 25000
rect 450954 -3814 451574 25000
rect 452354 -1894 452974 25000
rect 453274 -7654 453894 25000
rect 454674 -5734 455294 25000
rect 456074 -3814 456694 25000
rect 457474 -1894 458094 25000
rect 458394 -7654 459014 25000
rect 459794 -5734 460414 25000
rect 461194 -3814 461814 25000
rect 462594 -1894 463214 25000
rect 463514 -7654 464134 25000
rect 464914 -5734 465534 25000
rect 466314 -3814 466934 25000
rect 467714 -1894 468334 25000
rect 468634 -7654 469254 25000
rect 470034 -5734 470654 25000
rect 471434 -3814 472054 25000
rect 472834 -1894 473454 25000
rect 473754 -7654 474374 25000
rect 475154 -5734 475774 25000
rect 476554 -3814 477174 25000
rect 477954 -1894 478574 25000
rect 478874 -7654 479494 25000
rect 480274 -5734 480894 25000
rect 481674 -3814 482294 25000
rect 483074 -1894 483694 25000
rect 483994 -7654 484614 25000
rect 485394 -5734 486014 25000
rect 486794 -3814 487414 25000
rect 488194 -1894 488814 25000
rect 489114 -7654 489734 25000
rect 490514 -5734 491134 25000
rect 491914 -3814 492534 25000
rect 493314 -1894 493934 25000
rect 494234 -7654 494854 25000
rect 495634 -5734 496254 25000
rect 497034 -3814 497654 25000
rect 498434 -1894 499054 25000
rect 499354 -7654 499974 25000
rect 500754 -5734 501374 25000
rect 502154 -3814 502774 25000
rect 503554 -1894 504174 25000
rect 504474 -7654 505094 25000
rect 505874 -5734 506494 25000
rect 507274 -3814 507894 25000
rect 508674 -1894 509294 25000
rect 509594 -7654 510214 25000
rect 510994 -5734 511614 25000
rect 512394 -3814 513014 25000
rect 513794 -1894 514414 25000
rect 514714 -7654 515334 25000
rect 516114 -5734 516734 25000
rect 517514 -3814 518134 25000
rect 518914 -1894 519534 25000
rect 519834 -7654 520454 25000
rect 521234 -5734 521854 25000
rect 522634 -3814 523254 25000
rect 524034 -1894 524654 25000
rect 524954 -7654 525574 25000
rect 526354 -5734 526974 25000
rect 527754 -3814 528374 25000
rect 529154 -1894 529774 25000
rect 530074 -7654 530694 25000
rect 531474 -5734 532094 25000
rect 532874 -3814 533494 25000
rect 534274 -1894 534894 25000
rect 535194 -7654 535814 25000
rect 536594 -5734 537214 25000
rect 537994 -3814 538614 25000
rect 539394 -1894 540014 25000
rect 540314 -7654 540934 25000
rect 541714 -5734 542334 25000
rect 543114 -3814 543734 25000
rect 544514 -1894 545134 25000
rect 545434 -7654 546054 25000
rect 546834 -5734 547454 25000
rect 548234 -3814 548854 25000
rect 549634 -1894 550254 25000
rect 550554 -7654 551174 25000
rect 551954 -5734 552574 709670
rect 553354 -3814 553974 707750
rect 554754 -1894 555374 705830
rect 555674 -7654 556294 711590
rect 557074 -5734 557694 709670
rect 558474 -3814 559094 707750
rect 559874 -1894 560494 705830
rect 560794 -7654 561414 711590
rect 562194 -5734 562814 709670
rect 563594 -3814 564214 707750
rect 564994 -1894 565614 705830
rect 565914 -7654 566534 711590
rect 567314 -5734 567934 709670
rect 568714 -3814 569334 707750
rect 570114 -1894 570734 705830
rect 571034 -7654 571654 711590
rect 572434 -5734 573054 709670
rect 573834 -3814 574454 707750
rect 575234 -1894 575854 705830
rect 576154 -7654 576774 711590
rect 577554 -5734 578174 709670
rect 578954 -3814 579574 707750
rect 580354 -1894 580974 705830
rect 581274 -7654 581894 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 33243 29128 546669 664616
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -6806 694306 590730 694926
rect -4886 690586 588810 691206
rect -2966 686866 586890 687486
rect -8726 680026 592650 680646
rect -6806 676306 590730 676926
rect -4886 672586 588810 673206
rect -2966 668866 586890 669486
rect -8726 662026 592650 662646
rect -6806 658306 590730 658926
rect -4886 654586 588810 655206
rect -2966 650866 586890 651486
rect -8726 644026 592650 644646
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -2966 632866 586890 633486
rect -8726 626026 592650 626646
rect -6806 622306 590730 622926
rect -4886 618586 588810 619206
rect -2966 614866 586890 615486
rect -8726 608026 592650 608646
rect -6806 604306 590730 604926
rect -4886 600586 588810 601206
rect -2966 596866 586890 597486
rect -8726 590026 592650 590646
rect -6806 586306 590730 586926
rect -4886 582586 588810 583206
rect -2966 578866 586890 579486
rect -8726 572026 592650 572646
rect -6806 568306 590730 568926
rect -4886 564586 588810 565206
rect -2966 560866 586890 561486
rect -8726 554026 592650 554646
rect -6806 550306 590730 550926
rect -4886 546586 588810 547206
rect -2966 542866 586890 543486
rect -8726 536026 592650 536646
rect -6806 532306 590730 532926
rect -4886 528586 588810 529206
rect -2966 524866 586890 525486
rect -8726 518026 592650 518646
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -2966 506866 586890 507486
rect -8726 500026 592650 500646
rect -6806 496306 590730 496926
rect -4886 492586 588810 493206
rect -2966 488866 586890 489486
rect -8726 482026 592650 482646
rect -6806 478306 590730 478926
rect -4886 474586 588810 475206
rect -2966 470866 586890 471486
rect -8726 464026 592650 464646
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -2966 452866 586890 453486
rect -8726 446026 592650 446646
rect -6806 442306 590730 442926
rect -4886 438586 588810 439206
rect -2966 434866 586890 435486
rect -8726 428026 592650 428646
rect -6806 424306 590730 424926
rect -4886 420586 588810 421206
rect -2966 416866 586890 417486
rect -8726 410026 592650 410646
rect -6806 406306 590730 406926
rect -4886 402586 588810 403206
rect -2966 398866 586890 399486
rect -8726 392026 592650 392646
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -2966 380866 586890 381486
rect -8726 374026 592650 374646
rect -6806 370306 590730 370926
rect -4886 366586 588810 367206
rect -2966 362866 586890 363486
rect -8726 356026 592650 356646
rect -6806 352306 590730 352926
rect -4886 348586 588810 349206
rect -2966 344866 586890 345486
rect -8726 338026 592650 338646
rect -6806 334306 590730 334926
rect -4886 330586 588810 331206
rect -2966 326866 586890 327486
rect -8726 320026 592650 320646
rect -6806 316306 590730 316926
rect -4886 312586 588810 313206
rect -2966 308866 586890 309486
rect -8726 302026 592650 302646
rect -6806 298306 590730 298926
rect -4886 294586 588810 295206
rect -2966 290866 586890 291486
rect -8726 284026 592650 284646
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -2966 272866 586890 273486
rect -8726 266026 592650 266646
rect -6806 262306 590730 262926
rect -4886 258586 588810 259206
rect -2966 254866 586890 255486
rect -8726 248026 592650 248646
rect -6806 244306 590730 244926
rect -4886 240586 588810 241206
rect -2966 236866 586890 237486
rect -8726 230026 592650 230646
rect -6806 226306 590730 226926
rect -4886 222586 588810 223206
rect -2966 218866 586890 219486
rect -8726 212026 592650 212646
rect -6806 208306 590730 208926
rect -4886 204586 588810 205206
rect -2966 200866 586890 201486
rect -8726 194026 592650 194646
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -2966 182866 586890 183486
rect -8726 176026 592650 176646
rect -6806 172306 590730 172926
rect -4886 168586 588810 169206
rect -2966 164866 586890 165486
rect -8726 158026 592650 158646
rect -6806 154306 590730 154926
rect -4886 150586 588810 151206
rect -2966 146866 586890 147486
rect -8726 140026 592650 140646
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -2966 128866 586890 129486
rect -8726 122026 592650 122646
rect -6806 118306 590730 118926
rect -4886 114586 588810 115206
rect -2966 110866 586890 111486
rect -8726 104026 592650 104646
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -2966 92866 586890 93486
rect -8726 86026 592650 86646
rect -6806 82306 590730 82926
rect -4886 78586 588810 79206
rect -2966 74866 586890 75486
rect -8726 68026 592650 68646
rect -6806 64306 590730 64926
rect -4886 60586 588810 61206
rect -2966 56866 586890 57486
rect -8726 50026 592650 50646
rect -6806 46306 590730 46926
rect -4886 42586 588810 43206
rect -2966 38866 586890 39486
rect -8726 32026 592650 32646
rect -6806 28306 590730 28926
rect -4886 24586 588810 25206
rect -2966 20866 586890 21486
rect -8726 14026 592650 14646
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 32514 -1894 33134 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 42754 -1894 43374 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 52994 -1894 53614 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 63234 -1894 63854 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73474 -1894 74094 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 83714 -1894 84334 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 93954 -1894 94574 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 104194 -1894 104814 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 114434 -1894 115054 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 124674 -1894 125294 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 134914 -1894 135534 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145154 -1894 145774 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 155394 -1894 156014 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 165634 -1894 166254 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 175874 -1894 176494 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 186114 -1894 186734 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 196354 -1894 196974 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 206594 -1894 207214 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 216834 -1894 217454 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 227074 -1894 227694 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 237314 -1894 237934 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 247554 -1894 248174 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 257794 -1894 258414 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 268034 -1894 268654 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 278274 -1894 278894 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 288514 -1894 289134 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 298754 -1894 299374 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 308994 -1894 309614 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 319234 -1894 319854 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 329474 -1894 330094 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 339714 -1894 340334 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 349954 -1894 350574 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 360194 -1894 360814 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 370434 -1894 371054 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 380674 -1894 381294 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 390914 -1894 391534 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 401154 -1894 401774 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 411394 -1894 412014 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 421634 -1894 422254 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 431874 -1894 432494 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 442114 -1894 442734 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 452354 -1894 452974 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 462594 -1894 463214 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 472834 -1894 473454 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 483074 -1894 483694 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 493314 -1894 493934 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 503554 -1894 504174 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 513794 -1894 514414 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 524034 -1894 524654 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 534274 -1894 534894 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s 544514 -1894 545134 25000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 12034 -1894 12654 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 22274 -1894 22894 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 32514 669000 33134 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 42754 669000 43374 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 52994 669000 53614 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 63234 669000 63854 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 73474 669000 74094 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 83714 669000 84334 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 93954 669000 94574 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 104194 669000 104814 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 114434 669000 115054 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 124674 669000 125294 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 134914 669000 135534 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 145154 669000 145774 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 155394 669000 156014 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 165634 669000 166254 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 175874 669000 176494 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 186114 669000 186734 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 196354 669000 196974 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 206594 669000 207214 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 216834 669000 217454 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 227074 669000 227694 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 237314 669000 237934 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 247554 669000 248174 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 257794 669000 258414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 268034 669000 268654 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 278274 669000 278894 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 288514 669000 289134 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 298754 669000 299374 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 308994 669000 309614 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 319234 669000 319854 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 329474 669000 330094 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 339714 669000 340334 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 349954 669000 350574 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 360194 669000 360814 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 370434 669000 371054 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 380674 669000 381294 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 390914 669000 391534 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 401154 669000 401774 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 411394 669000 412014 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 421634 669000 422254 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 431874 669000 432494 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 442114 669000 442734 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 452354 669000 452974 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 462594 669000 463214 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 472834 669000 473454 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 483074 669000 483694 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 493314 669000 493934 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 503554 669000 504174 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 513794 669000 514414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 524034 669000 524654 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 534274 669000 534894 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 544514 669000 545134 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 554754 -1894 555374 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 564994 -1894 565614 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 575234 -1894 575854 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 36234 -3814 36854 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 46474 -3814 47094 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 56714 -3814 57334 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 66954 -3814 67574 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 77194 -3814 77814 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 87434 -3814 88054 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 97674 -3814 98294 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 107914 -3814 108534 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 118154 -3814 118774 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 128394 -3814 129014 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 138634 -3814 139254 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 148874 -3814 149494 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 159114 -3814 159734 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 169354 -3814 169974 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 179594 -3814 180214 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 189834 -3814 190454 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 200074 -3814 200694 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 210314 -3814 210934 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 220554 -3814 221174 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 230794 -3814 231414 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 241034 -3814 241654 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 251274 -3814 251894 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 261514 -3814 262134 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 271754 -3814 272374 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 281994 -3814 282614 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 292234 -3814 292854 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 302474 -3814 303094 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 312714 -3814 313334 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 322954 -3814 323574 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 333194 -3814 333814 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 343434 -3814 344054 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 353674 -3814 354294 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 363914 -3814 364534 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 374154 -3814 374774 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 384394 -3814 385014 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 394634 -3814 395254 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 404874 -3814 405494 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 415114 -3814 415734 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 425354 -3814 425974 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 435594 -3814 436214 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 445834 -3814 446454 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 456074 -3814 456694 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 466314 -3814 466934 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 476554 -3814 477174 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 486794 -3814 487414 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 497034 -3814 497654 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 507274 -3814 507894 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 517514 -3814 518134 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 527754 -3814 528374 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 537994 -3814 538614 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s 548234 -3814 548854 25000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 15754 -3814 16374 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 25994 -3814 26614 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 36234 669000 36854 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 46474 669000 47094 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 56714 669000 57334 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 66954 669000 67574 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 77194 669000 77814 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 87434 669000 88054 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 97674 669000 98294 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 107914 669000 108534 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 118154 669000 118774 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 128394 669000 129014 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 138634 669000 139254 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 148874 669000 149494 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 159114 669000 159734 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 169354 669000 169974 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 179594 669000 180214 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 189834 669000 190454 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 200074 669000 200694 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 210314 669000 210934 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 220554 669000 221174 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 230794 669000 231414 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 241034 669000 241654 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 251274 669000 251894 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 261514 669000 262134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 271754 669000 272374 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 281994 669000 282614 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 292234 669000 292854 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 302474 669000 303094 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 312714 669000 313334 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 322954 669000 323574 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 333194 669000 333814 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 343434 669000 344054 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 353674 669000 354294 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 363914 669000 364534 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 374154 669000 374774 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 384394 669000 385014 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 394634 669000 395254 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 404874 669000 405494 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 415114 669000 415734 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 425354 669000 425974 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 435594 669000 436214 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 445834 669000 446454 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 456074 669000 456694 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 466314 669000 466934 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 476554 669000 477174 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 486794 669000 487414 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 497034 669000 497654 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 507274 669000 507894 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 517514 669000 518134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 527754 669000 528374 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 537994 669000 538614 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 548234 669000 548854 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 558474 -3814 559094 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 568714 -3814 569334 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 578954 -3814 579574 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 29714 -5734 30334 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 39954 -5734 40574 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 50194 -5734 50814 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 60434 -5734 61054 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 70674 -5734 71294 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 80914 -5734 81534 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 91154 -5734 91774 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 101394 -5734 102014 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 111634 -5734 112254 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 121874 -5734 122494 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 132114 -5734 132734 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 142354 -5734 142974 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 152594 -5734 153214 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 162834 -5734 163454 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 173074 -5734 173694 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 183314 -5734 183934 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 193554 -5734 194174 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 203794 -5734 204414 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 214034 -5734 214654 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 224274 -5734 224894 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 234514 -5734 235134 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 244754 -5734 245374 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 254994 -5734 255614 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 265234 -5734 265854 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 275474 -5734 276094 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 285714 -5734 286334 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 295954 -5734 296574 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 306194 -5734 306814 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 316434 -5734 317054 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 326674 -5734 327294 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 336914 -5734 337534 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 347154 -5734 347774 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 357394 -5734 358014 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 367634 -5734 368254 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 377874 -5734 378494 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 388114 -5734 388734 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 398354 -5734 398974 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 408594 -5734 409214 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 418834 -5734 419454 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 429074 -5734 429694 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 439314 -5734 439934 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 449554 -5734 450174 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 459794 -5734 460414 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 470034 -5734 470654 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 480274 -5734 480894 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 490514 -5734 491134 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 500754 -5734 501374 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 510994 -5734 511614 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 521234 -5734 521854 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 531474 -5734 532094 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s 541714 -5734 542334 25000 6 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 19474 -5734 20094 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 29714 669000 30334 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 39954 669000 40574 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 50194 669000 50814 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 60434 669000 61054 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 70674 669000 71294 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 80914 669000 81534 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 91154 669000 91774 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 101394 669000 102014 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 111634 669000 112254 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 121874 669000 122494 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 132114 669000 132734 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 142354 669000 142974 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 152594 669000 153214 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 162834 669000 163454 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 173074 669000 173694 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 183314 669000 183934 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 193554 669000 194174 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 203794 669000 204414 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 214034 669000 214654 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 224274 669000 224894 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 234514 669000 235134 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 244754 669000 245374 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 254994 669000 255614 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 265234 669000 265854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 275474 669000 276094 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 285714 669000 286334 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 295954 669000 296574 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 306194 669000 306814 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 316434 669000 317054 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 326674 669000 327294 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 336914 669000 337534 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 347154 669000 347774 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 357394 669000 358014 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 367634 669000 368254 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 377874 669000 378494 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 388114 669000 388734 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 398354 669000 398974 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 408594 669000 409214 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 418834 669000 419454 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 429074 669000 429694 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 439314 669000 439934 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 449554 669000 450174 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 459794 669000 460414 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 470034 669000 470654 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 480274 669000 480894 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 490514 669000 491134 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 500754 669000 501374 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 510994 669000 511614 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 521234 669000 521854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 531474 669000 532094 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 541714 669000 542334 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 551954 -5734 552574 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 562194 -5734 562814 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 572434 -5734 573054 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 33434 -7654 34054 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 43674 -7654 44294 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 53914 -7654 54534 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 64154 -7654 64774 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 74394 -7654 75014 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 84634 -7654 85254 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 94874 -7654 95494 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 105114 -7654 105734 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 115354 -7654 115974 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 125594 -7654 126214 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 135834 -7654 136454 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 146074 -7654 146694 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 156314 -7654 156934 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 166554 -7654 167174 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 176794 -7654 177414 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 187034 -7654 187654 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 197274 -7654 197894 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 207514 -7654 208134 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 217754 -7654 218374 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 227994 -7654 228614 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 238234 -7654 238854 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 248474 -7654 249094 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 258714 -7654 259334 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 268954 -7654 269574 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 279194 -7654 279814 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 289434 -7654 290054 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 299674 -7654 300294 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 309914 -7654 310534 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 320154 -7654 320774 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 330394 -7654 331014 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 340634 -7654 341254 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 350874 -7654 351494 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 361114 -7654 361734 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 371354 -7654 371974 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 381594 -7654 382214 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 391834 -7654 392454 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 402074 -7654 402694 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 412314 -7654 412934 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 422554 -7654 423174 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 432794 -7654 433414 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 443034 -7654 443654 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 453274 -7654 453894 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 463514 -7654 464134 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 473754 -7654 474374 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 483994 -7654 484614 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 494234 -7654 494854 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 504474 -7654 505094 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 514714 -7654 515334 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 524954 -7654 525574 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 535194 -7654 535814 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s 545434 -7654 546054 25000 6 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 23194 -7654 23814 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 33434 669000 34054 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 43674 669000 44294 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 53914 669000 54534 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 64154 669000 64774 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 74394 669000 75014 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 84634 669000 85254 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 94874 669000 95494 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 105114 669000 105734 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 115354 669000 115974 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 125594 669000 126214 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 135834 669000 136454 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 146074 669000 146694 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 156314 669000 156934 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 166554 669000 167174 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 176794 669000 177414 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 187034 669000 187654 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 197274 669000 197894 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 207514 669000 208134 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 217754 669000 218374 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 227994 669000 228614 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 238234 669000 238854 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 248474 669000 249094 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 258714 669000 259334 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 268954 669000 269574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 279194 669000 279814 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 289434 669000 290054 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 299674 669000 300294 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 309914 669000 310534 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 320154 669000 320774 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 330394 669000 331014 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 340634 669000 341254 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 350874 669000 351494 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 361114 669000 361734 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 371354 669000 371974 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 381594 669000 382214 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 391834 669000 392454 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 402074 669000 402694 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 412314 669000 412934 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 422554 669000 423174 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 432794 669000 433414 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 443034 669000 443654 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 453274 669000 453894 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 463514 669000 464134 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 473754 669000 474374 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 483994 669000 484614 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 494234 669000 494854 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 504474 669000 505094 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 514714 669000 515334 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 524954 669000 525574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 535194 669000 535814 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 545434 669000 546054 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 555674 -7654 556294 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 565914 -7654 566534 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 576154 -7654 576774 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 34834 -5734 35454 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 45074 -5734 45694 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 55314 -5734 55934 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 65554 -5734 66174 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 75794 -5734 76414 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 86034 -5734 86654 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 96274 -5734 96894 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 106514 -5734 107134 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 116754 -5734 117374 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 126994 -5734 127614 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 137234 -5734 137854 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 147474 -5734 148094 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 157714 -5734 158334 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 167954 -5734 168574 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 178194 -5734 178814 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 188434 -5734 189054 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 198674 -5734 199294 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 208914 -5734 209534 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219154 -5734 219774 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229394 -5734 230014 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239634 -5734 240254 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 249874 -5734 250494 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 260114 -5734 260734 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 270354 -5734 270974 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 280594 -5734 281214 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 290834 -5734 291454 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 301074 -5734 301694 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 311314 -5734 311934 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 321554 -5734 322174 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 331794 -5734 332414 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 342034 -5734 342654 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 352274 -5734 352894 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 362514 -5734 363134 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 372754 -5734 373374 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 382994 -5734 383614 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 393234 -5734 393854 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 403474 -5734 404094 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 413714 -5734 414334 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423954 -5734 424574 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 434194 -5734 434814 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 444434 -5734 445054 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 454674 -5734 455294 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 464914 -5734 465534 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 475154 -5734 475774 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 485394 -5734 486014 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495634 -5734 496254 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 505874 -5734 506494 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 516114 -5734 516734 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 526354 -5734 526974 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 536594 -5734 537214 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 546834 -5734 547454 25000 6 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 14354 -5734 14974 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 24594 -5734 25214 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 34834 669000 35454 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 45074 669000 45694 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 55314 669000 55934 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 65554 669000 66174 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 75794 669000 76414 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 86034 669000 86654 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 96274 669000 96894 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 106514 669000 107134 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 116754 669000 117374 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 126994 669000 127614 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 137234 669000 137854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 147474 669000 148094 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 157714 669000 158334 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 167954 669000 168574 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 178194 669000 178814 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 188434 669000 189054 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 198674 669000 199294 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 208914 669000 209534 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 219154 669000 219774 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229394 669000 230014 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 239634 669000 240254 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 249874 669000 250494 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 260114 669000 260734 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 270354 669000 270974 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 280594 669000 281214 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 290834 669000 291454 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 301074 669000 301694 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 311314 669000 311934 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 321554 669000 322174 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 331794 669000 332414 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 342034 669000 342654 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 352274 669000 352894 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 362514 669000 363134 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 372754 669000 373374 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 382994 669000 383614 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 393234 669000 393854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 403474 669000 404094 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 413714 669000 414334 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423954 669000 424574 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 434194 669000 434814 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 444434 669000 445054 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 454674 669000 455294 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 464914 669000 465534 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 475154 669000 475774 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 485394 669000 486014 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495634 669000 496254 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 505874 669000 506494 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 516114 669000 516734 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 526354 669000 526974 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 536594 669000 537214 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 546834 669000 547454 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 557074 -5734 557694 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 567314 -5734 567934 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 577554 -5734 578174 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 28314 -7654 28934 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 38554 -7654 39174 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 48794 -7654 49414 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 59034 -7654 59654 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 69274 -7654 69894 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 79514 -7654 80134 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 89754 -7654 90374 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 99994 -7654 100614 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110234 -7654 110854 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 120474 -7654 121094 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 130714 -7654 131334 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 140954 -7654 141574 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 151194 -7654 151814 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 161434 -7654 162054 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 171674 -7654 172294 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 181914 -7654 182534 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 192154 -7654 192774 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 202394 -7654 203014 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 212634 -7654 213254 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222874 -7654 223494 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233114 -7654 233734 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 243354 -7654 243974 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 253594 -7654 254214 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 263834 -7654 264454 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 274074 -7654 274694 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 284314 -7654 284934 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 294554 -7654 295174 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 304794 -7654 305414 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 315034 -7654 315654 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 325274 -7654 325894 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 335514 -7654 336134 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 345754 -7654 346374 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 355994 -7654 356614 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 366234 -7654 366854 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 376474 -7654 377094 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 386714 -7654 387334 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 396954 -7654 397574 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 407194 -7654 407814 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 417434 -7654 418054 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 427674 -7654 428294 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 437914 -7654 438534 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 448154 -7654 448774 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 458394 -7654 459014 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 468634 -7654 469254 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 478874 -7654 479494 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 489114 -7654 489734 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 499354 -7654 499974 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 509594 -7654 510214 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 519834 -7654 520454 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 530074 -7654 530694 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 540314 -7654 540934 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 550554 -7654 551174 25000 6 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 18074 -7654 18694 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 28314 669000 28934 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 38554 669000 39174 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 48794 669000 49414 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 59034 669000 59654 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 69274 669000 69894 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 79514 669000 80134 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 89754 669000 90374 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 99994 669000 100614 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 110234 669000 110854 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 120474 669000 121094 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 130714 669000 131334 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 140954 669000 141574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 151194 669000 151814 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 161434 669000 162054 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 171674 669000 172294 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 181914 669000 182534 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 192154 669000 192774 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 202394 669000 203014 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 212634 669000 213254 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 222874 669000 223494 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 233114 669000 233734 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 243354 669000 243974 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 253594 669000 254214 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 263834 669000 264454 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 274074 669000 274694 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 284314 669000 284934 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 294554 669000 295174 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 304794 669000 305414 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 315034 669000 315654 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 325274 669000 325894 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 335514 669000 336134 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 345754 669000 346374 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 355994 669000 356614 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 366234 669000 366854 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 376474 669000 377094 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 386714 669000 387334 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 396954 669000 397574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 407194 669000 407814 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 417434 669000 418054 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 427674 669000 428294 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 437914 669000 438534 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 448154 669000 448774 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 458394 669000 459014 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 468634 669000 469254 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 478874 669000 479494 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 489114 669000 489734 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 499354 669000 499974 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 509594 669000 510214 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 519834 669000 520454 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 530074 669000 530694 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 540314 669000 540934 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 550554 669000 551174 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 560794 -7654 561414 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 571034 -7654 571654 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 581274 -7654 581894 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 27394 -1894 28014 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 37634 -1894 38254 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 47874 -1894 48494 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 58114 -1894 58734 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 68354 -1894 68974 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 78594 -1894 79214 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 88834 -1894 89454 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99074 -1894 99694 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 109314 -1894 109934 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 119554 -1894 120174 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 129794 -1894 130414 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 140034 -1894 140654 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 150274 -1894 150894 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 160514 -1894 161134 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 170754 -1894 171374 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 180994 -1894 181614 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191234 -1894 191854 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 201474 -1894 202094 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211714 -1894 212334 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 221954 -1894 222574 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 232194 -1894 232814 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 242434 -1894 243054 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 252674 -1894 253294 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 262914 -1894 263534 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 273154 -1894 273774 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 283394 -1894 284014 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 293634 -1894 294254 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 303874 -1894 304494 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 314114 -1894 314734 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 324354 -1894 324974 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 334594 -1894 335214 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 344834 -1894 345454 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 355074 -1894 355694 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 365314 -1894 365934 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 375554 -1894 376174 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 385794 -1894 386414 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 396034 -1894 396654 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 406274 -1894 406894 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 416514 -1894 417134 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 426754 -1894 427374 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 436994 -1894 437614 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 447234 -1894 447854 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 457474 -1894 458094 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 467714 -1894 468334 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 477954 -1894 478574 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 488194 -1894 488814 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 498434 -1894 499054 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 508674 -1894 509294 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 518914 -1894 519534 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 529154 -1894 529774 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 539394 -1894 540014 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 549634 -1894 550254 25000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 6914 -1894 7534 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 17154 -1894 17774 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 27394 669000 28014 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 37634 669000 38254 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 47874 669000 48494 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 58114 669000 58734 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 68354 669000 68974 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 78594 669000 79214 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 88834 669000 89454 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99074 669000 99694 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 109314 669000 109934 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 119554 669000 120174 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 129794 669000 130414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 140034 669000 140654 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 150274 669000 150894 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 160514 669000 161134 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 170754 669000 171374 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 180994 669000 181614 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 191234 669000 191854 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 201474 669000 202094 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 211714 669000 212334 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 221954 669000 222574 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 232194 669000 232814 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 242434 669000 243054 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 252674 669000 253294 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 262914 669000 263534 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 273154 669000 273774 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 283394 669000 284014 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 293634 669000 294254 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 303874 669000 304494 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 314114 669000 314734 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 324354 669000 324974 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 334594 669000 335214 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 344834 669000 345454 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 355074 669000 355694 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 365314 669000 365934 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 375554 669000 376174 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 385794 669000 386414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 396034 669000 396654 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 406274 669000 406894 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 416514 669000 417134 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 426754 669000 427374 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 436994 669000 437614 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 447234 669000 447854 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 457474 669000 458094 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 467714 669000 468334 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 477954 669000 478574 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 488194 669000 488814 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 498434 669000 499054 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 508674 669000 509294 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 518914 669000 519534 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 529154 669000 529774 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 539394 669000 540014 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 549634 669000 550254 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 559874 -1894 560494 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 570114 -1894 570734 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 580354 -1894 580974 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 31114 -3814 31734 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 41354 -3814 41974 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 51594 -3814 52214 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 61834 -3814 62454 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 72074 -3814 72694 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 82314 -3814 82934 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 92554 -3814 93174 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 102794 -3814 103414 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 113034 -3814 113654 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 123274 -3814 123894 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 133514 -3814 134134 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 143754 -3814 144374 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 153994 -3814 154614 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 164234 -3814 164854 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 174474 -3814 175094 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 184714 -3814 185334 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 194954 -3814 195574 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 205194 -3814 205814 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215434 -3814 216054 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 225674 -3814 226294 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235914 -3814 236534 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 246154 -3814 246774 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 256394 -3814 257014 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 266634 -3814 267254 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 276874 -3814 277494 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 287114 -3814 287734 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 297354 -3814 297974 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 307594 -3814 308214 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 317834 -3814 318454 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 328074 -3814 328694 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 338314 -3814 338934 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 348554 -3814 349174 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 358794 -3814 359414 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 369034 -3814 369654 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 379274 -3814 379894 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 389514 -3814 390134 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 399754 -3814 400374 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 409994 -3814 410614 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 420234 -3814 420854 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 430474 -3814 431094 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 440714 -3814 441334 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 450954 -3814 451574 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 461194 -3814 461814 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 471434 -3814 472054 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 481674 -3814 482294 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491914 -3814 492534 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 502154 -3814 502774 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 512394 -3814 513014 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 522634 -3814 523254 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 532874 -3814 533494 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 543114 -3814 543734 25000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 10634 -3814 11254 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 20874 -3814 21494 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 31114 669000 31734 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 41354 669000 41974 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 51594 669000 52214 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 61834 669000 62454 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 72074 669000 72694 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 82314 669000 82934 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 92554 669000 93174 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 102794 669000 103414 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 113034 669000 113654 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 123274 669000 123894 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 133514 669000 134134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 143754 669000 144374 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 153994 669000 154614 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 164234 669000 164854 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 174474 669000 175094 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 184714 669000 185334 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 194954 669000 195574 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 205194 669000 205814 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 215434 669000 216054 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 225674 669000 226294 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 235914 669000 236534 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 246154 669000 246774 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 256394 669000 257014 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 266634 669000 267254 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 276874 669000 277494 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 287114 669000 287734 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 297354 669000 297974 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 307594 669000 308214 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 317834 669000 318454 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 328074 669000 328694 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 338314 669000 338934 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 348554 669000 349174 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 358794 669000 359414 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 369034 669000 369654 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 379274 669000 379894 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 389514 669000 390134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 399754 669000 400374 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 409994 669000 410614 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 420234 669000 420854 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 430474 669000 431094 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 440714 669000 441334 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 450954 669000 451574 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 461194 669000 461814 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 471434 669000 472054 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 481674 669000 482294 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491914 669000 492534 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 502154 669000 502774 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 512394 669000 513014 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 522634 669000 523254 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 532874 669000 533494 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 543114 669000 543734 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 553354 -3814 553974 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 563594 -3814 564214 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 573834 -3814 574454 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 404076908
string GDS_FILE /home/angl/mpw6-prga/caravel/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 402623422
<< end >>

