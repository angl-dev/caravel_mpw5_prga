VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 2934.450 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 194.330 2934.450 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 374.330 2934.450 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 554.330 2934.450 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 734.330 2934.450 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 914.330 2934.450 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1094.330 2934.450 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1274.330 2934.450 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1454.330 2934.450 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1634.330 2934.450 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1814.330 2934.450 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1994.330 2934.450 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2174.330 2934.450 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2354.330 2934.450 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2534.330 2934.450 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2714.330 2934.450 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2894.330 2934.450 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3074.330 2934.450 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3254.330 2934.450 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3434.330 2934.450 3437.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 162.570 -9.470 165.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.770 -9.470 216.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.970 -9.470 268.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 -9.470 319.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 367.370 -9.470 370.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 418.570 -9.470 421.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.770 -9.470 472.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 520.970 -9.470 524.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 572.170 -9.470 575.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.370 -9.470 626.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.570 -9.470 677.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.770 -9.470 728.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 776.970 -9.470 780.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 828.170 -9.470 831.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 879.370 -9.470 882.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 930.570 -9.470 933.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.770 -9.470 984.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.970 -9.470 1036.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.170 -9.470 1087.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.370 -9.470 1138.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1186.570 -9.470 1189.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1237.770 -9.470 1240.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1288.970 -9.470 1292.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1340.170 -9.470 1343.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1391.370 -9.470 1394.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.570 -9.470 1445.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.770 -9.470 1496.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.970 -9.470 1548.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1596.170 -9.470 1599.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.370 -9.470 1650.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1698.570 -9.470 1701.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1749.770 -9.470 1752.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1800.970 -9.470 1804.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1852.170 -9.470 1855.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1903.370 -9.470 1906.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.570 -9.470 1957.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2005.770 -9.470 2008.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.970 -9.470 2060.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.170 -9.470 2111.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2159.370 -9.470 2162.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2210.570 -9.470 2213.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2261.770 -9.470 2264.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2312.970 -9.470 2316.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2364.170 -9.470 2367.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2415.370 -9.470 2418.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2466.570 -9.470 2469.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2517.770 -9.470 2520.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2568.970 -9.470 2572.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2620.170 -9.470 2623.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2671.370 -9.470 2674.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2722.570 -9.470 2725.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.170 -9.470 63.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.370 -9.470 114.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 162.570 3345.000 165.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.770 3345.000 216.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.970 3345.000 268.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 3345.000 319.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 367.370 3345.000 370.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 418.570 3345.000 421.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.770 3345.000 472.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 520.970 3345.000 524.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 572.170 3345.000 575.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.370 3345.000 626.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.570 3345.000 677.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.770 3345.000 728.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 776.970 3345.000 780.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 828.170 3345.000 831.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 879.370 3345.000 882.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 930.570 3345.000 933.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.770 3345.000 984.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.970 3345.000 1036.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.170 3345.000 1087.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.370 3345.000 1138.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1186.570 3345.000 1189.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1237.770 3345.000 1240.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1288.970 3345.000 1292.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1340.170 3345.000 1343.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1391.370 3345.000 1394.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.570 3345.000 1445.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.770 3345.000 1496.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.970 3345.000 1548.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1596.170 3345.000 1599.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.370 3345.000 1650.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1698.570 3345.000 1701.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1749.770 3345.000 1752.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1800.970 3345.000 1804.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1852.170 3345.000 1855.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1903.370 3345.000 1906.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.570 3345.000 1957.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2005.770 3345.000 2008.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.970 3345.000 2060.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.170 3345.000 2111.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2159.370 3345.000 2162.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2210.570 3345.000 2213.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2261.770 3345.000 2264.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2312.970 3345.000 2316.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2364.170 3345.000 2367.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2415.370 3345.000 2418.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2466.570 3345.000 2469.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2517.770 3345.000 2520.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2568.970 3345.000 2572.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2620.170 3345.000 2623.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2671.370 3345.000 2674.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2722.570 3345.000 2725.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2773.770 -9.470 2776.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2824.970 -9.470 2828.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2876.170 -9.470 2879.270 3529.150 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 32.930 2944.050 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 212.930 2944.050 216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 392.930 2944.050 396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 572.930 2944.050 576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 752.930 2944.050 756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 932.930 2944.050 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.170 -19.070 184.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.370 -19.070 235.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 283.570 -19.070 286.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 -19.070 337.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 385.970 -19.070 389.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 437.170 -19.070 440.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.370 -19.070 491.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 539.570 -19.070 542.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 590.770 -19.070 593.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 641.970 -19.070 645.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.170 -19.070 696.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.370 -19.070 747.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 795.570 -19.070 798.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.770 -19.070 849.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 897.970 -19.070 901.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 949.170 -19.070 952.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1000.370 -19.070 1003.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1051.570 -19.070 1054.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1102.770 -19.070 1105.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1153.970 -19.070 1157.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1205.170 -19.070 1208.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.370 -19.070 1259.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1307.570 -19.070 1310.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.770 -19.070 1361.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1409.970 -19.070 1413.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1461.170 -19.070 1464.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1512.370 -19.070 1515.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1563.570 -19.070 1566.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.770 -19.070 1617.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1665.970 -19.070 1669.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1717.170 -19.070 1720.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.370 -19.070 1771.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1819.570 -19.070 1822.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1870.770 -19.070 1873.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.970 -19.070 1925.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1973.170 -19.070 1976.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.370 -19.070 2027.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.570 -19.070 2078.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2126.770 -19.070 2129.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.970 -19.070 2181.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2229.170 -19.070 2232.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.370 -19.070 2283.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2331.570 -19.070 2334.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2382.770 -19.070 2385.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2433.970 -19.070 2437.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2485.170 -19.070 2488.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.370 -19.070 2539.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2587.570 -19.070 2590.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2638.770 -19.070 2641.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2689.970 -19.070 2693.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2741.170 -19.070 2744.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.770 -19.070 81.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.970 -19.070 133.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.170 3345.000 184.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.370 3345.000 235.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 283.570 3345.000 286.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 3345.000 337.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 385.970 3345.000 389.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 437.170 3345.000 440.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.370 3345.000 491.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 539.570 3345.000 542.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 590.770 3345.000 593.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 641.970 3345.000 645.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.170 3345.000 696.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.370 3345.000 747.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 795.570 3345.000 798.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.770 3345.000 849.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 897.970 3345.000 901.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 949.170 3345.000 952.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1000.370 3345.000 1003.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1051.570 3345.000 1054.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1102.770 3345.000 1105.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1153.970 3345.000 1157.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1205.170 3345.000 1208.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.370 3345.000 1259.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1307.570 3345.000 1310.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.770 3345.000 1361.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1409.970 3345.000 1413.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1461.170 3345.000 1464.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1512.370 3345.000 1515.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1563.570 3345.000 1566.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.770 3345.000 1617.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1665.970 3345.000 1669.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1717.170 3345.000 1720.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.370 3345.000 1771.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1819.570 3345.000 1822.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1870.770 3345.000 1873.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.970 3345.000 1925.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1973.170 3345.000 1976.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.370 3345.000 2027.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.570 3345.000 2078.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2126.770 3345.000 2129.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.970 3345.000 2181.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2229.170 3345.000 2232.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.370 3345.000 2283.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2331.570 3345.000 2334.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2382.770 3345.000 2385.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2433.970 3345.000 2437.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2485.170 3345.000 2488.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.370 3345.000 2539.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2587.570 3345.000 2590.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2638.770 3345.000 2641.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2689.970 3345.000 2693.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2741.170 3345.000 2744.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2792.370 -19.070 2795.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2843.570 -19.070 2846.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2894.770 -19.070 2897.870 3538.750 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 51.530 2953.650 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 231.530 2953.650 234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 411.530 2953.650 414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 591.530 2953.650 594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 771.530 2953.650 774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 951.530 2953.650 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 148.570 -28.670 151.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 199.770 -28.670 202.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.970 -28.670 254.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 302.170 -28.670 305.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 353.370 -28.670 356.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.570 -28.670 407.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 455.770 -28.670 458.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 506.970 -28.670 510.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.170 -28.670 561.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 609.370 -28.670 612.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 660.570 -28.670 663.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.770 -28.670 714.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 762.970 -28.670 766.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.170 -28.670 817.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.370 -28.670 868.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 916.570 -28.670 919.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 967.770 -28.670 970.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1018.970 -28.670 1022.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1070.170 -28.670 1073.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.370 -28.670 1124.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1172.570 -28.670 1175.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.770 -28.670 1226.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1274.970 -28.670 1278.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.170 -28.670 1329.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.370 -28.670 1380.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1428.570 -28.670 1431.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1479.770 -28.670 1482.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1530.970 -28.670 1534.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1582.170 -28.670 1585.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.370 -28.670 1636.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.570 -28.670 1687.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.770 -28.670 1738.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.970 -28.670 1790.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1838.170 -28.670 1841.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1889.370 -28.670 1892.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1940.570 -28.670 1943.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.770 -28.670 1994.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2042.970 -28.670 2046.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.170 -28.670 2097.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.370 -28.670 2148.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2196.570 -28.670 2199.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2247.770 -28.670 2250.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2298.970 -28.670 2302.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2350.170 -28.670 2353.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.370 -28.670 2404.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2452.570 -28.670 2455.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2503.770 -28.670 2506.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.970 -28.670 2558.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2606.170 -28.670 2609.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2657.370 -28.670 2660.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.570 -28.670 2711.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.370 -28.670 100.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 148.570 3345.000 151.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 199.770 3345.000 202.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.970 3345.000 254.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 302.170 3345.000 305.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 353.370 3345.000 356.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.570 3345.000 407.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 455.770 3345.000 458.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 506.970 3345.000 510.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.170 3345.000 561.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 609.370 3345.000 612.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 660.570 3345.000 663.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.770 3345.000 714.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 762.970 3345.000 766.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.170 3345.000 817.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.370 3345.000 868.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 916.570 3345.000 919.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 967.770 3345.000 970.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1018.970 3345.000 1022.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1070.170 3345.000 1073.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.370 3345.000 1124.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1172.570 3345.000 1175.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.770 3345.000 1226.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1274.970 3345.000 1278.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.170 3345.000 1329.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.370 3345.000 1380.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1428.570 3345.000 1431.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1479.770 3345.000 1482.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1530.970 3345.000 1534.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1582.170 3345.000 1585.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.370 3345.000 1636.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.570 3345.000 1687.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.770 3345.000 1738.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.970 3345.000 1790.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1838.170 3345.000 1841.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1889.370 3345.000 1892.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1940.570 3345.000 1943.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.770 3345.000 1994.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2042.970 3345.000 2046.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.170 3345.000 2097.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.370 3345.000 2148.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2196.570 3345.000 2199.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2247.770 3345.000 2250.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2298.970 3345.000 2302.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2350.170 3345.000 2353.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.370 3345.000 2404.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2452.570 3345.000 2455.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2503.770 3345.000 2506.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.970 3345.000 2558.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2606.170 3345.000 2609.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2657.370 3345.000 2660.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.570 3345.000 2711.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2759.770 -28.670 2762.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2810.970 -28.670 2814.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2862.170 -28.670 2865.270 3548.350 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.130 2963.250 253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.130 2963.250 433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.130 2963.250 613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 167.170 -38.270 170.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.370 -38.270 221.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.570 -38.270 272.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.770 -38.270 323.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.970 -38.270 375.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.170 -38.270 426.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.370 -38.270 477.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.570 -38.270 528.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.770 -38.270 579.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.970 -38.270 631.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.170 -38.270 682.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 730.370 -38.270 733.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 781.570 -38.270 784.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.770 -38.270 835.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 883.970 -38.270 887.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.170 -38.270 938.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 986.370 -38.270 989.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1037.570 -38.270 1040.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.770 -38.270 1091.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1139.970 -38.270 1143.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1191.170 -38.270 1194.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1242.370 -38.270 1245.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.570 -38.270 1296.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1344.770 -38.270 1347.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.970 -38.270 1399.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1447.170 -38.270 1450.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1498.370 -38.270 1501.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1549.570 -38.270 1552.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1600.770 -38.270 1603.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.970 -38.270 1655.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1703.170 -38.270 1706.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1754.370 -38.270 1757.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1805.570 -38.270 1808.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.770 -38.270 1859.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1907.970 -38.270 1911.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1959.170 -38.270 1962.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2010.370 -38.270 2013.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.570 -38.270 2064.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2112.770 -38.270 2115.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.970 -38.270 2167.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.170 -38.270 2218.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2266.370 -38.270 2269.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2317.570 -38.270 2320.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2368.770 -38.270 2371.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2419.970 -38.270 2423.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2471.170 -38.270 2474.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2522.370 -38.270 2525.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2573.570 -38.270 2576.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.770 -38.270 2627.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2675.970 -38.270 2679.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.170 -38.270 2730.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.970 -38.270 119.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 167.170 3345.000 170.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.370 3345.000 221.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.570 3345.000 272.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.770 3345.000 323.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.970 3345.000 375.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.170 3345.000 426.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.370 3345.000 477.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.570 3345.000 528.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.770 3345.000 579.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.970 3345.000 631.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.170 3345.000 682.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 730.370 3345.000 733.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 781.570 3345.000 784.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.770 3345.000 835.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 883.970 3345.000 887.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.170 3345.000 938.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 986.370 3345.000 989.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1037.570 3345.000 1040.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.770 3345.000 1091.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1139.970 3345.000 1143.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1191.170 3345.000 1194.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1242.370 3345.000 1245.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.570 3345.000 1296.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1344.770 3345.000 1347.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.970 3345.000 1399.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1447.170 3345.000 1450.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1498.370 3345.000 1501.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1549.570 3345.000 1552.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1600.770 3345.000 1603.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.970 3345.000 1655.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1703.170 3345.000 1706.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1754.370 3345.000 1757.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1805.570 3345.000 1808.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.770 3345.000 1859.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1907.970 3345.000 1911.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1959.170 3345.000 1962.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2010.370 3345.000 2013.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.570 3345.000 2064.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2112.770 3345.000 2115.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.970 3345.000 2167.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.170 3345.000 2218.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2266.370 3345.000 2269.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2317.570 3345.000 2320.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2368.770 3345.000 2371.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2419.970 3345.000 2423.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2471.170 3345.000 2474.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2522.370 3345.000 2525.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2573.570 3345.000 2576.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.770 3345.000 2627.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2675.970 3345.000 2679.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.170 3345.000 2730.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2778.370 -38.270 2781.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.570 -38.270 2832.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2880.770 -38.270 2883.870 3557.950 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 141.530 2953.650 144.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 321.530 2953.650 324.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 501.530 2953.650 504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 681.530 2953.650 684.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 861.530 2953.650 864.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.170 -28.670 177.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.370 -28.670 228.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.570 -28.670 279.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.770 -28.670 330.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.970 -28.670 382.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 430.170 -28.670 433.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.370 -28.670 484.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.570 -28.670 535.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 583.770 -28.670 586.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 634.970 -28.670 638.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 686.170 -28.670 689.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 737.370 -28.670 740.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 788.570 -28.670 791.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 839.770 -28.670 842.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 890.970 -28.670 894.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.170 -28.670 945.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 993.370 -28.670 996.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1044.570 -28.670 1047.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.770 -28.670 1098.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.970 -28.670 1150.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.170 -28.670 1201.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.370 -28.670 1252.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.570 -28.670 1303.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1351.770 -28.670 1354.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1402.970 -28.670 1406.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.170 -28.670 1457.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1505.370 -28.670 1508.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1556.570 -28.670 1559.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1607.770 -28.670 1610.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.970 -28.670 1662.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.170 -28.670 1713.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1761.370 -28.670 1764.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1812.570 -28.670 1815.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1863.770 -28.670 1866.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1914.970 -28.670 1918.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.170 -28.670 1969.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.370 -28.670 2020.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2068.570 -28.670 2071.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2119.770 -28.670 2122.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2170.970 -28.670 2174.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2222.170 -28.670 2225.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2273.370 -28.670 2276.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2324.570 -28.670 2327.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.770 -28.670 2378.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.970 -28.670 2430.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.170 -28.670 2481.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2529.370 -28.670 2532.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2580.570 -28.670 2583.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.770 -28.670 2634.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2682.970 -28.670 2686.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2734.170 -28.670 2737.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.770 -28.670 74.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.970 -28.670 126.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.170 3345.000 177.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.370 3345.000 228.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.570 3345.000 279.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.770 3345.000 330.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.970 3345.000 382.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 430.170 3345.000 433.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.370 3345.000 484.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.570 3345.000 535.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 583.770 3345.000 586.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 634.970 3345.000 638.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 686.170 3345.000 689.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 737.370 3345.000 740.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 788.570 3345.000 791.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 839.770 3345.000 842.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 890.970 3345.000 894.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.170 3345.000 945.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 993.370 3345.000 996.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1044.570 3345.000 1047.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.770 3345.000 1098.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.970 3345.000 1150.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.170 3345.000 1201.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.370 3345.000 1252.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.570 3345.000 1303.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1351.770 3345.000 1354.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1402.970 3345.000 1406.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.170 3345.000 1457.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1505.370 3345.000 1508.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1556.570 3345.000 1559.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1607.770 3345.000 1610.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.970 3345.000 1662.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.170 3345.000 1713.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1761.370 3345.000 1764.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1812.570 3345.000 1815.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1863.770 3345.000 1866.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1914.970 3345.000 1918.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.170 3345.000 1969.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.370 3345.000 2020.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2068.570 3345.000 2071.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2119.770 3345.000 2122.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2170.970 3345.000 2174.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2222.170 3345.000 2225.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2273.370 3345.000 2276.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2324.570 3345.000 2327.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.770 3345.000 2378.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2426.970 3345.000 2430.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.170 3345.000 2481.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2529.370 3345.000 2532.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2580.570 3345.000 2583.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.770 3345.000 2634.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2682.970 3345.000 2686.070 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2734.170 3345.000 2737.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.370 -28.670 2788.470 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.570 -28.670 2839.670 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2887.770 -28.670 2890.870 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 160.130 2963.250 163.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 340.130 2963.250 343.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 520.130 2963.250 523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 700.130 2963.250 703.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 880.130 2963.250 883.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.570 -38.270 144.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 192.770 -38.270 195.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.970 -38.270 247.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 295.170 -38.270 298.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.370 -38.270 349.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 397.570 -38.270 400.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.770 -38.270 451.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 499.970 -38.270 503.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 551.170 -38.270 554.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 602.370 -38.270 605.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.570 -38.270 656.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.770 -38.270 707.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 755.970 -38.270 759.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.170 -38.270 810.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.370 -38.270 861.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 909.570 -38.270 912.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 960.770 -38.270 963.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.970 -38.270 1015.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1063.170 -38.270 1066.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.370 -38.270 1117.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.570 -38.270 1168.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.770 -38.270 1219.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1267.970 -38.270 1271.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1319.170 -38.270 1322.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1370.370 -38.270 1373.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.570 -38.270 1424.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.770 -38.270 1475.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.970 -38.270 1527.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.170 -38.270 1578.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1626.370 -38.270 1629.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1677.570 -38.270 1680.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.770 -38.270 1731.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.970 -38.270 1783.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.170 -38.270 1834.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1882.370 -38.270 1885.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.570 -38.270 1936.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.770 -38.270 1987.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.970 -38.270 2039.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2087.170 -38.270 2090.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2138.370 -38.270 2141.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2189.570 -38.270 2192.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.770 -38.270 2243.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2291.970 -38.270 2295.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2343.170 -38.270 2346.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.370 -38.270 2397.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2445.570 -38.270 2448.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.770 -38.270 2499.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.970 -38.270 2551.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2599.170 -38.270 2602.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2650.370 -38.270 2653.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2701.570 -38.270 2704.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2752.770 -38.270 2755.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.370 -38.270 93.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.570 3345.000 144.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 192.770 3345.000 195.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.970 3345.000 247.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 295.170 3345.000 298.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.370 3345.000 349.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 397.570 3345.000 400.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.770 3345.000 451.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 499.970 3345.000 503.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 551.170 3345.000 554.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 602.370 3345.000 605.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.570 3345.000 656.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.770 3345.000 707.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 755.970 3345.000 759.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.170 3345.000 810.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.370 3345.000 861.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 909.570 3345.000 912.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 960.770 3345.000 963.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.970 3345.000 1015.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1063.170 3345.000 1066.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.370 3345.000 1117.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.570 3345.000 1168.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.770 3345.000 1219.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1267.970 3345.000 1271.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1319.170 3345.000 1322.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1370.370 3345.000 1373.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.570 3345.000 1424.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.770 3345.000 1475.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.970 3345.000 1527.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.170 3345.000 1578.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1626.370 3345.000 1629.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1677.570 3345.000 1680.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.770 3345.000 1731.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.970 3345.000 1783.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.170 3345.000 1834.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1882.370 3345.000 1885.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.570 3345.000 1936.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.770 3345.000 1987.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.970 3345.000 2039.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2087.170 3345.000 2090.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2138.370 3345.000 2141.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2189.570 3345.000 2192.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.770 3345.000 2243.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2291.970 3345.000 2295.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2343.170 3345.000 2346.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.370 3345.000 2397.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2445.570 3345.000 2448.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2496.770 3345.000 2499.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.970 3345.000 2551.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2599.170 3345.000 2602.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2650.370 3345.000 2653.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2701.570 3345.000 2704.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2752.770 3345.000 2755.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2803.970 -38.270 2807.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2855.170 -38.270 2858.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2906.370 -38.270 2909.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 104.330 2934.450 107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 284.330 2934.450 287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 464.330 2934.450 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 644.330 2934.450 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 824.330 2934.450 827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1004.330 2934.450 1007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1184.330 2934.450 1187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1364.330 2934.450 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1544.330 2934.450 1547.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1724.330 2934.450 1727.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1904.330 2934.450 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2084.330 2934.450 2087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2264.330 2934.450 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2444.330 2934.450 2447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2624.330 2934.450 2627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2804.330 2934.450 2807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2984.330 2934.450 2987.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3344.330 2934.450 3347.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.970 -9.470 140.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.170 -9.470 191.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.370 -9.470 242.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.570 -9.470 293.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.770 -9.470 344.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 392.970 -9.470 396.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 444.170 -9.470 447.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.370 -9.470 498.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.570 -9.470 549.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 597.770 -9.470 600.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.970 -9.470 652.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.170 -9.470 703.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.370 -9.470 754.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 802.570 -9.470 805.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 853.770 -9.470 856.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.970 -9.470 908.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.170 -9.470 959.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.370 -9.470 1010.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.570 -9.470 1061.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1109.770 -9.470 1112.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1160.970 -9.470 1164.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1212.170 -9.470 1215.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.370 -9.470 1266.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.570 -9.470 1317.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1365.770 -9.470 1368.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1416.970 -9.470 1420.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1468.170 -9.470 1471.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1519.370 -9.470 1522.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1570.570 -9.470 1573.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1621.770 -9.470 1624.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1672.970 -9.470 1676.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1724.170 -9.470 1727.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.370 -9.470 1778.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1826.570 -9.470 1829.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1877.770 -9.470 1880.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1928.970 -9.470 1932.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.170 -9.470 1983.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.370 -9.470 2034.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2082.570 -9.470 2085.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2133.770 -9.470 2136.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.970 -9.470 2188.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.170 -9.470 2239.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2287.370 -9.470 2290.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2338.570 -9.470 2341.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2389.770 -9.470 2392.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2440.970 -9.470 2444.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2492.170 -9.470 2495.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2543.370 -9.470 2546.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2594.570 -9.470 2597.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2645.770 -9.470 2648.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2696.970 -9.470 2700.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2748.170 -9.470 2751.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.570 -9.470 37.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.770 -9.470 88.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.970 3345.000 140.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.170 3345.000 191.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.370 3345.000 242.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.570 3345.000 293.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.770 3345.000 344.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 392.970 3345.000 396.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 444.170 3345.000 447.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.370 3345.000 498.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.570 3345.000 549.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 597.770 3345.000 600.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.970 3345.000 652.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.170 3345.000 703.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.370 3345.000 754.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 802.570 3345.000 805.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 853.770 3345.000 856.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.970 3345.000 908.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.170 3345.000 959.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.370 3345.000 1010.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.570 3345.000 1061.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1109.770 3345.000 1112.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1160.970 3345.000 1164.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1212.170 3345.000 1215.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.370 3345.000 1266.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.570 3345.000 1317.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1365.770 3345.000 1368.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1416.970 3345.000 1420.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1468.170 3345.000 1471.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1519.370 3345.000 1522.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1570.570 3345.000 1573.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1621.770 3345.000 1624.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1672.970 3345.000 1676.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1724.170 3345.000 1727.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.370 3345.000 1778.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1826.570 3345.000 1829.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1877.770 3345.000 1880.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1928.970 3345.000 1932.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.170 3345.000 1983.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.370 3345.000 2034.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2082.570 3345.000 2085.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2133.770 3345.000 2136.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.970 3345.000 2188.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.170 3345.000 2239.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2287.370 3345.000 2290.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2338.570 3345.000 2341.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2389.770 3345.000 2392.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2440.970 3345.000 2444.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2492.170 3345.000 2495.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2543.370 3345.000 2546.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2594.570 3345.000 2597.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2645.770 3345.000 2648.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2696.970 3345.000 2700.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2748.170 3345.000 2751.270 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2799.370 -9.470 2802.470 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2850.570 -9.470 2853.670 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2901.770 -9.470 2904.870 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 122.930 2944.050 126.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 302.930 2944.050 306.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 482.930 2944.050 486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 662.930 2944.050 666.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 842.930 2944.050 846.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 155.570 -19.070 158.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 206.770 -19.070 209.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 257.970 -19.070 261.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.170 -19.070 312.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 360.370 -19.070 363.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.570 -19.070 414.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 462.770 -19.070 465.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.970 -19.070 517.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.170 -19.070 568.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.370 -19.070 619.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 667.570 -19.070 670.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 718.770 -19.070 721.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 769.970 -19.070 773.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.170 -19.070 824.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 872.370 -19.070 875.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.570 -19.070 926.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.770 -19.070 977.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.970 -19.070 1029.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.170 -19.070 1080.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.370 -19.070 1131.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1179.570 -19.070 1182.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1230.770 -19.070 1233.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.970 -19.070 1285.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1333.170 -19.070 1336.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1384.370 -19.070 1387.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.570 -19.070 1438.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.770 -19.070 1489.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1537.970 -19.070 1541.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1589.170 -19.070 1592.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1640.370 -19.070 1643.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1691.570 -19.070 1694.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1742.770 -19.070 1745.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1793.970 -19.070 1797.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1845.170 -19.070 1848.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1896.370 -19.070 1899.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.570 -19.070 1950.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1998.770 -19.070 2001.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2049.970 -19.070 2053.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2101.170 -19.070 2104.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.370 -19.070 2155.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2203.570 -19.070 2206.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.770 -19.070 2257.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2305.970 -19.070 2309.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2357.170 -19.070 2360.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.370 -19.070 2411.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2459.570 -19.070 2462.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2510.770 -19.070 2513.870 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2561.970 -19.070 2565.070 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2613.170 -19.070 2616.270 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.370 -19.070 2667.470 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2715.570 -19.070 2718.670 125.000 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.170 -19.070 56.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.370 -19.070 107.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 155.570 3345.000 158.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 206.770 3345.000 209.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 257.970 3345.000 261.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.170 3345.000 312.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 360.370 3345.000 363.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.570 3345.000 414.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 462.770 3345.000 465.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.970 3345.000 517.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.170 3345.000 568.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.370 3345.000 619.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 667.570 3345.000 670.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 718.770 3345.000 721.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 769.970 3345.000 773.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.170 3345.000 824.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 872.370 3345.000 875.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.570 3345.000 926.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.770 3345.000 977.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.970 3345.000 1029.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.170 3345.000 1080.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.370 3345.000 1131.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1179.570 3345.000 1182.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1230.770 3345.000 1233.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.970 3345.000 1285.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1333.170 3345.000 1336.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1384.370 3345.000 1387.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.570 3345.000 1438.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.770 3345.000 1489.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1537.970 3345.000 1541.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1589.170 3345.000 1592.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1640.370 3345.000 1643.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1691.570 3345.000 1694.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1742.770 3345.000 1745.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1793.970 3345.000 1797.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1845.170 3345.000 1848.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1896.370 3345.000 1899.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.570 3345.000 1950.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1998.770 3345.000 2001.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2049.970 3345.000 2053.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2101.170 3345.000 2104.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.370 3345.000 2155.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2203.570 3345.000 2206.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.770 3345.000 2257.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2305.970 3345.000 2309.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2357.170 3345.000 2360.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.370 3345.000 2411.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2459.570 3345.000 2462.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2510.770 3345.000 2513.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2561.970 3345.000 2565.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2613.170 3345.000 2616.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.370 3345.000 2667.470 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2715.570 3345.000 2718.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2766.770 -19.070 2769.870 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.970 -19.070 2821.070 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2869.170 -19.070 2872.270 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 152.120 145.795 2741.000 3322.925 ;
      LAYER met1 ;
        RECT 13.870 103.060 2903.450 3515.220 ;
      LAYER met2 ;
        RECT 13.890 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2903.430 3518.050 ;
        RECT 13.890 98.755 2903.430 3517.320 ;
      LAYER met3 ;
        RECT 2.800 3485.700 2917.200 3486.185 ;
        RECT 2.400 3485.020 2917.200 3485.700 ;
        RECT 2.400 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 2.400 3420.380 2917.600 3420.420 ;
        RECT 2.400 3418.380 2917.200 3420.380 ;
        RECT 2.400 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 2.400 3354.420 2917.600 3355.140 ;
        RECT 2.400 3352.420 2917.200 3354.420 ;
        RECT 2.400 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 2.400 3287.780 2917.600 3289.860 ;
        RECT 2.400 3285.780 2917.200 3287.780 ;
        RECT 2.400 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 2.400 3221.140 2917.600 3224.580 ;
        RECT 2.400 3219.140 2917.200 3221.140 ;
        RECT 2.400 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 2.400 3155.180 2917.600 3159.300 ;
        RECT 2.400 3153.180 2917.200 3155.180 ;
        RECT 2.400 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 2.400 3088.540 2917.600 3094.700 ;
        RECT 2.400 3086.540 2917.200 3088.540 ;
        RECT 2.400 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 2.400 3021.900 2917.600 3029.420 ;
        RECT 2.400 3019.900 2917.200 3021.900 ;
        RECT 2.400 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 2.400 2955.940 2917.600 2964.140 ;
        RECT 2.400 2953.940 2917.200 2955.940 ;
        RECT 2.400 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 2.400 2889.300 2917.600 2898.860 ;
        RECT 2.400 2887.300 2917.200 2889.300 ;
        RECT 2.400 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 2.400 2822.660 2917.600 2833.580 ;
        RECT 2.400 2820.660 2917.200 2822.660 ;
        RECT 2.400 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 2.400 2756.700 2917.600 2768.300 ;
        RECT 2.400 2754.700 2917.200 2756.700 ;
        RECT 2.400 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 2.400 2690.060 2917.600 2703.020 ;
        RECT 2.400 2688.060 2917.200 2690.060 ;
        RECT 2.400 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 2.400 2623.420 2917.600 2638.420 ;
        RECT 2.400 2621.420 2917.200 2623.420 ;
        RECT 2.400 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 2.400 2557.460 2917.600 2573.140 ;
        RECT 2.400 2555.460 2917.200 2557.460 ;
        RECT 2.400 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 2.400 2490.820 2917.600 2507.860 ;
        RECT 2.400 2488.820 2917.200 2490.820 ;
        RECT 2.400 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 2.400 2424.180 2917.600 2442.580 ;
        RECT 2.400 2422.180 2917.200 2424.180 ;
        RECT 2.400 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 2.400 2358.220 2917.600 2377.300 ;
        RECT 2.400 2356.220 2917.200 2358.220 ;
        RECT 2.400 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 2.400 2291.580 2917.600 2312.020 ;
        RECT 2.400 2289.580 2917.200 2291.580 ;
        RECT 2.400 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 2.400 2224.940 2917.600 2246.740 ;
        RECT 2.400 2222.940 2917.200 2224.940 ;
        RECT 2.400 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 2.400 2158.980 2917.600 2182.140 ;
        RECT 2.400 2156.980 2917.200 2158.980 ;
        RECT 2.400 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 2.400 2092.340 2917.600 2116.860 ;
        RECT 2.400 2090.340 2917.200 2092.340 ;
        RECT 2.400 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 2.400 2025.700 2917.600 2051.580 ;
        RECT 2.400 2023.700 2917.200 2025.700 ;
        RECT 2.400 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 2.400 1959.740 2917.600 1986.300 ;
        RECT 2.400 1957.740 2917.200 1959.740 ;
        RECT 2.400 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 2.400 1893.100 2917.600 1921.020 ;
        RECT 2.400 1891.100 2917.200 1893.100 ;
        RECT 2.400 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.400 1826.460 2917.600 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.400 1760.500 2917.600 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 2.400 1693.860 2917.600 1725.860 ;
        RECT 2.400 1691.860 2917.200 1693.860 ;
        RECT 2.400 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 2.400 1627.220 2917.600 1660.580 ;
        RECT 2.400 1625.220 2917.200 1627.220 ;
        RECT 2.400 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 2.400 1561.260 2917.600 1595.300 ;
        RECT 2.400 1559.260 2917.200 1561.260 ;
        RECT 2.400 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 2.400 1494.620 2917.600 1530.020 ;
        RECT 2.400 1492.620 2917.200 1494.620 ;
        RECT 2.400 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 2.400 1427.980 2917.600 1464.740 ;
        RECT 2.400 1425.980 2917.200 1427.980 ;
        RECT 2.400 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 2.400 1362.020 2917.600 1399.460 ;
        RECT 2.400 1360.020 2917.200 1362.020 ;
        RECT 2.400 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 2.400 1295.380 2917.600 1334.860 ;
        RECT 2.400 1293.380 2917.200 1295.380 ;
        RECT 2.400 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 2.400 1228.740 2917.600 1269.580 ;
        RECT 2.400 1226.740 2917.200 1228.740 ;
        RECT 2.400 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 2.400 1162.780 2917.600 1204.300 ;
        RECT 2.400 1160.780 2917.200 1162.780 ;
        RECT 2.400 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 2.400 1096.140 2917.600 1139.020 ;
        RECT 2.400 1094.140 2917.200 1096.140 ;
        RECT 2.400 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 2.400 1029.500 2917.600 1073.740 ;
        RECT 2.400 1027.500 2917.200 1029.500 ;
        RECT 2.400 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 2.400 963.540 2917.600 1008.460 ;
        RECT 2.400 961.540 2917.200 963.540 ;
        RECT 2.400 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 2.400 896.900 2917.600 943.180 ;
        RECT 2.400 894.900 2917.200 896.900 ;
        RECT 2.400 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 2.400 830.260 2917.600 878.580 ;
        RECT 2.400 828.260 2917.200 830.260 ;
        RECT 2.400 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 2.400 764.300 2917.600 813.300 ;
        RECT 2.400 762.300 2917.200 764.300 ;
        RECT 2.400 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 2.400 697.660 2917.600 748.020 ;
        RECT 2.400 695.660 2917.200 697.660 ;
        RECT 2.400 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 2.400 631.020 2917.600 682.740 ;
        RECT 2.400 629.020 2917.200 631.020 ;
        RECT 2.400 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 2.400 565.060 2917.600 617.460 ;
        RECT 2.400 563.060 2917.200 565.060 ;
        RECT 2.400 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 2.400 498.420 2917.600 552.180 ;
        RECT 2.400 496.420 2917.200 498.420 ;
        RECT 2.400 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 2.400 431.780 2917.600 486.900 ;
        RECT 2.400 429.780 2917.200 431.780 ;
        RECT 2.400 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 2.400 365.820 2917.600 422.300 ;
        RECT 2.400 363.820 2917.200 365.820 ;
        RECT 2.400 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 2.400 299.180 2917.600 357.020 ;
        RECT 2.400 297.180 2917.200 299.180 ;
        RECT 2.400 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 2.400 232.540 2917.600 291.740 ;
        RECT 2.400 230.540 2917.200 232.540 ;
        RECT 2.400 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 2.400 166.580 2917.600 226.460 ;
        RECT 2.400 164.580 2917.200 166.580 ;
        RECT 2.400 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 2.400 99.940 2917.600 161.180 ;
        RECT 2.400 98.775 2917.200 99.940 ;
      LAYER met4 ;
        RECT 166.215 145.640 2733.345 3323.080 ;
  END
END user_project_wrapper
END LIBRARY

